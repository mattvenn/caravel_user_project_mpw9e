VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO rgb_mixer
  CLASS BLOCK ;
  FOREIGN rgb_mixer ;
  ORIGIN 0.000 0.000 ;
  SIZE 180.000 BY 210.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 144.850 206.000 145.410 210.000 ;
    END
  END clk
  PIN enc0_a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 74.010 206.000 74.570 210.000 ;
    END
  END enc0_a
  PIN enc0_b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 176.000 173.140 180.000 174.340 ;
    END
  END enc0_b
  PIN enc1_a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 176.000 64.340 180.000 65.540 ;
    END
  END enc1_a
  PIN enc1_b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 41.810 206.000 42.370 210.000 ;
    END
  END enc1_b
  PIN enc2_a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 142.540 4.000 143.740 ;
    END
  END enc2_a
  PIN enc2_b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 71.140 4.000 72.340 ;
    END
  END enc2_b
  PIN io_oeb_high[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 176.000 26.940 180.000 28.140 ;
    END
  END io_oeb_high[0]
  PIN io_oeb_high[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.190 0.000 135.750 4.000 ;
    END
  END io_oeb_high[1]
  PIN io_oeb_high[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT -0.050 0.000 0.510 4.000 ;
    END
  END io_oeb_high[2]
  PIN io_oeb_high[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.050 206.000 177.610 210.000 ;
    END
  END io_oeb_high[3]
  PIN io_oeb_high[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.150 0.000 32.710 4.000 ;
    END
  END io_oeb_high[4]
  PIN io_oeb_high[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.610 0.000 171.170 4.000 ;
    END
  END io_oeb_high[5]
  PIN io_oeb_low[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.570 0.000 68.130 4.000 ;
    END
  END io_oeb_low[0]
  PIN io_oeb_low[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 33.740 4.000 34.940 ;
    END
  END io_oeb_low[1]
  PIN io_oeb_low[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 176.000 135.740 180.000 136.940 ;
    END
  END io_oeb_low[2]
  PIN io_oeb_low[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 179.940 4.000 181.140 ;
    END
  END io_oeb_low[3]
  PIN pwm0_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 109.430 206.000 109.990 210.000 ;
    END
  END pwm0_out
  PIN pwm1_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 102.990 0.000 103.550 4.000 ;
    END
  END pwm1_out
  PIN pwm2_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.540 4.000 109.740 ;
    END
  END pwm2_out
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 6.390 206.000 6.950 210.000 ;
    END
  END reset
  PIN sync
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 176.000 98.340 180.000 99.540 ;
    END
  END sync
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 25.820 10.640 27.420 198.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 68.025 10.640 69.625 198.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 110.230 10.640 111.830 198.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 152.435 10.640 154.035 198.800 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 46.920 10.640 48.520 198.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 89.125 10.640 90.725 198.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 131.330 10.640 132.930 198.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 173.535 10.640 175.135 198.800 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 174.340 198.645 ;
      LAYER met1 ;
        RECT 0.070 10.640 177.490 198.800 ;
      LAYER met2 ;
        RECT 0.100 205.720 6.110 206.000 ;
        RECT 7.230 205.720 41.530 206.000 ;
        RECT 42.650 205.720 73.730 206.000 ;
        RECT 74.850 205.720 109.150 206.000 ;
        RECT 110.270 205.720 144.570 206.000 ;
        RECT 145.690 205.720 176.770 206.000 ;
        RECT 0.100 4.280 177.460 205.720 ;
        RECT 0.790 4.000 31.870 4.280 ;
        RECT 32.990 4.000 67.290 4.280 ;
        RECT 68.410 4.000 102.710 4.280 ;
        RECT 103.830 4.000 134.910 4.280 ;
        RECT 136.030 4.000 170.330 4.280 ;
        RECT 171.450 4.000 177.460 4.280 ;
      LAYER met3 ;
        RECT 3.990 181.540 176.100 198.725 ;
        RECT 4.400 179.540 176.100 181.540 ;
        RECT 3.990 174.740 176.100 179.540 ;
        RECT 3.990 172.740 175.600 174.740 ;
        RECT 3.990 144.140 176.100 172.740 ;
        RECT 4.400 142.140 176.100 144.140 ;
        RECT 3.990 137.340 176.100 142.140 ;
        RECT 3.990 135.340 175.600 137.340 ;
        RECT 3.990 110.140 176.100 135.340 ;
        RECT 4.400 108.140 176.100 110.140 ;
        RECT 3.990 99.940 176.100 108.140 ;
        RECT 3.990 97.940 175.600 99.940 ;
        RECT 3.990 72.740 176.100 97.940 ;
        RECT 4.400 70.740 176.100 72.740 ;
        RECT 3.990 65.940 176.100 70.740 ;
        RECT 3.990 63.940 175.600 65.940 ;
        RECT 3.990 35.340 176.100 63.940 ;
        RECT 4.400 33.340 176.100 35.340 ;
        RECT 3.990 28.540 176.100 33.340 ;
        RECT 3.990 26.540 175.600 28.540 ;
        RECT 3.990 10.715 176.100 26.540 ;
  END
END rgb_mixer
END LIBRARY

