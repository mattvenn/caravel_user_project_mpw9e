// This is the unpowered netlist.
module rgb_mixer (clk,
    enc0_a,
    enc0_b,
    enc1_a,
    enc1_b,
    enc2_a,
    enc2_b,
    pwm0_out,
    pwm1_out,
    pwm2_out,
    reset,
    sync,
    io_oeb_high,
    io_oeb_low);
 input clk;
 input enc0_a;
 input enc0_b;
 input enc1_a;
 input enc1_b;
 input enc2_a;
 input enc2_b;
 output pwm0_out;
 output pwm1_out;
 output pwm2_out;
 input reset;
 output sync;
 output [5:0] io_oeb_high;
 output [3:0] io_oeb_low;

 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire _277_;
 wire _278_;
 wire _279_;
 wire _280_;
 wire _281_;
 wire _282_;
 wire _283_;
 wire _284_;
 wire _285_;
 wire _286_;
 wire _287_;
 wire _288_;
 wire _289_;
 wire _290_;
 wire _291_;
 wire _292_;
 wire _293_;
 wire _294_;
 wire _295_;
 wire _296_;
 wire _297_;
 wire _298_;
 wire _299_;
 wire _300_;
 wire _301_;
 wire _302_;
 wire _303_;
 wire _304_;
 wire _305_;
 wire _306_;
 wire _307_;
 wire _308_;
 wire _309_;
 wire _310_;
 wire _311_;
 wire _312_;
 wire _313_;
 wire _314_;
 wire _315_;
 wire _316_;
 wire _317_;
 wire _318_;
 wire _319_;
 wire _320_;
 wire _321_;
 wire _322_;
 wire _323_;
 wire _324_;
 wire _325_;
 wire _326_;
 wire _327_;
 wire _328_;
 wire _329_;
 wire _330_;
 wire _331_;
 wire _332_;
 wire _333_;
 wire _334_;
 wire _335_;
 wire _336_;
 wire _337_;
 wire _338_;
 wire _339_;
 wire _340_;
 wire _341_;
 wire _342_;
 wire _343_;
 wire _344_;
 wire _345_;
 wire _346_;
 wire _347_;
 wire _348_;
 wire _349_;
 wire _350_;
 wire _351_;
 wire _352_;
 wire _353_;
 wire _354_;
 wire _355_;
 wire _356_;
 wire _357_;
 wire _358_;
 wire _359_;
 wire _360_;
 wire _361_;
 wire _362_;
 wire _363_;
 wire _364_;
 wire _365_;
 wire _366_;
 wire _367_;
 wire _368_;
 wire _369_;
 wire _370_;
 wire _371_;
 wire _372_;
 wire _373_;
 wire _374_;
 wire _375_;
 wire _376_;
 wire _377_;
 wire _378_;
 wire _379_;
 wire _380_;
 wire _381_;
 wire _382_;
 wire _383_;
 wire _384_;
 wire _385_;
 wire _386_;
 wire _387_;
 wire _388_;
 wire _389_;
 wire _390_;
 wire _391_;
 wire _392_;
 wire _393_;
 wire _394_;
 wire _395_;
 wire _396_;
 wire _397_;
 wire _398_;
 wire _399_;
 wire _400_;
 wire _401_;
 wire _402_;
 wire _403_;
 wire _404_;
 wire _405_;
 wire _406_;
 wire _407_;
 wire _408_;
 wire _409_;
 wire _410_;
 wire _411_;
 wire _412_;
 wire _413_;
 wire _414_;
 wire _415_;
 wire _416_;
 wire _417_;
 wire _418_;
 wire _419_;
 wire _420_;
 wire _421_;
 wire _422_;
 wire _423_;
 wire _424_;
 wire _425_;
 wire clknet_0_clk;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire \debounce0_a.button_hist[0] ;
 wire \debounce0_a.button_hist[1] ;
 wire \debounce0_a.button_hist[2] ;
 wire \debounce0_a.button_hist[3] ;
 wire \debounce0_a.button_hist[4] ;
 wire \debounce0_a.button_hist[5] ;
 wire \debounce0_a.button_hist[6] ;
 wire \debounce0_a.button_hist[7] ;
 wire \debounce0_a.debounced ;
 wire \debounce0_a.reset ;
 wire \debounce0_b.button_hist[0] ;
 wire \debounce0_b.button_hist[1] ;
 wire \debounce0_b.button_hist[2] ;
 wire \debounce0_b.button_hist[3] ;
 wire \debounce0_b.button_hist[4] ;
 wire \debounce0_b.button_hist[5] ;
 wire \debounce0_b.button_hist[6] ;
 wire \debounce0_b.button_hist[7] ;
 wire \debounce0_b.debounced ;
 wire \debounce1_a.button_hist[0] ;
 wire \debounce1_a.button_hist[1] ;
 wire \debounce1_a.button_hist[2] ;
 wire \debounce1_a.button_hist[3] ;
 wire \debounce1_a.button_hist[4] ;
 wire \debounce1_a.button_hist[5] ;
 wire \debounce1_a.button_hist[6] ;
 wire \debounce1_a.button_hist[7] ;
 wire \debounce1_a.debounced ;
 wire \debounce1_b.button_hist[0] ;
 wire \debounce1_b.button_hist[1] ;
 wire \debounce1_b.button_hist[2] ;
 wire \debounce1_b.button_hist[3] ;
 wire \debounce1_b.button_hist[4] ;
 wire \debounce1_b.button_hist[5] ;
 wire \debounce1_b.button_hist[6] ;
 wire \debounce1_b.button_hist[7] ;
 wire \debounce1_b.debounced ;
 wire \debounce2_a.button_hist[0] ;
 wire \debounce2_a.button_hist[1] ;
 wire \debounce2_a.button_hist[2] ;
 wire \debounce2_a.button_hist[3] ;
 wire \debounce2_a.button_hist[4] ;
 wire \debounce2_a.button_hist[5] ;
 wire \debounce2_a.button_hist[6] ;
 wire \debounce2_a.button_hist[7] ;
 wire \debounce2_a.debounced ;
 wire \debounce2_b.button_hist[0] ;
 wire \debounce2_b.button_hist[1] ;
 wire \debounce2_b.button_hist[2] ;
 wire \debounce2_b.button_hist[3] ;
 wire \debounce2_b.button_hist[4] ;
 wire \debounce2_b.button_hist[5] ;
 wire \debounce2_b.button_hist[6] ;
 wire \debounce2_b.button_hist[7] ;
 wire \debounce2_b.debounced ;
 wire \encoder0.old_a ;
 wire \encoder0.old_b ;
 wire \encoder0.value[0] ;
 wire \encoder0.value[1] ;
 wire \encoder0.value[2] ;
 wire \encoder0.value[3] ;
 wire \encoder0.value[4] ;
 wire \encoder0.value[5] ;
 wire \encoder0.value[6] ;
 wire \encoder0.value[7] ;
 wire \encoder1.old_a ;
 wire \encoder1.old_b ;
 wire \encoder1.value[0] ;
 wire \encoder1.value[1] ;
 wire \encoder1.value[2] ;
 wire \encoder1.value[3] ;
 wire \encoder1.value[4] ;
 wire \encoder1.value[5] ;
 wire \encoder1.value[6] ;
 wire \encoder1.value[7] ;
 wire \encoder2.old_a ;
 wire \encoder2.old_b ;
 wire \encoder2.value[0] ;
 wire \encoder2.value[1] ;
 wire \encoder2.value[2] ;
 wire \encoder2.value[3] ;
 wire \encoder2.value[4] ;
 wire \encoder2.value[5] ;
 wire \encoder2.value[6] ;
 wire \encoder2.value[7] ;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net2;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net3;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net4;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net5;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire \pwm0.count[0] ;
 wire \pwm0.count[1] ;
 wire \pwm0.count[2] ;
 wire \pwm0.count[3] ;
 wire \pwm0.count[4] ;
 wire \pwm0.count[5] ;
 wire \pwm0.count[6] ;
 wire \pwm0.count[7] ;
 wire \pwm1.count[0] ;
 wire \pwm1.count[1] ;
 wire \pwm1.count[2] ;
 wire \pwm1.count[3] ;
 wire \pwm1.count[4] ;
 wire \pwm1.count[5] ;
 wire \pwm1.count[6] ;
 wire \pwm1.count[7] ;
 wire \pwm2.count[0] ;
 wire \pwm2.count[1] ;
 wire \pwm2.count[2] ;
 wire \pwm2.count[3] ;
 wire \pwm2.count[4] ;
 wire \pwm2.count[5] ;
 wire \pwm2.count[6] ;
 wire \pwm2.count[7] ;

 sky130_fd_sc_hd__decap_3 FILLER_0_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_18 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_142 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_187 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_174 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_171 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_210 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_184 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_49 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_61 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_168 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_95 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_61 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_87 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_60 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_93 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__inv_2 _427_ (.A(\pwm0.count[7] ),
    .Y(_109_));
 sky130_fd_sc_hd__inv_2 _428_ (.A(\pwm0.count[6] ),
    .Y(_110_));
 sky130_fd_sc_hd__a22o_1 _429_ (.A1(\encoder0.value[7] ),
    .A2(_109_),
    .B1(_110_),
    .B2(\encoder0.value[6] ),
    .X(_111_));
 sky130_fd_sc_hd__inv_2 _430_ (.A(\pwm0.count[5] ),
    .Y(_112_));
 sky130_fd_sc_hd__inv_2 _431_ (.A(\pwm0.count[4] ),
    .Y(_113_));
 sky130_fd_sc_hd__inv_2 _432_ (.A(\pwm0.count[3] ),
    .Y(_114_));
 sky130_fd_sc_hd__inv_2 _433_ (.A(\pwm0.count[2] ),
    .Y(_115_));
 sky130_fd_sc_hd__or2_1 _434_ (.A(\encoder0.value[2] ),
    .B(_115_),
    .X(_116_));
 sky130_fd_sc_hd__inv_2 _435_ (.A(net54),
    .Y(_117_));
 sky130_fd_sc_hd__or2_1 _436_ (.A(\encoder0.value[1] ),
    .B(_117_),
    .X(_118_));
 sky130_fd_sc_hd__inv_2 _437_ (.A(net26),
    .Y(_119_));
 sky130_fd_sc_hd__a22o_1 _438_ (.A1(\encoder0.value[1] ),
    .A2(_117_),
    .B1(_119_),
    .B2(\encoder0.value[0] ),
    .X(_120_));
 sky130_fd_sc_hd__a22o_1 _439_ (.A1(\encoder0.value[2] ),
    .A2(_115_),
    .B1(_118_),
    .B2(_120_),
    .X(_121_));
 sky130_fd_sc_hd__a22o_1 _440_ (.A1(\encoder0.value[3] ),
    .A2(_114_),
    .B1(_116_),
    .B2(_121_),
    .X(_122_));
 sky130_fd_sc_hd__o221a_1 _441_ (.A1(\encoder0.value[4] ),
    .A2(_113_),
    .B1(_114_),
    .B2(\encoder0.value[3] ),
    .C1(_122_),
    .X(_123_));
 sky130_fd_sc_hd__a221o_1 _442_ (.A1(\encoder0.value[5] ),
    .A2(_112_),
    .B1(_113_),
    .B2(\encoder0.value[4] ),
    .C1(_123_),
    .X(_124_));
 sky130_fd_sc_hd__o221a_1 _443_ (.A1(\encoder0.value[6] ),
    .A2(_110_),
    .B1(_112_),
    .B2(\encoder0.value[5] ),
    .C1(_124_),
    .X(_125_));
 sky130_fd_sc_hd__clkbuf_4 _444_ (.A(net68),
    .X(_126_));
 sky130_fd_sc_hd__inv_2 _445_ (.A(_126_),
    .Y(_127_));
 sky130_fd_sc_hd__buf_2 _446_ (.A(_127_),
    .X(_128_));
 sky130_fd_sc_hd__clkbuf_4 _447_ (.A(_128_),
    .X(_129_));
 sky130_fd_sc_hd__o221a_1 _448_ (.A1(\encoder0.value[7] ),
    .A2(_109_),
    .B1(_111_),
    .B2(_125_),
    .C1(_129_),
    .X(net8));
 sky130_fd_sc_hd__inv_2 _449_ (.A(\encoder1.value[7] ),
    .Y(_130_));
 sky130_fd_sc_hd__inv_2 _450_ (.A(net153),
    .Y(_131_));
 sky130_fd_sc_hd__inv_2 _451_ (.A(\encoder1.value[5] ),
    .Y(_132_));
 sky130_fd_sc_hd__inv_2 _452_ (.A(\encoder1.value[4] ),
    .Y(_133_));
 sky130_fd_sc_hd__inv_2 _453_ (.A(\encoder1.value[3] ),
    .Y(_134_));
 sky130_fd_sc_hd__or2_1 _454_ (.A(_134_),
    .B(\pwm1.count[3] ),
    .X(_135_));
 sky130_fd_sc_hd__inv_2 _455_ (.A(\encoder1.value[2] ),
    .Y(_136_));
 sky130_fd_sc_hd__inv_2 _456_ (.A(\encoder1.value[0] ),
    .Y(_137_));
 sky130_fd_sc_hd__inv_2 _457_ (.A(\encoder1.value[1] ),
    .Y(_138_));
 sky130_fd_sc_hd__a21o_1 _458_ (.A1(_138_),
    .A2(\pwm1.count[1] ),
    .B1(\pwm1.count[0] ),
    .X(_139_));
 sky130_fd_sc_hd__o22a_1 _459_ (.A1(_136_),
    .A2(\pwm1.count[2] ),
    .B1(\pwm1.count[1] ),
    .B2(_138_),
    .X(_140_));
 sky130_fd_sc_hd__o21a_1 _460_ (.A1(_137_),
    .A2(_139_),
    .B1(_140_),
    .X(_141_));
 sky130_fd_sc_hd__a221o_1 _461_ (.A1(_134_),
    .A2(\pwm1.count[3] ),
    .B1(\pwm1.count[2] ),
    .B2(_136_),
    .C1(_141_),
    .X(_142_));
 sky130_fd_sc_hd__a22o_1 _462_ (.A1(_133_),
    .A2(\pwm1.count[4] ),
    .B1(_135_),
    .B2(_142_),
    .X(_143_));
 sky130_fd_sc_hd__o221a_1 _463_ (.A1(_132_),
    .A2(\pwm1.count[5] ),
    .B1(\pwm1.count[4] ),
    .B2(_133_),
    .C1(_143_),
    .X(_144_));
 sky130_fd_sc_hd__a221o_1 _464_ (.A1(_131_),
    .A2(\pwm1.count[6] ),
    .B1(\pwm1.count[5] ),
    .B2(_132_),
    .C1(_144_),
    .X(_145_));
 sky130_fd_sc_hd__o221a_1 _465_ (.A1(_130_),
    .A2(\pwm1.count[7] ),
    .B1(\pwm1.count[6] ),
    .B2(_131_),
    .C1(_145_),
    .X(_146_));
 sky130_fd_sc_hd__buf_4 _466_ (.A(_126_),
    .X(_147_));
 sky130_fd_sc_hd__a211oi_4 _467_ (.A1(_130_),
    .A2(\pwm1.count[7] ),
    .B1(_146_),
    .C1(_147_),
    .Y(net9));
 sky130_fd_sc_hd__inv_2 _468_ (.A(\encoder2.value[7] ),
    .Y(_148_));
 sky130_fd_sc_hd__inv_2 _469_ (.A(net159),
    .Y(_149_));
 sky130_fd_sc_hd__inv_2 _470_ (.A(\encoder2.value[5] ),
    .Y(_150_));
 sky130_fd_sc_hd__inv_2 _471_ (.A(\encoder2.value[4] ),
    .Y(_151_));
 sky130_fd_sc_hd__inv_2 _472_ (.A(\encoder2.value[3] ),
    .Y(_152_));
 sky130_fd_sc_hd__or2_1 _473_ (.A(_152_),
    .B(\pwm2.count[3] ),
    .X(_153_));
 sky130_fd_sc_hd__inv_2 _474_ (.A(\encoder2.value[2] ),
    .Y(_154_));
 sky130_fd_sc_hd__inv_2 _475_ (.A(\encoder2.value[0] ),
    .Y(_155_));
 sky130_fd_sc_hd__inv_2 _476_ (.A(\encoder2.value[1] ),
    .Y(_156_));
 sky130_fd_sc_hd__a21o_1 _477_ (.A1(_156_),
    .A2(\pwm2.count[1] ),
    .B1(\pwm2.count[0] ),
    .X(_157_));
 sky130_fd_sc_hd__o22a_1 _478_ (.A1(_154_),
    .A2(\pwm2.count[2] ),
    .B1(\pwm2.count[1] ),
    .B2(_156_),
    .X(_158_));
 sky130_fd_sc_hd__o21a_1 _479_ (.A1(_155_),
    .A2(_157_),
    .B1(_158_),
    .X(_159_));
 sky130_fd_sc_hd__a221o_1 _480_ (.A1(_152_),
    .A2(\pwm2.count[3] ),
    .B1(\pwm2.count[2] ),
    .B2(_154_),
    .C1(_159_),
    .X(_160_));
 sky130_fd_sc_hd__a22o_1 _481_ (.A1(_151_),
    .A2(\pwm2.count[4] ),
    .B1(_153_),
    .B2(_160_),
    .X(_161_));
 sky130_fd_sc_hd__o221a_1 _482_ (.A1(_150_),
    .A2(\pwm2.count[5] ),
    .B1(\pwm2.count[4] ),
    .B2(_151_),
    .C1(_161_),
    .X(_162_));
 sky130_fd_sc_hd__a221o_1 _483_ (.A1(_149_),
    .A2(\pwm2.count[6] ),
    .B1(\pwm2.count[5] ),
    .B2(_150_),
    .C1(_162_),
    .X(_163_));
 sky130_fd_sc_hd__o221a_1 _484_ (.A1(_148_),
    .A2(\pwm2.count[7] ),
    .B1(\pwm2.count[6] ),
    .B2(_149_),
    .C1(_163_),
    .X(_164_));
 sky130_fd_sc_hd__a211oi_2 _485_ (.A1(_148_),
    .A2(\pwm2.count[7] ),
    .B1(_164_),
    .C1(_147_),
    .Y(net10));
 sky130_fd_sc_hd__inv_2 _486_ (.A(net24),
    .Y(_000_));
 sky130_fd_sc_hd__or4_1 _487_ (.A(\debounce0_a.button_hist[1] ),
    .B(\debounce0_a.button_hist[0] ),
    .C(\debounce0_a.button_hist[3] ),
    .D(\debounce0_a.button_hist[2] ),
    .X(_165_));
 sky130_fd_sc_hd__o41a_1 _488_ (.A1(\debounce0_a.button_hist[4] ),
    .A2(\debounce0_a.button_hist[7] ),
    .A3(\debounce0_a.button_hist[6] ),
    .A4(_165_),
    .B1(\debounce0_a.debounced ),
    .X(_166_));
 sky130_fd_sc_hd__and4_1 _489_ (.A(\debounce0_a.button_hist[1] ),
    .B(\debounce0_a.button_hist[0] ),
    .C(\debounce0_a.button_hist[3] ),
    .D(\debounce0_a.button_hist[2] ),
    .X(_167_));
 sky130_fd_sc_hd__a41o_1 _490_ (.A1(\debounce0_a.button_hist[4] ),
    .A2(\debounce0_a.button_hist[7] ),
    .A3(\debounce0_a.button_hist[6] ),
    .A4(_167_),
    .B1(\debounce0_a.debounced ),
    .X(_168_));
 sky130_fd_sc_hd__clkbuf_4 _491_ (.A(_128_),
    .X(_169_));
 sky130_fd_sc_hd__o211a_1 _492_ (.A1(net36),
    .A2(_166_),
    .B1(_168_),
    .C1(_169_),
    .X(_001_));
 sky130_fd_sc_hd__clkbuf_4 _493_ (.A(_128_),
    .X(_170_));
 sky130_fd_sc_hd__and2_1 _494_ (.A(_170_),
    .B(net1),
    .X(_171_));
 sky130_fd_sc_hd__clkbuf_1 _495_ (.A(_171_),
    .X(_002_));
 sky130_fd_sc_hd__and2_1 _496_ (.A(net110),
    .B(_170_),
    .X(_172_));
 sky130_fd_sc_hd__clkbuf_1 _497_ (.A(_172_),
    .X(_003_));
 sky130_fd_sc_hd__and2_1 _498_ (.A(net100),
    .B(_170_),
    .X(_173_));
 sky130_fd_sc_hd__clkbuf_1 _499_ (.A(_173_),
    .X(_004_));
 sky130_fd_sc_hd__and2_1 _500_ (.A(net77),
    .B(_170_),
    .X(_174_));
 sky130_fd_sc_hd__clkbuf_1 _501_ (.A(_174_),
    .X(_005_));
 sky130_fd_sc_hd__clkbuf_2 _502_ (.A(_128_),
    .X(_175_));
 sky130_fd_sc_hd__and2_1 _503_ (.A(net89),
    .B(_175_),
    .X(_176_));
 sky130_fd_sc_hd__clkbuf_1 _504_ (.A(_176_),
    .X(_006_));
 sky130_fd_sc_hd__and2_1 _505_ (.A(net117),
    .B(_175_),
    .X(_177_));
 sky130_fd_sc_hd__clkbuf_1 _506_ (.A(_177_),
    .X(_007_));
 sky130_fd_sc_hd__and2_1 _507_ (.A(net36),
    .B(_175_),
    .X(_178_));
 sky130_fd_sc_hd__clkbuf_1 _508_ (.A(_178_),
    .X(_008_));
 sky130_fd_sc_hd__and2_1 _509_ (.A(net137),
    .B(_175_),
    .X(_179_));
 sky130_fd_sc_hd__clkbuf_1 _510_ (.A(_179_),
    .X(_009_));
 sky130_fd_sc_hd__or4_1 _511_ (.A(\debounce0_b.button_hist[1] ),
    .B(\debounce0_b.button_hist[0] ),
    .C(\debounce0_b.button_hist[3] ),
    .D(\debounce0_b.button_hist[2] ),
    .X(_180_));
 sky130_fd_sc_hd__o41a_1 _512_ (.A1(\debounce0_b.button_hist[4] ),
    .A2(\debounce0_b.button_hist[7] ),
    .A3(\debounce0_b.button_hist[6] ),
    .A4(_180_),
    .B1(\debounce0_b.debounced ),
    .X(_181_));
 sky130_fd_sc_hd__and4_1 _513_ (.A(\debounce0_b.button_hist[1] ),
    .B(\debounce0_b.button_hist[0] ),
    .C(\debounce0_b.button_hist[3] ),
    .D(\debounce0_b.button_hist[2] ),
    .X(_182_));
 sky130_fd_sc_hd__a41o_1 _514_ (.A1(\debounce0_b.button_hist[4] ),
    .A2(\debounce0_b.button_hist[7] ),
    .A3(\debounce0_b.button_hist[6] ),
    .A4(_182_),
    .B1(\debounce0_b.debounced ),
    .X(_183_));
 sky130_fd_sc_hd__o211a_1 _515_ (.A1(net32),
    .A2(_181_),
    .B1(_183_),
    .C1(_169_),
    .X(_010_));
 sky130_fd_sc_hd__and2_1 _516_ (.A(_170_),
    .B(net2),
    .X(_184_));
 sky130_fd_sc_hd__clkbuf_1 _517_ (.A(_184_),
    .X(_011_));
 sky130_fd_sc_hd__and2_1 _518_ (.A(net118),
    .B(_175_),
    .X(_185_));
 sky130_fd_sc_hd__clkbuf_1 _519_ (.A(_185_),
    .X(_012_));
 sky130_fd_sc_hd__and2_1 _520_ (.A(net90),
    .B(_175_),
    .X(_186_));
 sky130_fd_sc_hd__clkbuf_1 _521_ (.A(_186_),
    .X(_013_));
 sky130_fd_sc_hd__and2_1 _522_ (.A(net97),
    .B(_175_),
    .X(_187_));
 sky130_fd_sc_hd__clkbuf_1 _523_ (.A(_187_),
    .X(_014_));
 sky130_fd_sc_hd__and2_1 _524_ (.A(net82),
    .B(_175_),
    .X(_188_));
 sky130_fd_sc_hd__clkbuf_1 _525_ (.A(_188_),
    .X(_015_));
 sky130_fd_sc_hd__and2_1 _526_ (.A(net121),
    .B(_175_),
    .X(_189_));
 sky130_fd_sc_hd__clkbuf_1 _527_ (.A(_189_),
    .X(_016_));
 sky130_fd_sc_hd__and2_1 _528_ (.A(net32),
    .B(_175_),
    .X(_190_));
 sky130_fd_sc_hd__clkbuf_1 _529_ (.A(_190_),
    .X(_017_));
 sky130_fd_sc_hd__buf_2 _530_ (.A(_127_),
    .X(_191_));
 sky130_fd_sc_hd__and2_1 _531_ (.A(net109),
    .B(_191_),
    .X(_192_));
 sky130_fd_sc_hd__clkbuf_1 _532_ (.A(_192_),
    .X(_018_));
 sky130_fd_sc_hd__or4_1 _533_ (.A(\debounce1_a.button_hist[1] ),
    .B(\debounce1_a.button_hist[0] ),
    .C(\debounce1_a.button_hist[3] ),
    .D(\debounce1_a.button_hist[2] ),
    .X(_193_));
 sky130_fd_sc_hd__o41a_1 _534_ (.A1(\debounce1_a.button_hist[4] ),
    .A2(\debounce1_a.button_hist[7] ),
    .A3(\debounce1_a.button_hist[6] ),
    .A4(_193_),
    .B1(\debounce1_a.debounced ),
    .X(_194_));
 sky130_fd_sc_hd__and4_1 _535_ (.A(\debounce1_a.button_hist[1] ),
    .B(\debounce1_a.button_hist[0] ),
    .C(\debounce1_a.button_hist[3] ),
    .D(\debounce1_a.button_hist[2] ),
    .X(_195_));
 sky130_fd_sc_hd__a41o_1 _536_ (.A1(\debounce1_a.button_hist[4] ),
    .A2(\debounce1_a.button_hist[7] ),
    .A3(\debounce1_a.button_hist[6] ),
    .A4(_195_),
    .B1(\debounce1_a.debounced ),
    .X(_196_));
 sky130_fd_sc_hd__o211a_1 _537_ (.A1(net30),
    .A2(_194_),
    .B1(_196_),
    .C1(_169_),
    .X(_019_));
 sky130_fd_sc_hd__and2_1 _538_ (.A(_170_),
    .B(net3),
    .X(_197_));
 sky130_fd_sc_hd__clkbuf_1 _539_ (.A(_197_),
    .X(_020_));
 sky130_fd_sc_hd__and2_1 _540_ (.A(net94),
    .B(_191_),
    .X(_198_));
 sky130_fd_sc_hd__clkbuf_1 _541_ (.A(_198_),
    .X(_021_));
 sky130_fd_sc_hd__and2_1 _542_ (.A(net91),
    .B(_191_),
    .X(_199_));
 sky130_fd_sc_hd__clkbuf_1 _543_ (.A(_199_),
    .X(_022_));
 sky130_fd_sc_hd__and2_1 _544_ (.A(net95),
    .B(_191_),
    .X(_200_));
 sky130_fd_sc_hd__clkbuf_1 _545_ (.A(_200_),
    .X(_023_));
 sky130_fd_sc_hd__and2_1 _546_ (.A(net92),
    .B(_191_),
    .X(_201_));
 sky130_fd_sc_hd__clkbuf_1 _547_ (.A(_201_),
    .X(_024_));
 sky130_fd_sc_hd__and2_1 _548_ (.A(net116),
    .B(_191_),
    .X(_202_));
 sky130_fd_sc_hd__clkbuf_1 _549_ (.A(_202_),
    .X(_025_));
 sky130_fd_sc_hd__and2_1 _550_ (.A(net30),
    .B(_191_),
    .X(_203_));
 sky130_fd_sc_hd__clkbuf_1 _551_ (.A(_203_),
    .X(_026_));
 sky130_fd_sc_hd__and2_1 _552_ (.A(net126),
    .B(_191_),
    .X(_204_));
 sky130_fd_sc_hd__clkbuf_1 _553_ (.A(_204_),
    .X(_027_));
 sky130_fd_sc_hd__or4_1 _554_ (.A(\debounce1_b.button_hist[1] ),
    .B(\debounce1_b.button_hist[0] ),
    .C(\debounce1_b.button_hist[3] ),
    .D(\debounce1_b.button_hist[2] ),
    .X(_205_));
 sky130_fd_sc_hd__o41a_1 _555_ (.A1(\debounce1_b.button_hist[4] ),
    .A2(\debounce1_b.button_hist[7] ),
    .A3(\debounce1_b.button_hist[6] ),
    .A4(_205_),
    .B1(\debounce1_b.debounced ),
    .X(_206_));
 sky130_fd_sc_hd__and4_1 _556_ (.A(\debounce1_b.button_hist[1] ),
    .B(\debounce1_b.button_hist[0] ),
    .C(\debounce1_b.button_hist[3] ),
    .D(\debounce1_b.button_hist[2] ),
    .X(_207_));
 sky130_fd_sc_hd__a41o_1 _557_ (.A1(\debounce1_b.button_hist[4] ),
    .A2(\debounce1_b.button_hist[7] ),
    .A3(\debounce1_b.button_hist[6] ),
    .A4(_207_),
    .B1(\debounce1_b.debounced ),
    .X(_208_));
 sky130_fd_sc_hd__o211a_1 _558_ (.A1(net38),
    .A2(_206_),
    .B1(_208_),
    .C1(_169_),
    .X(_028_));
 sky130_fd_sc_hd__and2_1 _559_ (.A(_170_),
    .B(net4),
    .X(_209_));
 sky130_fd_sc_hd__clkbuf_1 _560_ (.A(_209_),
    .X(_029_));
 sky130_fd_sc_hd__and2_1 _561_ (.A(net111),
    .B(_191_),
    .X(_210_));
 sky130_fd_sc_hd__clkbuf_1 _562_ (.A(_210_),
    .X(_030_));
 sky130_fd_sc_hd__and2_1 _563_ (.A(net86),
    .B(_191_),
    .X(_211_));
 sky130_fd_sc_hd__clkbuf_1 _564_ (.A(_211_),
    .X(_031_));
 sky130_fd_sc_hd__buf_2 _565_ (.A(_127_),
    .X(_212_));
 sky130_fd_sc_hd__and2_1 _566_ (.A(net98),
    .B(_212_),
    .X(_213_));
 sky130_fd_sc_hd__clkbuf_1 _567_ (.A(_213_),
    .X(_032_));
 sky130_fd_sc_hd__and2_1 _568_ (.A(net96),
    .B(_212_),
    .X(_214_));
 sky130_fd_sc_hd__clkbuf_1 _569_ (.A(_214_),
    .X(_033_));
 sky130_fd_sc_hd__and2_1 _570_ (.A(net113),
    .B(_212_),
    .X(_215_));
 sky130_fd_sc_hd__clkbuf_1 _571_ (.A(_215_),
    .X(_034_));
 sky130_fd_sc_hd__and2_1 _572_ (.A(net38),
    .B(_212_),
    .X(_216_));
 sky130_fd_sc_hd__clkbuf_1 _573_ (.A(_216_),
    .X(_035_));
 sky130_fd_sc_hd__and2_1 _574_ (.A(net123),
    .B(_212_),
    .X(_217_));
 sky130_fd_sc_hd__clkbuf_1 _575_ (.A(_217_),
    .X(_036_));
 sky130_fd_sc_hd__or4_1 _576_ (.A(\debounce2_a.button_hist[1] ),
    .B(\debounce2_a.button_hist[0] ),
    .C(\debounce2_a.button_hist[3] ),
    .D(\debounce2_a.button_hist[2] ),
    .X(_218_));
 sky130_fd_sc_hd__o41a_1 _577_ (.A1(\debounce2_a.button_hist[4] ),
    .A2(\debounce2_a.button_hist[7] ),
    .A3(\debounce2_a.button_hist[6] ),
    .A4(_218_),
    .B1(\debounce2_a.debounced ),
    .X(_219_));
 sky130_fd_sc_hd__and4_1 _578_ (.A(\debounce2_a.button_hist[1] ),
    .B(\debounce2_a.button_hist[0] ),
    .C(\debounce2_a.button_hist[3] ),
    .D(\debounce2_a.button_hist[2] ),
    .X(_220_));
 sky130_fd_sc_hd__a41o_1 _579_ (.A1(\debounce2_a.button_hist[4] ),
    .A2(\debounce2_a.button_hist[7] ),
    .A3(\debounce2_a.button_hist[6] ),
    .A4(_220_),
    .B1(\debounce2_a.debounced ),
    .X(_221_));
 sky130_fd_sc_hd__o211a_1 _580_ (.A1(net42),
    .A2(_219_),
    .B1(_221_),
    .C1(_169_),
    .X(_037_));
 sky130_fd_sc_hd__and2_1 _581_ (.A(_170_),
    .B(net5),
    .X(_222_));
 sky130_fd_sc_hd__clkbuf_1 _582_ (.A(_222_),
    .X(_038_));
 sky130_fd_sc_hd__and2_1 _583_ (.A(net106),
    .B(_212_),
    .X(_223_));
 sky130_fd_sc_hd__clkbuf_1 _584_ (.A(_223_),
    .X(_039_));
 sky130_fd_sc_hd__and2_1 _585_ (.A(net103),
    .B(_212_),
    .X(_224_));
 sky130_fd_sc_hd__clkbuf_1 _586_ (.A(_224_),
    .X(_040_));
 sky130_fd_sc_hd__and2_1 _587_ (.A(net93),
    .B(_212_),
    .X(_225_));
 sky130_fd_sc_hd__clkbuf_1 _588_ (.A(_225_),
    .X(_041_));
 sky130_fd_sc_hd__and2_1 _589_ (.A(net88),
    .B(_212_),
    .X(_226_));
 sky130_fd_sc_hd__clkbuf_1 _590_ (.A(_226_),
    .X(_042_));
 sky130_fd_sc_hd__and2_1 _591_ (.A(net122),
    .B(_212_),
    .X(_227_));
 sky130_fd_sc_hd__clkbuf_1 _592_ (.A(_227_),
    .X(_043_));
 sky130_fd_sc_hd__clkbuf_2 _593_ (.A(_127_),
    .X(_228_));
 sky130_fd_sc_hd__and2_1 _594_ (.A(net42),
    .B(_228_),
    .X(_229_));
 sky130_fd_sc_hd__clkbuf_1 _595_ (.A(_229_),
    .X(_044_));
 sky130_fd_sc_hd__and2_1 _596_ (.A(net83),
    .B(_228_),
    .X(_230_));
 sky130_fd_sc_hd__clkbuf_1 _597_ (.A(_230_),
    .X(_045_));
 sky130_fd_sc_hd__or4_1 _598_ (.A(\debounce2_b.button_hist[1] ),
    .B(\debounce2_b.button_hist[0] ),
    .C(\debounce2_b.button_hist[3] ),
    .D(\debounce2_b.button_hist[2] ),
    .X(_231_));
 sky130_fd_sc_hd__o41a_1 _599_ (.A1(\debounce2_b.button_hist[4] ),
    .A2(\debounce2_b.button_hist[7] ),
    .A3(\debounce2_b.button_hist[6] ),
    .A4(_231_),
    .B1(\debounce2_b.debounced ),
    .X(_232_));
 sky130_fd_sc_hd__and4_1 _600_ (.A(\debounce2_b.button_hist[1] ),
    .B(\debounce2_b.button_hist[0] ),
    .C(\debounce2_b.button_hist[3] ),
    .D(\debounce2_b.button_hist[2] ),
    .X(_233_));
 sky130_fd_sc_hd__a41o_1 _601_ (.A1(\debounce2_b.button_hist[4] ),
    .A2(\debounce2_b.button_hist[7] ),
    .A3(\debounce2_b.button_hist[6] ),
    .A4(_233_),
    .B1(\debounce2_b.debounced ),
    .X(_234_));
 sky130_fd_sc_hd__o211a_1 _602_ (.A1(net34),
    .A2(_232_),
    .B1(_234_),
    .C1(_169_),
    .X(_046_));
 sky130_fd_sc_hd__nor2_1 _603_ (.A(_147_),
    .B(net28),
    .Y(_047_));
 sky130_fd_sc_hd__clkbuf_4 _604_ (.A(_128_),
    .X(_235_));
 sky130_fd_sc_hd__o21ai_1 _605_ (.A1(net60),
    .A2(net28),
    .B1(_235_),
    .Y(_236_));
 sky130_fd_sc_hd__a21oi_1 _606_ (.A1(net60),
    .A2(net28),
    .B1(_236_),
    .Y(_048_));
 sky130_fd_sc_hd__and3_1 _607_ (.A(net64),
    .B(net60),
    .C(net28),
    .X(_237_));
 sky130_fd_sc_hd__a21oi_1 _608_ (.A1(net60),
    .A2(net28),
    .B1(net64),
    .Y(_238_));
 sky130_fd_sc_hd__nor3_1 _609_ (.A(_147_),
    .B(_237_),
    .C(_238_),
    .Y(_049_));
 sky130_fd_sc_hd__and2_1 _610_ (.A(net85),
    .B(_237_),
    .X(_239_));
 sky130_fd_sc_hd__o21ai_1 _611_ (.A1(net85),
    .A2(_237_),
    .B1(_235_),
    .Y(_240_));
 sky130_fd_sc_hd__nor2_1 _612_ (.A(_239_),
    .B(_240_),
    .Y(_050_));
 sky130_fd_sc_hd__clkbuf_4 _613_ (.A(_126_),
    .X(_241_));
 sky130_fd_sc_hd__and3_1 _614_ (.A(net50),
    .B(\pwm2.count[3] ),
    .C(_237_),
    .X(_242_));
 sky130_fd_sc_hd__nor2_1 _615_ (.A(_241_),
    .B(_242_),
    .Y(_243_));
 sky130_fd_sc_hd__o21a_1 _616_ (.A1(net50),
    .A2(_239_),
    .B1(_243_),
    .X(_051_));
 sky130_fd_sc_hd__and2_1 _617_ (.A(net71),
    .B(_242_),
    .X(_244_));
 sky130_fd_sc_hd__nor2_1 _618_ (.A(_241_),
    .B(_244_),
    .Y(_245_));
 sky130_fd_sc_hd__o21a_1 _619_ (.A1(net71),
    .A2(_242_),
    .B1(_245_),
    .X(_052_));
 sky130_fd_sc_hd__and3_1 _620_ (.A(net52),
    .B(net71),
    .C(_242_),
    .X(_246_));
 sky130_fd_sc_hd__nor2_1 _621_ (.A(_241_),
    .B(_246_),
    .Y(_247_));
 sky130_fd_sc_hd__o21a_1 _622_ (.A1(net52),
    .A2(_244_),
    .B1(_247_),
    .X(_053_));
 sky130_fd_sc_hd__a21oi_1 _623_ (.A1(net75),
    .A2(_246_),
    .B1(_241_),
    .Y(_248_));
 sky130_fd_sc_hd__o21a_1 _624_ (.A1(net75),
    .A2(_246_),
    .B1(_248_),
    .X(_054_));
 sky130_fd_sc_hd__and2_1 _625_ (.A(net155),
    .B(_228_),
    .X(_249_));
 sky130_fd_sc_hd__clkbuf_1 _626_ (.A(_249_),
    .X(_055_));
 sky130_fd_sc_hd__and2_1 _627_ (.A(_170_),
    .B(net6),
    .X(_250_));
 sky130_fd_sc_hd__clkbuf_1 _628_ (.A(_250_),
    .X(_056_));
 sky130_fd_sc_hd__and2_1 _629_ (.A(net84),
    .B(_228_),
    .X(_251_));
 sky130_fd_sc_hd__clkbuf_1 _630_ (.A(_251_),
    .X(_057_));
 sky130_fd_sc_hd__and2_1 _631_ (.A(net87),
    .B(_228_),
    .X(_252_));
 sky130_fd_sc_hd__clkbuf_1 _632_ (.A(_252_),
    .X(_058_));
 sky130_fd_sc_hd__and2_1 _633_ (.A(net80),
    .B(_228_),
    .X(_253_));
 sky130_fd_sc_hd__clkbuf_1 _634_ (.A(_253_),
    .X(_059_));
 sky130_fd_sc_hd__and2_1 _635_ (.A(net79),
    .B(_228_),
    .X(_254_));
 sky130_fd_sc_hd__clkbuf_1 _636_ (.A(_254_),
    .X(_060_));
 sky130_fd_sc_hd__and2_1 _637_ (.A(net78),
    .B(_228_),
    .X(_255_));
 sky130_fd_sc_hd__clkbuf_1 _638_ (.A(_255_),
    .X(_061_));
 sky130_fd_sc_hd__and2_1 _639_ (.A(net34),
    .B(_228_),
    .X(_256_));
 sky130_fd_sc_hd__clkbuf_1 _640_ (.A(_256_),
    .X(_062_));
 sky130_fd_sc_hd__and2_1 _641_ (.A(net112),
    .B(_228_),
    .X(_257_));
 sky130_fd_sc_hd__clkbuf_1 _642_ (.A(_257_),
    .X(_063_));
 sky130_fd_sc_hd__and2b_1 _643_ (.A_N(net155),
    .B(net163),
    .X(_258_));
 sky130_fd_sc_hd__and2b_1 _644_ (.A_N(net163),
    .B(net155),
    .X(_259_));
 sky130_fd_sc_hd__and2_1 _645_ (.A(\encoder0.old_b ),
    .B(\encoder0.old_a ),
    .X(_260_));
 sky130_fd_sc_hd__nor2_1 _646_ (.A(\encoder0.old_b ),
    .B(\encoder0.old_a ),
    .Y(_261_));
 sky130_fd_sc_hd__o22a_2 _647_ (.A1(_258_),
    .A2(_259_),
    .B1(_260_),
    .B2(_261_),
    .X(_262_));
 sky130_fd_sc_hd__clkbuf_4 _648_ (.A(_262_),
    .X(_263_));
 sky130_fd_sc_hd__a21oi_1 _649_ (.A1(net129),
    .A2(_262_),
    .B1(_241_),
    .Y(_264_));
 sky130_fd_sc_hd__o21a_1 _650_ (.A1(net129),
    .A2(_263_),
    .B1(_264_),
    .X(_064_));
 sky130_fd_sc_hd__o22a_1 _651_ (.A1(_258_),
    .A2(_260_),
    .B1(_261_),
    .B2(_259_),
    .X(_265_));
 sky130_fd_sc_hd__or2_1 _652_ (.A(net101),
    .B(_265_),
    .X(_266_));
 sky130_fd_sc_hd__nand2_1 _653_ (.A(net101),
    .B(_265_),
    .Y(_267_));
 sky130_fd_sc_hd__a21oi_1 _654_ (.A1(_266_),
    .A2(_267_),
    .B1(\encoder0.value[0] ),
    .Y(_268_));
 sky130_fd_sc_hd__and3_1 _655_ (.A(\encoder0.value[0] ),
    .B(_266_),
    .C(_267_),
    .X(_269_));
 sky130_fd_sc_hd__o21ai_1 _656_ (.A1(_268_),
    .A2(_269_),
    .B1(_263_),
    .Y(_270_));
 sky130_fd_sc_hd__o211a_1 _657_ (.A1(net101),
    .A2(_263_),
    .B1(_270_),
    .C1(_169_),
    .X(_065_));
 sky130_fd_sc_hd__a21boi_2 _658_ (.A1(net129),
    .A2(_266_),
    .B1_N(_267_),
    .Y(_271_));
 sky130_fd_sc_hd__or2_1 _659_ (.A(net141),
    .B(_265_),
    .X(_272_));
 sky130_fd_sc_hd__clkbuf_4 _660_ (.A(_265_),
    .X(_273_));
 sky130_fd_sc_hd__nand2_1 _661_ (.A(net141),
    .B(_273_),
    .Y(_274_));
 sky130_fd_sc_hd__nand2_1 _662_ (.A(_272_),
    .B(_274_),
    .Y(_275_));
 sky130_fd_sc_hd__xnor2_1 _663_ (.A(_271_),
    .B(_275_),
    .Y(_276_));
 sky130_fd_sc_hd__nand2_1 _664_ (.A(_263_),
    .B(_276_),
    .Y(_277_));
 sky130_fd_sc_hd__o211a_1 _665_ (.A1(net141),
    .A2(_263_),
    .B1(_277_),
    .C1(_169_),
    .X(_066_));
 sky130_fd_sc_hd__xnor2_1 _666_ (.A(net143),
    .B(_273_),
    .Y(_278_));
 sky130_fd_sc_hd__o21ai_1 _667_ (.A1(_271_),
    .A2(_275_),
    .B1(_274_),
    .Y(_279_));
 sky130_fd_sc_hd__o21ai_1 _668_ (.A1(_278_),
    .A2(_279_),
    .B1(_262_),
    .Y(_280_));
 sky130_fd_sc_hd__a21o_1 _669_ (.A1(_278_),
    .A2(_279_),
    .B1(_280_),
    .X(_281_));
 sky130_fd_sc_hd__o211a_1 _670_ (.A1(net143),
    .A2(_263_),
    .B1(_281_),
    .C1(_169_),
    .X(_067_));
 sky130_fd_sc_hd__o21ai_1 _671_ (.A1(net143),
    .A2(net141),
    .B1(_273_),
    .Y(_282_));
 sky130_fd_sc_hd__o31a_1 _672_ (.A1(_271_),
    .A2(_275_),
    .A3(_278_),
    .B1(_282_),
    .X(_283_));
 sky130_fd_sc_hd__xnor2_1 _673_ (.A(net165),
    .B(_273_),
    .Y(_284_));
 sky130_fd_sc_hd__and2_1 _674_ (.A(_283_),
    .B(_284_),
    .X(_285_));
 sky130_fd_sc_hd__nor2_1 _675_ (.A(_283_),
    .B(_284_),
    .Y(_286_));
 sky130_fd_sc_hd__o21ai_1 _676_ (.A1(_285_),
    .A2(_286_),
    .B1(_263_),
    .Y(_287_));
 sky130_fd_sc_hd__o211a_1 _677_ (.A1(net165),
    .A2(_263_),
    .B1(_287_),
    .C1(_169_),
    .X(_068_));
 sky130_fd_sc_hd__xnor2_1 _678_ (.A(net161),
    .B(_273_),
    .Y(_288_));
 sky130_fd_sc_hd__a21o_1 _679_ (.A1(\encoder0.value[4] ),
    .A2(_273_),
    .B1(_286_),
    .X(_289_));
 sky130_fd_sc_hd__nor2_1 _680_ (.A(_288_),
    .B(_289_),
    .Y(_290_));
 sky130_fd_sc_hd__a21bo_1 _681_ (.A1(_288_),
    .A2(_289_),
    .B1_N(_262_),
    .X(_291_));
 sky130_fd_sc_hd__o221a_1 _682_ (.A1(net161),
    .A2(_263_),
    .B1(_290_),
    .B2(_291_),
    .C1(_129_),
    .X(_069_));
 sky130_fd_sc_hd__inv_2 _683_ (.A(net169),
    .Y(_292_));
 sky130_fd_sc_hd__nor2_1 _684_ (.A(net169),
    .B(_273_),
    .Y(_293_));
 sky130_fd_sc_hd__and2_1 _685_ (.A(\encoder0.value[6] ),
    .B(_273_),
    .X(_294_));
 sky130_fd_sc_hd__or2_1 _686_ (.A(_293_),
    .B(_294_),
    .X(_295_));
 sky130_fd_sc_hd__o21ai_1 _687_ (.A1(net161),
    .A2(net165),
    .B1(_273_),
    .Y(_296_));
 sky130_fd_sc_hd__o31a_1 _688_ (.A1(_283_),
    .A2(_284_),
    .A3(_288_),
    .B1(_296_),
    .X(_297_));
 sky130_fd_sc_hd__nor2_1 _689_ (.A(_295_),
    .B(_297_),
    .Y(_298_));
 sky130_fd_sc_hd__a21bo_1 _690_ (.A1(_295_),
    .A2(_297_),
    .B1_N(_262_),
    .X(_299_));
 sky130_fd_sc_hd__o22ai_1 _691_ (.A1(_292_),
    .A2(_262_),
    .B1(_298_),
    .B2(_299_),
    .Y(_300_));
 sky130_fd_sc_hd__and2_1 _692_ (.A(_170_),
    .B(net170),
    .X(_301_));
 sky130_fd_sc_hd__clkbuf_1 _693_ (.A(_301_),
    .X(_070_));
 sky130_fd_sc_hd__xnor2_1 _694_ (.A(net124),
    .B(_273_),
    .Y(_302_));
 sky130_fd_sc_hd__o21a_1 _695_ (.A1(_294_),
    .A2(_298_),
    .B1(_302_),
    .X(_303_));
 sky130_fd_sc_hd__o31ai_1 _696_ (.A1(_294_),
    .A2(_298_),
    .A3(_302_),
    .B1(_262_),
    .Y(_304_));
 sky130_fd_sc_hd__o221a_1 _697_ (.A1(net124),
    .A2(_263_),
    .B1(_303_),
    .B2(_304_),
    .C1(_235_),
    .X(_071_));
 sky130_fd_sc_hd__and2_1 _698_ (.A(net164),
    .B(_128_),
    .X(_305_));
 sky130_fd_sc_hd__clkbuf_1 _699_ (.A(_305_),
    .X(_072_));
 sky130_fd_sc_hd__and2_1 _700_ (.A(net163),
    .B(_128_),
    .X(_306_));
 sky130_fd_sc_hd__clkbuf_1 _701_ (.A(_306_),
    .X(_073_));
 sky130_fd_sc_hd__and2b_1 _702_ (.A_N(\debounce1_a.debounced ),
    .B(\debounce1_b.debounced ),
    .X(_307_));
 sky130_fd_sc_hd__and2b_1 _703_ (.A_N(\debounce1_b.debounced ),
    .B(\debounce1_a.debounced ),
    .X(_308_));
 sky130_fd_sc_hd__and2_1 _704_ (.A(\encoder1.old_b ),
    .B(\encoder1.old_a ),
    .X(_309_));
 sky130_fd_sc_hd__nor2_1 _705_ (.A(\encoder1.old_b ),
    .B(\encoder1.old_a ),
    .Y(_310_));
 sky130_fd_sc_hd__o22a_2 _706_ (.A1(_307_),
    .A2(_308_),
    .B1(_309_),
    .B2(_310_),
    .X(_311_));
 sky130_fd_sc_hd__buf_2 _707_ (.A(_311_),
    .X(_312_));
 sky130_fd_sc_hd__a21oi_1 _708_ (.A1(net151),
    .A2(_311_),
    .B1(_241_),
    .Y(_313_));
 sky130_fd_sc_hd__o21a_1 _709_ (.A1(net151),
    .A2(_312_),
    .B1(_313_),
    .X(_074_));
 sky130_fd_sc_hd__o22a_1 _710_ (.A1(_307_),
    .A2(_309_),
    .B1(_310_),
    .B2(_308_),
    .X(_314_));
 sky130_fd_sc_hd__or2_1 _711_ (.A(net107),
    .B(_314_),
    .X(_315_));
 sky130_fd_sc_hd__nand2_1 _712_ (.A(net107),
    .B(_314_),
    .Y(_316_));
 sky130_fd_sc_hd__a21oi_1 _713_ (.A1(_315_),
    .A2(_316_),
    .B1(\encoder1.value[0] ),
    .Y(_317_));
 sky130_fd_sc_hd__and3_1 _714_ (.A(\encoder1.value[0] ),
    .B(_315_),
    .C(_316_),
    .X(_318_));
 sky130_fd_sc_hd__o21ai_1 _715_ (.A1(_317_),
    .A2(_318_),
    .B1(_312_),
    .Y(_319_));
 sky130_fd_sc_hd__o211a_1 _716_ (.A1(net107),
    .A2(_312_),
    .B1(_319_),
    .C1(_129_),
    .X(_075_));
 sky130_fd_sc_hd__a21boi_2 _717_ (.A1(\encoder1.value[0] ),
    .A2(_315_),
    .B1_N(_316_),
    .Y(_320_));
 sky130_fd_sc_hd__or2_1 _718_ (.A(net131),
    .B(_314_),
    .X(_321_));
 sky130_fd_sc_hd__clkbuf_4 _719_ (.A(_314_),
    .X(_322_));
 sky130_fd_sc_hd__nand2_1 _720_ (.A(net131),
    .B(_322_),
    .Y(_323_));
 sky130_fd_sc_hd__nand2_1 _721_ (.A(_321_),
    .B(_323_),
    .Y(_324_));
 sky130_fd_sc_hd__xnor2_1 _722_ (.A(_320_),
    .B(_324_),
    .Y(_325_));
 sky130_fd_sc_hd__nand2_1 _723_ (.A(_312_),
    .B(_325_),
    .Y(_326_));
 sky130_fd_sc_hd__o211a_1 _724_ (.A1(net131),
    .A2(_312_),
    .B1(_326_),
    .C1(_129_),
    .X(_076_));
 sky130_fd_sc_hd__xnor2_1 _725_ (.A(net145),
    .B(_322_),
    .Y(_327_));
 sky130_fd_sc_hd__o21ai_1 _726_ (.A1(_320_),
    .A2(_324_),
    .B1(_323_),
    .Y(_328_));
 sky130_fd_sc_hd__o21ai_1 _727_ (.A1(_327_),
    .A2(_328_),
    .B1(_311_),
    .Y(_329_));
 sky130_fd_sc_hd__a21o_1 _728_ (.A1(_327_),
    .A2(_328_),
    .B1(_329_),
    .X(_330_));
 sky130_fd_sc_hd__o211a_1 _729_ (.A1(net145),
    .A2(_312_),
    .B1(_330_),
    .C1(_129_),
    .X(_077_));
 sky130_fd_sc_hd__o21ai_1 _730_ (.A1(net145),
    .A2(net131),
    .B1(_322_),
    .Y(_331_));
 sky130_fd_sc_hd__o31a_1 _731_ (.A1(_320_),
    .A2(_324_),
    .A3(_327_),
    .B1(_331_),
    .X(_332_));
 sky130_fd_sc_hd__nor2_1 _732_ (.A(net133),
    .B(_322_),
    .Y(_333_));
 sky130_fd_sc_hd__and2_1 _733_ (.A(net133),
    .B(_322_),
    .X(_334_));
 sky130_fd_sc_hd__or2_1 _734_ (.A(_333_),
    .B(_334_),
    .X(_335_));
 sky130_fd_sc_hd__and2_1 _735_ (.A(_332_),
    .B(_335_),
    .X(_336_));
 sky130_fd_sc_hd__nor2_1 _736_ (.A(_332_),
    .B(_335_),
    .Y(_337_));
 sky130_fd_sc_hd__o21ai_1 _737_ (.A1(_336_),
    .A2(_337_),
    .B1(_312_),
    .Y(_338_));
 sky130_fd_sc_hd__o211a_1 _738_ (.A1(net133),
    .A2(_312_),
    .B1(_338_),
    .C1(_129_),
    .X(_078_));
 sky130_fd_sc_hd__xnor2_1 _739_ (.A(net149),
    .B(_322_),
    .Y(_339_));
 sky130_fd_sc_hd__o21a_1 _740_ (.A1(_334_),
    .A2(_337_),
    .B1(_339_),
    .X(_340_));
 sky130_fd_sc_hd__o31ai_1 _741_ (.A1(_334_),
    .A2(_337_),
    .A3(_339_),
    .B1(_311_),
    .Y(_341_));
 sky130_fd_sc_hd__o221a_1 _742_ (.A1(net149),
    .A2(_312_),
    .B1(_340_),
    .B2(_341_),
    .C1(_235_),
    .X(_079_));
 sky130_fd_sc_hd__nor2_1 _743_ (.A(net153),
    .B(_322_),
    .Y(_342_));
 sky130_fd_sc_hd__and2_1 _744_ (.A(net153),
    .B(_322_),
    .X(_343_));
 sky130_fd_sc_hd__or2_1 _745_ (.A(_342_),
    .B(_343_),
    .X(_344_));
 sky130_fd_sc_hd__o21ai_1 _746_ (.A1(net149),
    .A2(net133),
    .B1(_322_),
    .Y(_345_));
 sky130_fd_sc_hd__o31a_1 _747_ (.A1(_332_),
    .A2(_335_),
    .A3(_339_),
    .B1(_345_),
    .X(_346_));
 sky130_fd_sc_hd__nor2_1 _748_ (.A(_344_),
    .B(_346_),
    .Y(_347_));
 sky130_fd_sc_hd__a21bo_1 _749_ (.A1(_344_),
    .A2(_346_),
    .B1_N(_311_),
    .X(_348_));
 sky130_fd_sc_hd__o22a_1 _750_ (.A1(_131_),
    .A2(_311_),
    .B1(_347_),
    .B2(_348_),
    .X(_349_));
 sky130_fd_sc_hd__nor2_1 _751_ (.A(_147_),
    .B(net154),
    .Y(_080_));
 sky130_fd_sc_hd__xnor2_1 _752_ (.A(net119),
    .B(_322_),
    .Y(_350_));
 sky130_fd_sc_hd__o21a_1 _753_ (.A1(_343_),
    .A2(_347_),
    .B1(_350_),
    .X(_351_));
 sky130_fd_sc_hd__o31ai_1 _754_ (.A1(_343_),
    .A2(_347_),
    .A3(_350_),
    .B1(_311_),
    .Y(_352_));
 sky130_fd_sc_hd__o221a_1 _755_ (.A1(net119),
    .A2(_312_),
    .B1(_351_),
    .B2(_352_),
    .C1(_235_),
    .X(_081_));
 sky130_fd_sc_hd__and2_1 _756_ (.A(net167),
    .B(_128_),
    .X(_353_));
 sky130_fd_sc_hd__clkbuf_1 _757_ (.A(_353_),
    .X(_082_));
 sky130_fd_sc_hd__and2_1 _758_ (.A(net168),
    .B(_128_),
    .X(_354_));
 sky130_fd_sc_hd__clkbuf_1 _759_ (.A(_354_),
    .X(_083_));
 sky130_fd_sc_hd__and2b_1 _760_ (.A_N(\debounce2_a.debounced ),
    .B(net156),
    .X(_355_));
 sky130_fd_sc_hd__and2b_1 _761_ (.A_N(net156),
    .B(\debounce2_a.debounced ),
    .X(_356_));
 sky130_fd_sc_hd__and2_1 _762_ (.A(\encoder2.old_b ),
    .B(\encoder2.old_a ),
    .X(_357_));
 sky130_fd_sc_hd__nor2_1 _763_ (.A(\encoder2.old_b ),
    .B(\encoder2.old_a ),
    .Y(_358_));
 sky130_fd_sc_hd__o22a_2 _764_ (.A1(_355_),
    .A2(_356_),
    .B1(_357_),
    .B2(_358_),
    .X(_359_));
 sky130_fd_sc_hd__buf_2 _765_ (.A(_359_),
    .X(_360_));
 sky130_fd_sc_hd__a21oi_1 _766_ (.A1(net147),
    .A2(_359_),
    .B1(_241_),
    .Y(_361_));
 sky130_fd_sc_hd__o21a_1 _767_ (.A1(net147),
    .A2(_360_),
    .B1(_361_),
    .X(_084_));
 sky130_fd_sc_hd__o22a_1 _768_ (.A1(_355_),
    .A2(_357_),
    .B1(_358_),
    .B2(_356_),
    .X(_362_));
 sky130_fd_sc_hd__or2_1 _769_ (.A(net104),
    .B(_362_),
    .X(_363_));
 sky130_fd_sc_hd__nand2_1 _770_ (.A(net104),
    .B(_362_),
    .Y(_364_));
 sky130_fd_sc_hd__a21oi_1 _771_ (.A1(_363_),
    .A2(_364_),
    .B1(\encoder2.value[0] ),
    .Y(_365_));
 sky130_fd_sc_hd__and3_1 _772_ (.A(\encoder2.value[0] ),
    .B(_363_),
    .C(_364_),
    .X(_366_));
 sky130_fd_sc_hd__o21ai_1 _773_ (.A1(_365_),
    .A2(_366_),
    .B1(_360_),
    .Y(_367_));
 sky130_fd_sc_hd__o211a_1 _774_ (.A1(net104),
    .A2(_360_),
    .B1(_367_),
    .C1(_129_),
    .X(_085_));
 sky130_fd_sc_hd__a21boi_2 _775_ (.A1(\encoder2.value[0] ),
    .A2(_363_),
    .B1_N(_364_),
    .Y(_368_));
 sky130_fd_sc_hd__or2_1 _776_ (.A(net135),
    .B(_362_),
    .X(_369_));
 sky130_fd_sc_hd__clkbuf_4 _777_ (.A(_362_),
    .X(_370_));
 sky130_fd_sc_hd__nand2_1 _778_ (.A(net135),
    .B(_370_),
    .Y(_371_));
 sky130_fd_sc_hd__nand2_1 _779_ (.A(_369_),
    .B(_371_),
    .Y(_372_));
 sky130_fd_sc_hd__xnor2_1 _780_ (.A(_368_),
    .B(_372_),
    .Y(_373_));
 sky130_fd_sc_hd__nand2_1 _781_ (.A(_360_),
    .B(_373_),
    .Y(_374_));
 sky130_fd_sc_hd__o211a_1 _782_ (.A1(net135),
    .A2(_360_),
    .B1(_374_),
    .C1(_129_),
    .X(_086_));
 sky130_fd_sc_hd__xnor2_1 _783_ (.A(net127),
    .B(_370_),
    .Y(_375_));
 sky130_fd_sc_hd__o21ai_1 _784_ (.A1(_368_),
    .A2(_372_),
    .B1(_371_),
    .Y(_376_));
 sky130_fd_sc_hd__o21ai_1 _785_ (.A1(_375_),
    .A2(_376_),
    .B1(_359_),
    .Y(_377_));
 sky130_fd_sc_hd__a21o_1 _786_ (.A1(_375_),
    .A2(_376_),
    .B1(_377_),
    .X(_378_));
 sky130_fd_sc_hd__o211a_1 _787_ (.A1(net127),
    .A2(_360_),
    .B1(_378_),
    .C1(_129_),
    .X(_087_));
 sky130_fd_sc_hd__o21ai_1 _788_ (.A1(net127),
    .A2(net135),
    .B1(_370_),
    .Y(_379_));
 sky130_fd_sc_hd__o31a_1 _789_ (.A1(_368_),
    .A2(_372_),
    .A3(_375_),
    .B1(_379_),
    .X(_380_));
 sky130_fd_sc_hd__nor2_1 _790_ (.A(net139),
    .B(_370_),
    .Y(_381_));
 sky130_fd_sc_hd__and2_1 _791_ (.A(net139),
    .B(_370_),
    .X(_382_));
 sky130_fd_sc_hd__or2_1 _792_ (.A(_381_),
    .B(_382_),
    .X(_383_));
 sky130_fd_sc_hd__and2_1 _793_ (.A(_380_),
    .B(_383_),
    .X(_384_));
 sky130_fd_sc_hd__nor2_1 _794_ (.A(_380_),
    .B(_383_),
    .Y(_385_));
 sky130_fd_sc_hd__o21ai_1 _795_ (.A1(_384_),
    .A2(_385_),
    .B1(_360_),
    .Y(_386_));
 sky130_fd_sc_hd__o211a_1 _796_ (.A1(net139),
    .A2(_360_),
    .B1(_386_),
    .C1(_129_),
    .X(_088_));
 sky130_fd_sc_hd__xnor2_1 _797_ (.A(net157),
    .B(_370_),
    .Y(_387_));
 sky130_fd_sc_hd__o21a_1 _798_ (.A1(_382_),
    .A2(_385_),
    .B1(_387_),
    .X(_388_));
 sky130_fd_sc_hd__o31ai_1 _799_ (.A1(_382_),
    .A2(_385_),
    .A3(_387_),
    .B1(_359_),
    .Y(_389_));
 sky130_fd_sc_hd__o221a_1 _800_ (.A1(net157),
    .A2(_360_),
    .B1(_388_),
    .B2(_389_),
    .C1(_235_),
    .X(_089_));
 sky130_fd_sc_hd__nor2_1 _801_ (.A(net159),
    .B(_370_),
    .Y(_390_));
 sky130_fd_sc_hd__and2_1 _802_ (.A(net159),
    .B(_370_),
    .X(_391_));
 sky130_fd_sc_hd__or2_1 _803_ (.A(_390_),
    .B(_391_),
    .X(_392_));
 sky130_fd_sc_hd__o21ai_1 _804_ (.A1(net157),
    .A2(net139),
    .B1(_370_),
    .Y(_393_));
 sky130_fd_sc_hd__o31a_1 _805_ (.A1(_380_),
    .A2(_383_),
    .A3(_387_),
    .B1(_393_),
    .X(_394_));
 sky130_fd_sc_hd__nor2_1 _806_ (.A(_392_),
    .B(_394_),
    .Y(_395_));
 sky130_fd_sc_hd__a21bo_1 _807_ (.A1(_392_),
    .A2(_394_),
    .B1_N(_359_),
    .X(_396_));
 sky130_fd_sc_hd__o22a_1 _808_ (.A1(_149_),
    .A2(_359_),
    .B1(_395_),
    .B2(_396_),
    .X(_397_));
 sky130_fd_sc_hd__nor2_1 _809_ (.A(_147_),
    .B(net160),
    .Y(_090_));
 sky130_fd_sc_hd__xnor2_1 _810_ (.A(net114),
    .B(_370_),
    .Y(_398_));
 sky130_fd_sc_hd__o21a_1 _811_ (.A1(_391_),
    .A2(_395_),
    .B1(_398_),
    .X(_399_));
 sky130_fd_sc_hd__o31ai_1 _812_ (.A1(_391_),
    .A2(_395_),
    .A3(_398_),
    .B1(_359_),
    .Y(_400_));
 sky130_fd_sc_hd__o221a_1 _813_ (.A1(net114),
    .A2(_360_),
    .B1(_399_),
    .B2(_400_),
    .C1(_235_),
    .X(_091_));
 sky130_fd_sc_hd__and2_1 _814_ (.A(net156),
    .B(_128_),
    .X(_401_));
 sky130_fd_sc_hd__clkbuf_1 _815_ (.A(_401_),
    .X(_092_));
 sky130_fd_sc_hd__nor2_1 _816_ (.A(_147_),
    .B(net26),
    .Y(_093_));
 sky130_fd_sc_hd__a21oi_1 _817_ (.A1(_117_),
    .A2(_119_),
    .B1(_241_),
    .Y(_402_));
 sky130_fd_sc_hd__o21a_1 _818_ (.A1(_117_),
    .A2(_119_),
    .B1(_402_),
    .X(_094_));
 sky130_fd_sc_hd__and3_1 _819_ (.A(net58),
    .B(net54),
    .C(net26),
    .X(_403_));
 sky130_fd_sc_hd__a21oi_1 _820_ (.A1(net54),
    .A2(net26),
    .B1(net58),
    .Y(_404_));
 sky130_fd_sc_hd__nor3_1 _821_ (.A(_147_),
    .B(_403_),
    .C(_404_),
    .Y(_095_));
 sky130_fd_sc_hd__and2_1 _822_ (.A(net99),
    .B(_403_),
    .X(_405_));
 sky130_fd_sc_hd__o21ai_1 _823_ (.A1(net99),
    .A2(_403_),
    .B1(_235_),
    .Y(_406_));
 sky130_fd_sc_hd__nor2_1 _824_ (.A(_405_),
    .B(_406_),
    .Y(_096_));
 sky130_fd_sc_hd__and3_1 _825_ (.A(net46),
    .B(\pwm0.count[3] ),
    .C(_403_),
    .X(_407_));
 sky130_fd_sc_hd__nor2_1 _826_ (.A(_126_),
    .B(_407_),
    .Y(_408_));
 sky130_fd_sc_hd__o21a_1 _827_ (.A1(net46),
    .A2(_405_),
    .B1(_408_),
    .X(_097_));
 sky130_fd_sc_hd__and2_1 _828_ (.A(net69),
    .B(_407_),
    .X(_409_));
 sky130_fd_sc_hd__nor2_1 _829_ (.A(_126_),
    .B(_409_),
    .Y(_410_));
 sky130_fd_sc_hd__o21a_1 _830_ (.A1(net69),
    .A2(_407_),
    .B1(_410_),
    .X(_098_));
 sky130_fd_sc_hd__and3_1 _831_ (.A(net44),
    .B(\pwm0.count[5] ),
    .C(_407_),
    .X(_411_));
 sky130_fd_sc_hd__nor2_1 _832_ (.A(_126_),
    .B(_411_),
    .Y(_412_));
 sky130_fd_sc_hd__o21a_1 _833_ (.A1(net44),
    .A2(_409_),
    .B1(_412_),
    .X(_099_));
 sky130_fd_sc_hd__a21oi_1 _834_ (.A1(net56),
    .A2(_411_),
    .B1(_241_),
    .Y(_413_));
 sky130_fd_sc_hd__o21a_1 _835_ (.A1(net56),
    .A2(_411_),
    .B1(_413_),
    .X(_100_));
 sky130_fd_sc_hd__nor2_1 _836_ (.A(_147_),
    .B(net40),
    .Y(_101_));
 sky130_fd_sc_hd__o21ai_1 _837_ (.A1(net63),
    .A2(net40),
    .B1(_235_),
    .Y(_414_));
 sky130_fd_sc_hd__a21oi_1 _838_ (.A1(net63),
    .A2(net40),
    .B1(_414_),
    .Y(_102_));
 sky130_fd_sc_hd__and3_1 _839_ (.A(net66),
    .B(net63),
    .C(net40),
    .X(_415_));
 sky130_fd_sc_hd__a21oi_1 _840_ (.A1(net63),
    .A2(net40),
    .B1(net66),
    .Y(_416_));
 sky130_fd_sc_hd__nor3_1 _841_ (.A(_147_),
    .B(_415_),
    .C(_416_),
    .Y(_103_));
 sky130_fd_sc_hd__and2_1 _842_ (.A(net81),
    .B(_415_),
    .X(_417_));
 sky130_fd_sc_hd__o21ai_1 _843_ (.A1(net81),
    .A2(_415_),
    .B1(_235_),
    .Y(_418_));
 sky130_fd_sc_hd__nor2_1 _844_ (.A(_417_),
    .B(_418_),
    .Y(_104_));
 sky130_fd_sc_hd__and3_1 _845_ (.A(net61),
    .B(net81),
    .C(_415_),
    .X(_419_));
 sky130_fd_sc_hd__nor2_1 _846_ (.A(_126_),
    .B(_419_),
    .Y(_420_));
 sky130_fd_sc_hd__o21a_1 _847_ (.A1(net61),
    .A2(_417_),
    .B1(_420_),
    .X(_105_));
 sky130_fd_sc_hd__and2_1 _848_ (.A(net73),
    .B(_419_),
    .X(_421_));
 sky130_fd_sc_hd__nor2_1 _849_ (.A(_126_),
    .B(_421_),
    .Y(_422_));
 sky130_fd_sc_hd__o21a_1 _850_ (.A1(net73),
    .A2(_419_),
    .B1(_422_),
    .X(_106_));
 sky130_fd_sc_hd__and3_1 _851_ (.A(net48),
    .B(net73),
    .C(_419_),
    .X(_423_));
 sky130_fd_sc_hd__nor2_1 _852_ (.A(_126_),
    .B(_423_),
    .Y(_424_));
 sky130_fd_sc_hd__o21a_1 _853_ (.A1(net48),
    .A2(_421_),
    .B1(_424_),
    .X(_107_));
 sky130_fd_sc_hd__a21oi_1 _854_ (.A1(net138),
    .A2(_423_),
    .B1(_241_),
    .Y(_425_));
 sky130_fd_sc_hd__o21a_1 _855_ (.A1(net138),
    .A2(_423_),
    .B1(_425_),
    .X(_108_));
 sky130_fd_sc_hd__dfstp_1 _856_ (.CLK(clknet_3_5__leaf_clk),
    .D(net12),
    .SET_B(net25),
    .Q(\debounce0_a.reset ));
 sky130_fd_sc_hd__conb_1 _856__12 (.LO(net12));
 sky130_fd_sc_hd__dfxtp_1 _857_ (.CLK(clknet_3_7__leaf_clk),
    .D(net37),
    .Q(\debounce0_a.debounced ));
 sky130_fd_sc_hd__dfxtp_1 _858_ (.CLK(clknet_3_5__leaf_clk),
    .D(_002_),
    .Q(\debounce0_a.button_hist[0] ));
 sky130_fd_sc_hd__dfxtp_1 _859_ (.CLK(clknet_3_5__leaf_clk),
    .D(_003_),
    .Q(\debounce0_a.button_hist[1] ));
 sky130_fd_sc_hd__dfxtp_1 _860_ (.CLK(clknet_3_5__leaf_clk),
    .D(_004_),
    .Q(\debounce0_a.button_hist[2] ));
 sky130_fd_sc_hd__dfxtp_1 _861_ (.CLK(clknet_3_7__leaf_clk),
    .D(_005_),
    .Q(\debounce0_a.button_hist[3] ));
 sky130_fd_sc_hd__dfxtp_1 _862_ (.CLK(clknet_3_7__leaf_clk),
    .D(_006_),
    .Q(\debounce0_a.button_hist[4] ));
 sky130_fd_sc_hd__dfxtp_1 _863_ (.CLK(clknet_3_7__leaf_clk),
    .D(_007_),
    .Q(\debounce0_a.button_hist[5] ));
 sky130_fd_sc_hd__dfxtp_1 _864_ (.CLK(clknet_3_7__leaf_clk),
    .D(_008_),
    .Q(\debounce0_a.button_hist[6] ));
 sky130_fd_sc_hd__dfxtp_1 _865_ (.CLK(clknet_3_7__leaf_clk),
    .D(_009_),
    .Q(\debounce0_a.button_hist[7] ));
 sky130_fd_sc_hd__dfxtp_1 _866_ (.CLK(clknet_3_7__leaf_clk),
    .D(net33),
    .Q(\debounce0_b.debounced ));
 sky130_fd_sc_hd__dfxtp_1 _867_ (.CLK(clknet_3_7__leaf_clk),
    .D(_011_),
    .Q(\debounce0_b.button_hist[0] ));
 sky130_fd_sc_hd__dfxtp_1 _868_ (.CLK(clknet_3_7__leaf_clk),
    .D(_012_),
    .Q(\debounce0_b.button_hist[1] ));
 sky130_fd_sc_hd__dfxtp_1 _869_ (.CLK(clknet_3_7__leaf_clk),
    .D(_013_),
    .Q(\debounce0_b.button_hist[2] ));
 sky130_fd_sc_hd__dfxtp_1 _870_ (.CLK(clknet_3_7__leaf_clk),
    .D(_014_),
    .Q(\debounce0_b.button_hist[3] ));
 sky130_fd_sc_hd__dfxtp_1 _871_ (.CLK(clknet_3_7__leaf_clk),
    .D(_015_),
    .Q(\debounce0_b.button_hist[4] ));
 sky130_fd_sc_hd__dfxtp_1 _872_ (.CLK(clknet_3_7__leaf_clk),
    .D(_016_),
    .Q(\debounce0_b.button_hist[5] ));
 sky130_fd_sc_hd__dfxtp_1 _873_ (.CLK(clknet_3_7__leaf_clk),
    .D(_017_),
    .Q(\debounce0_b.button_hist[6] ));
 sky130_fd_sc_hd__dfxtp_1 _874_ (.CLK(clknet_3_7__leaf_clk),
    .D(_018_),
    .Q(\debounce0_b.button_hist[7] ));
 sky130_fd_sc_hd__dfxtp_1 _875_ (.CLK(clknet_3_6__leaf_clk),
    .D(net31),
    .Q(\debounce1_a.debounced ));
 sky130_fd_sc_hd__dfxtp_1 _876_ (.CLK(clknet_3_6__leaf_clk),
    .D(_020_),
    .Q(\debounce1_a.button_hist[0] ));
 sky130_fd_sc_hd__dfxtp_1 _877_ (.CLK(clknet_3_6__leaf_clk),
    .D(_021_),
    .Q(\debounce1_a.button_hist[1] ));
 sky130_fd_sc_hd__dfxtp_1 _878_ (.CLK(clknet_3_6__leaf_clk),
    .D(_022_),
    .Q(\debounce1_a.button_hist[2] ));
 sky130_fd_sc_hd__dfxtp_1 _879_ (.CLK(clknet_3_6__leaf_clk),
    .D(_023_),
    .Q(\debounce1_a.button_hist[3] ));
 sky130_fd_sc_hd__dfxtp_1 _880_ (.CLK(clknet_3_6__leaf_clk),
    .D(_024_),
    .Q(\debounce1_a.button_hist[4] ));
 sky130_fd_sc_hd__dfxtp_1 _881_ (.CLK(clknet_3_6__leaf_clk),
    .D(_025_),
    .Q(\debounce1_a.button_hist[5] ));
 sky130_fd_sc_hd__dfxtp_1 _882_ (.CLK(clknet_3_6__leaf_clk),
    .D(_026_),
    .Q(\debounce1_a.button_hist[6] ));
 sky130_fd_sc_hd__dfxtp_1 _883_ (.CLK(clknet_3_6__leaf_clk),
    .D(_027_),
    .Q(\debounce1_a.button_hist[7] ));
 sky130_fd_sc_hd__dfxtp_1 _884_ (.CLK(clknet_3_5__leaf_clk),
    .D(net39),
    .Q(\debounce1_b.debounced ));
 sky130_fd_sc_hd__dfxtp_1 _885_ (.CLK(clknet_3_5__leaf_clk),
    .D(_029_),
    .Q(\debounce1_b.button_hist[0] ));
 sky130_fd_sc_hd__dfxtp_1 _886_ (.CLK(clknet_3_5__leaf_clk),
    .D(_030_),
    .Q(\debounce1_b.button_hist[1] ));
 sky130_fd_sc_hd__dfxtp_1 _887_ (.CLK(clknet_3_5__leaf_clk),
    .D(_031_),
    .Q(\debounce1_b.button_hist[2] ));
 sky130_fd_sc_hd__dfxtp_1 _888_ (.CLK(clknet_3_5__leaf_clk),
    .D(_032_),
    .Q(\debounce1_b.button_hist[3] ));
 sky130_fd_sc_hd__dfxtp_1 _889_ (.CLK(clknet_3_5__leaf_clk),
    .D(_033_),
    .Q(\debounce1_b.button_hist[4] ));
 sky130_fd_sc_hd__dfxtp_1 _890_ (.CLK(clknet_3_5__leaf_clk),
    .D(_034_),
    .Q(\debounce1_b.button_hist[5] ));
 sky130_fd_sc_hd__dfxtp_1 _891_ (.CLK(clknet_3_5__leaf_clk),
    .D(_035_),
    .Q(\debounce1_b.button_hist[6] ));
 sky130_fd_sc_hd__dfxtp_1 _892_ (.CLK(clknet_3_5__leaf_clk),
    .D(_036_),
    .Q(\debounce1_b.button_hist[7] ));
 sky130_fd_sc_hd__dfxtp_1 _893_ (.CLK(clknet_3_4__leaf_clk),
    .D(net43),
    .Q(\debounce2_a.debounced ));
 sky130_fd_sc_hd__dfxtp_1 _894_ (.CLK(clknet_3_4__leaf_clk),
    .D(_038_),
    .Q(\debounce2_a.button_hist[0] ));
 sky130_fd_sc_hd__dfxtp_1 _895_ (.CLK(clknet_3_4__leaf_clk),
    .D(_039_),
    .Q(\debounce2_a.button_hist[1] ));
 sky130_fd_sc_hd__dfxtp_1 _896_ (.CLK(clknet_3_4__leaf_clk),
    .D(_040_),
    .Q(\debounce2_a.button_hist[2] ));
 sky130_fd_sc_hd__dfxtp_1 _897_ (.CLK(clknet_3_4__leaf_clk),
    .D(_041_),
    .Q(\debounce2_a.button_hist[3] ));
 sky130_fd_sc_hd__dfxtp_1 _898_ (.CLK(clknet_3_4__leaf_clk),
    .D(_042_),
    .Q(\debounce2_a.button_hist[4] ));
 sky130_fd_sc_hd__dfxtp_1 _899_ (.CLK(clknet_3_4__leaf_clk),
    .D(_043_),
    .Q(\debounce2_a.button_hist[5] ));
 sky130_fd_sc_hd__dfxtp_1 _900_ (.CLK(clknet_3_5__leaf_clk),
    .D(_044_),
    .Q(\debounce2_a.button_hist[6] ));
 sky130_fd_sc_hd__dfxtp_1 _901_ (.CLK(clknet_3_4__leaf_clk),
    .D(_045_),
    .Q(\debounce2_a.button_hist[7] ));
 sky130_fd_sc_hd__dfxtp_1 _902_ (.CLK(clknet_3_1__leaf_clk),
    .D(net35),
    .Q(\debounce2_b.debounced ));
 sky130_fd_sc_hd__dfxtp_1 _903_ (.CLK(clknet_3_2__leaf_clk),
    .D(net29),
    .Q(\pwm2.count[0] ));
 sky130_fd_sc_hd__dfxtp_1 _904_ (.CLK(clknet_3_2__leaf_clk),
    .D(net174),
    .Q(\pwm2.count[1] ));
 sky130_fd_sc_hd__dfxtp_1 _905_ (.CLK(clknet_3_0__leaf_clk),
    .D(net65),
    .Q(\pwm2.count[2] ));
 sky130_fd_sc_hd__dfxtp_1 _906_ (.CLK(clknet_3_0__leaf_clk),
    .D(_050_),
    .Q(\pwm2.count[3] ));
 sky130_fd_sc_hd__dfxtp_1 _907_ (.CLK(clknet_3_0__leaf_clk),
    .D(net51),
    .Q(\pwm2.count[4] ));
 sky130_fd_sc_hd__dfxtp_1 _908_ (.CLK(clknet_3_0__leaf_clk),
    .D(net72),
    .Q(\pwm2.count[5] ));
 sky130_fd_sc_hd__dfxtp_1 _909_ (.CLK(clknet_3_0__leaf_clk),
    .D(net53),
    .Q(\pwm2.count[6] ));
 sky130_fd_sc_hd__dfxtp_1 _910_ (.CLK(clknet_3_0__leaf_clk),
    .D(net76),
    .Q(\pwm2.count[7] ));
 sky130_fd_sc_hd__dfxtp_1 _911_ (.CLK(clknet_3_5__leaf_clk),
    .D(_055_),
    .Q(\encoder0.old_a ));
 sky130_fd_sc_hd__dfxtp_1 _912_ (.CLK(clknet_3_1__leaf_clk),
    .D(_056_),
    .Q(\debounce2_b.button_hist[0] ));
 sky130_fd_sc_hd__dfxtp_1 _913_ (.CLK(clknet_3_1__leaf_clk),
    .D(_057_),
    .Q(\debounce2_b.button_hist[1] ));
 sky130_fd_sc_hd__dfxtp_1 _914_ (.CLK(clknet_3_1__leaf_clk),
    .D(_058_),
    .Q(\debounce2_b.button_hist[2] ));
 sky130_fd_sc_hd__dfxtp_1 _915_ (.CLK(clknet_3_1__leaf_clk),
    .D(_059_),
    .Q(\debounce2_b.button_hist[3] ));
 sky130_fd_sc_hd__dfxtp_1 _916_ (.CLK(clknet_3_1__leaf_clk),
    .D(_060_),
    .Q(\debounce2_b.button_hist[4] ));
 sky130_fd_sc_hd__dfxtp_1 _917_ (.CLK(clknet_3_4__leaf_clk),
    .D(_061_),
    .Q(\debounce2_b.button_hist[5] ));
 sky130_fd_sc_hd__dfxtp_1 _918_ (.CLK(clknet_3_4__leaf_clk),
    .D(_062_),
    .Q(\debounce2_b.button_hist[6] ));
 sky130_fd_sc_hd__dfxtp_1 _919_ (.CLK(clknet_3_1__leaf_clk),
    .D(_063_),
    .Q(\debounce2_b.button_hist[7] ));
 sky130_fd_sc_hd__dfxtp_1 _920_ (.CLK(clknet_3_4__leaf_clk),
    .D(net130),
    .Q(\encoder0.value[0] ));
 sky130_fd_sc_hd__dfxtp_1 _921_ (.CLK(clknet_3_4__leaf_clk),
    .D(net102),
    .Q(\encoder0.value[1] ));
 sky130_fd_sc_hd__dfxtp_1 _922_ (.CLK(clknet_3_5__leaf_clk),
    .D(net142),
    .Q(\encoder0.value[2] ));
 sky130_fd_sc_hd__dfxtp_1 _923_ (.CLK(clknet_3_4__leaf_clk),
    .D(net144),
    .Q(\encoder0.value[3] ));
 sky130_fd_sc_hd__dfxtp_1 _924_ (.CLK(clknet_3_7__leaf_clk),
    .D(net166),
    .Q(\encoder0.value[4] ));
 sky130_fd_sc_hd__dfxtp_1 _925_ (.CLK(clknet_3_6__leaf_clk),
    .D(net162),
    .Q(\encoder0.value[5] ));
 sky130_fd_sc_hd__dfxtp_1 _926_ (.CLK(clknet_3_7__leaf_clk),
    .D(_070_),
    .Q(\encoder0.value[6] ));
 sky130_fd_sc_hd__dfxtp_1 _927_ (.CLK(clknet_3_6__leaf_clk),
    .D(net125),
    .Q(\encoder0.value[7] ));
 sky130_fd_sc_hd__dfxtp_1 _928_ (.CLK(clknet_3_6__leaf_clk),
    .D(_072_),
    .Q(\encoder1.old_a ));
 sky130_fd_sc_hd__dfxtp_1 _929_ (.CLK(clknet_3_5__leaf_clk),
    .D(_073_),
    .Q(\encoder0.old_b ));
 sky130_fd_sc_hd__dfxtp_1 _930_ (.CLK(clknet_3_3__leaf_clk),
    .D(net152),
    .Q(\encoder1.value[0] ));
 sky130_fd_sc_hd__dfxtp_1 _931_ (.CLK(clknet_3_3__leaf_clk),
    .D(net108),
    .Q(\encoder1.value[1] ));
 sky130_fd_sc_hd__dfxtp_1 _932_ (.CLK(clknet_3_3__leaf_clk),
    .D(net132),
    .Q(\encoder1.value[2] ));
 sky130_fd_sc_hd__dfxtp_1 _933_ (.CLK(clknet_3_3__leaf_clk),
    .D(net146),
    .Q(\encoder1.value[3] ));
 sky130_fd_sc_hd__dfxtp_1 _934_ (.CLK(clknet_3_2__leaf_clk),
    .D(net134),
    .Q(\encoder1.value[4] ));
 sky130_fd_sc_hd__dfxtp_1 _935_ (.CLK(clknet_3_2__leaf_clk),
    .D(net150),
    .Q(\encoder1.value[5] ));
 sky130_fd_sc_hd__dfxtp_1 _936_ (.CLK(clknet_3_2__leaf_clk),
    .D(_080_),
    .Q(\encoder1.value[6] ));
 sky130_fd_sc_hd__dfxtp_1 _937_ (.CLK(clknet_3_2__leaf_clk),
    .D(net120),
    .Q(\encoder1.value[7] ));
 sky130_fd_sc_hd__dfxtp_1 _938_ (.CLK(clknet_3_4__leaf_clk),
    .D(_082_),
    .Q(\encoder2.old_a ));
 sky130_fd_sc_hd__dfxtp_1 _939_ (.CLK(clknet_3_3__leaf_clk),
    .D(_083_),
    .Q(\encoder1.old_b ));
 sky130_fd_sc_hd__dfxtp_1 _940_ (.CLK(clknet_3_0__leaf_clk),
    .D(net148),
    .Q(\encoder2.value[0] ));
 sky130_fd_sc_hd__dfxtp_1 _941_ (.CLK(clknet_3_2__leaf_clk),
    .D(net105),
    .Q(\encoder2.value[1] ));
 sky130_fd_sc_hd__dfxtp_1 _942_ (.CLK(clknet_3_3__leaf_clk),
    .D(net136),
    .Q(\encoder2.value[2] ));
 sky130_fd_sc_hd__dfxtp_1 _943_ (.CLK(clknet_3_0__leaf_clk),
    .D(net128),
    .Q(\encoder2.value[3] ));
 sky130_fd_sc_hd__dfxtp_1 _944_ (.CLK(clknet_3_1__leaf_clk),
    .D(net140),
    .Q(\encoder2.value[4] ));
 sky130_fd_sc_hd__dfxtp_1 _945_ (.CLK(clknet_3_1__leaf_clk),
    .D(net158),
    .Q(\encoder2.value[5] ));
 sky130_fd_sc_hd__dfxtp_1 _946_ (.CLK(clknet_3_0__leaf_clk),
    .D(_090_),
    .Q(\encoder2.value[6] ));
 sky130_fd_sc_hd__dfxtp_1 _947_ (.CLK(clknet_3_0__leaf_clk),
    .D(net115),
    .Q(\encoder2.value[7] ));
 sky130_fd_sc_hd__dfxtp_1 _948_ (.CLK(clknet_3_1__leaf_clk),
    .D(_092_),
    .Q(\encoder2.old_b ));
 sky130_fd_sc_hd__dfxtp_1 _949_ (.CLK(clknet_3_1__leaf_clk),
    .D(net27),
    .Q(\pwm0.count[0] ));
 sky130_fd_sc_hd__dfxtp_1 _950_ (.CLK(clknet_3_4__leaf_clk),
    .D(net55),
    .Q(\pwm0.count[1] ));
 sky130_fd_sc_hd__dfxtp_1 _951_ (.CLK(clknet_3_3__leaf_clk),
    .D(net59),
    .Q(\pwm0.count[2] ));
 sky130_fd_sc_hd__dfxtp_1 _952_ (.CLK(clknet_3_3__leaf_clk),
    .D(_096_),
    .Q(\pwm0.count[3] ));
 sky130_fd_sc_hd__dfxtp_1 _953_ (.CLK(clknet_3_3__leaf_clk),
    .D(net47),
    .Q(\pwm0.count[4] ));
 sky130_fd_sc_hd__dfxtp_1 _954_ (.CLK(clknet_3_3__leaf_clk),
    .D(net70),
    .Q(\pwm0.count[5] ));
 sky130_fd_sc_hd__dfxtp_1 _955_ (.CLK(clknet_3_3__leaf_clk),
    .D(net45),
    .Q(\pwm0.count[6] ));
 sky130_fd_sc_hd__dfxtp_1 _956_ (.CLK(clknet_3_3__leaf_clk),
    .D(net57),
    .Q(\pwm0.count[7] ));
 sky130_fd_sc_hd__dfxtp_1 _957_ (.CLK(clknet_3_3__leaf_clk),
    .D(net41),
    .Q(\pwm1.count[0] ));
 sky130_fd_sc_hd__dfxtp_1 _958_ (.CLK(clknet_3_3__leaf_clk),
    .D(net176),
    .Q(\pwm1.count[1] ));
 sky130_fd_sc_hd__dfxtp_1 _959_ (.CLK(clknet_3_3__leaf_clk),
    .D(net67),
    .Q(\pwm1.count[2] ));
 sky130_fd_sc_hd__dfxtp_1 _960_ (.CLK(clknet_3_2__leaf_clk),
    .D(_104_),
    .Q(\pwm1.count[3] ));
 sky130_fd_sc_hd__dfxtp_1 _961_ (.CLK(clknet_3_2__leaf_clk),
    .D(net62),
    .Q(\pwm1.count[4] ));
 sky130_fd_sc_hd__dfxtp_1 _962_ (.CLK(clknet_3_2__leaf_clk),
    .D(net74),
    .Q(\pwm1.count[5] ));
 sky130_fd_sc_hd__dfxtp_1 _963_ (.CLK(clknet_3_2__leaf_clk),
    .D(net49),
    .Q(\pwm1.count[6] ));
 sky130_fd_sc_hd__dfxtp_1 _964_ (.CLK(clknet_3_2__leaf_clk),
    .D(_108_),
    .Q(\pwm1.count[7] ));
 sky130_fd_sc_hd__buf_2 _976_ (.A(net7),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(net171),
    .X(net23));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(\debounce0_b.button_hist[5] ),
    .X(net32));
 sky130_fd_sc_hd__dlygate4sd3_1 hold100 (.A(\debounce2_a.button_hist[4] ),
    .X(net122));
 sky130_fd_sc_hd__dlygate4sd3_1 hold101 (.A(\debounce1_b.button_hist[6] ),
    .X(net123));
 sky130_fd_sc_hd__dlygate4sd3_1 hold102 (.A(\encoder0.value[7] ),
    .X(net124));
 sky130_fd_sc_hd__dlygate4sd3_1 hold103 (.A(_071_),
    .X(net125));
 sky130_fd_sc_hd__dlygate4sd3_1 hold104 (.A(\debounce1_a.button_hist[6] ),
    .X(net126));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold105 (.A(\encoder2.value[3] ),
    .X(net127));
 sky130_fd_sc_hd__dlygate4sd3_1 hold106 (.A(_087_),
    .X(net128));
 sky130_fd_sc_hd__buf_1 hold107 (.A(\encoder0.value[0] ),
    .X(net129));
 sky130_fd_sc_hd__dlygate4sd3_1 hold108 (.A(_064_),
    .X(net130));
 sky130_fd_sc_hd__buf_1 hold109 (.A(\encoder1.value[2] ),
    .X(net131));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(_010_),
    .X(net33));
 sky130_fd_sc_hd__dlygate4sd3_1 hold110 (.A(_076_),
    .X(net132));
 sky130_fd_sc_hd__buf_1 hold111 (.A(\encoder1.value[4] ),
    .X(net133));
 sky130_fd_sc_hd__dlygate4sd3_1 hold112 (.A(_078_),
    .X(net134));
 sky130_fd_sc_hd__buf_1 hold113 (.A(\encoder2.value[2] ),
    .X(net135));
 sky130_fd_sc_hd__dlygate4sd3_1 hold114 (.A(_086_),
    .X(net136));
 sky130_fd_sc_hd__dlygate4sd3_1 hold115 (.A(\debounce0_a.button_hist[6] ),
    .X(net137));
 sky130_fd_sc_hd__dlygate4sd3_1 hold116 (.A(\pwm1.count[7] ),
    .X(net138));
 sky130_fd_sc_hd__buf_1 hold117 (.A(\encoder2.value[4] ),
    .X(net139));
 sky130_fd_sc_hd__dlygate4sd3_1 hold118 (.A(_088_),
    .X(net140));
 sky130_fd_sc_hd__buf_1 hold119 (.A(\encoder0.value[2] ),
    .X(net141));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(\debounce2_b.button_hist[5] ),
    .X(net34));
 sky130_fd_sc_hd__dlygate4sd3_1 hold120 (.A(_066_),
    .X(net142));
 sky130_fd_sc_hd__buf_1 hold121 (.A(\encoder0.value[3] ),
    .X(net143));
 sky130_fd_sc_hd__dlygate4sd3_1 hold122 (.A(_067_),
    .X(net144));
 sky130_fd_sc_hd__buf_1 hold123 (.A(\encoder1.value[3] ),
    .X(net145));
 sky130_fd_sc_hd__dlygate4sd3_1 hold124 (.A(_077_),
    .X(net146));
 sky130_fd_sc_hd__dlygate4sd3_1 hold125 (.A(\encoder2.value[0] ),
    .X(net147));
 sky130_fd_sc_hd__dlygate4sd3_1 hold126 (.A(_084_),
    .X(net148));
 sky130_fd_sc_hd__buf_1 hold127 (.A(\encoder1.value[5] ),
    .X(net149));
 sky130_fd_sc_hd__dlygate4sd3_1 hold128 (.A(_079_),
    .X(net150));
 sky130_fd_sc_hd__dlygate4sd3_1 hold129 (.A(\encoder1.value[0] ),
    .X(net151));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(_046_),
    .X(net35));
 sky130_fd_sc_hd__dlygate4sd3_1 hold130 (.A(_074_),
    .X(net152));
 sky130_fd_sc_hd__buf_1 hold131 (.A(\encoder1.value[6] ),
    .X(net153));
 sky130_fd_sc_hd__dlygate4sd3_1 hold132 (.A(_349_),
    .X(net154));
 sky130_fd_sc_hd__dlygate4sd3_1 hold133 (.A(\debounce0_a.debounced ),
    .X(net155));
 sky130_fd_sc_hd__dlygate4sd3_1 hold134 (.A(\debounce2_b.debounced ),
    .X(net156));
 sky130_fd_sc_hd__buf_1 hold135 (.A(\encoder2.value[5] ),
    .X(net157));
 sky130_fd_sc_hd__dlygate4sd3_1 hold136 (.A(_089_),
    .X(net158));
 sky130_fd_sc_hd__buf_1 hold137 (.A(\encoder2.value[6] ),
    .X(net159));
 sky130_fd_sc_hd__dlygate4sd3_1 hold138 (.A(_397_),
    .X(net160));
 sky130_fd_sc_hd__buf_1 hold139 (.A(\encoder0.value[5] ),
    .X(net161));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(\debounce0_a.button_hist[5] ),
    .X(net36));
 sky130_fd_sc_hd__dlygate4sd3_1 hold140 (.A(_069_),
    .X(net162));
 sky130_fd_sc_hd__dlygate4sd3_1 hold141 (.A(\debounce0_b.debounced ),
    .X(net163));
 sky130_fd_sc_hd__dlygate4sd3_1 hold142 (.A(\debounce1_a.debounced ),
    .X(net164));
 sky130_fd_sc_hd__buf_1 hold143 (.A(\encoder0.value[4] ),
    .X(net165));
 sky130_fd_sc_hd__dlygate4sd3_1 hold144 (.A(_068_),
    .X(net166));
 sky130_fd_sc_hd__dlygate4sd3_1 hold145 (.A(\debounce2_a.debounced ),
    .X(net167));
 sky130_fd_sc_hd__dlygate4sd3_1 hold146 (.A(\debounce1_b.debounced ),
    .X(net168));
 sky130_fd_sc_hd__dlygate4sd3_1 hold147 (.A(\encoder0.value[6] ),
    .X(net169));
 sky130_fd_sc_hd__dlygate4sd3_1 hold148 (.A(_300_),
    .X(net170));
 sky130_fd_sc_hd__dlygate4sd3_1 hold149 (.A(reset),
    .X(net171));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(_001_),
    .X(net37));
 sky130_fd_sc_hd__dlygate4sd3_1 hold150 (.A(net23),
    .X(net172));
 sky130_fd_sc_hd__dlygate4sd3_1 hold151 (.A(\pwm2.count[1] ),
    .X(net173));
 sky130_fd_sc_hd__dlygate4sd3_1 hold152 (.A(_048_),
    .X(net174));
 sky130_fd_sc_hd__dlygate4sd3_1 hold153 (.A(\pwm1.count[1] ),
    .X(net175));
 sky130_fd_sc_hd__dlygate4sd3_1 hold154 (.A(_102_),
    .X(net176));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(\debounce1_b.button_hist[5] ),
    .X(net38));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(_028_),
    .X(net39));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold18 (.A(\pwm1.count[0] ),
    .X(net40));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(_101_),
    .X(net41));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(net7),
    .X(net24));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(\debounce2_a.button_hist[5] ),
    .X(net42));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(_037_),
    .X(net43));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(\pwm0.count[6] ),
    .X(net44));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(_099_),
    .X(net45));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(\pwm0.count[4] ),
    .X(net46));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(_097_),
    .X(net47));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(\pwm1.count[6] ),
    .X(net48));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(_107_),
    .X(net49));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(\pwm2.count[4] ),
    .X(net50));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(_051_),
    .X(net51));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(_000_),
    .X(net25));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(\pwm2.count[6] ),
    .X(net52));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(_053_),
    .X(net53));
 sky130_fd_sc_hd__buf_1 hold32 (.A(\pwm0.count[1] ),
    .X(net54));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(_094_),
    .X(net55));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(\pwm0.count[7] ),
    .X(net56));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(_100_),
    .X(net57));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(\pwm0.count[2] ),
    .X(net58));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(_095_),
    .X(net59));
 sky130_fd_sc_hd__buf_1 hold38 (.A(net173),
    .X(net60));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(\pwm1.count[4] ),
    .X(net61));
 sky130_fd_sc_hd__buf_1 hold4 (.A(\pwm0.count[0] ),
    .X(net26));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(_105_),
    .X(net62));
 sky130_fd_sc_hd__buf_1 hold41 (.A(net175),
    .X(net63));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(\pwm2.count[2] ),
    .X(net64));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(_049_),
    .X(net65));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(\pwm1.count[2] ),
    .X(net66));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(_103_),
    .X(net67));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(\debounce0_a.reset ),
    .X(net68));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(\pwm0.count[5] ),
    .X(net69));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(_098_),
    .X(net70));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(\pwm2.count[5] ),
    .X(net71));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(_093_),
    .X(net27));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(_052_),
    .X(net72));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(\pwm1.count[5] ),
    .X(net73));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(_106_),
    .X(net74));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(\pwm2.count[7] ),
    .X(net75));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(_054_),
    .X(net76));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(\debounce0_a.button_hist[2] ),
    .X(net77));
 sky130_fd_sc_hd__dlygate4sd3_1 hold56 (.A(\debounce2_b.button_hist[4] ),
    .X(net78));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(\debounce2_b.button_hist[3] ),
    .X(net79));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(\debounce2_b.button_hist[2] ),
    .X(net80));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(\pwm1.count[3] ),
    .X(net81));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold6 (.A(\pwm2.count[0] ),
    .X(net28));
 sky130_fd_sc_hd__dlygate4sd3_1 hold60 (.A(\debounce0_b.button_hist[3] ),
    .X(net82));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(\debounce2_a.button_hist[6] ),
    .X(net83));
 sky130_fd_sc_hd__dlygate4sd3_1 hold62 (.A(\debounce2_b.button_hist[0] ),
    .X(net84));
 sky130_fd_sc_hd__dlygate4sd3_1 hold63 (.A(\pwm2.count[3] ),
    .X(net85));
 sky130_fd_sc_hd__dlygate4sd3_1 hold64 (.A(\debounce1_b.button_hist[1] ),
    .X(net86));
 sky130_fd_sc_hd__dlygate4sd3_1 hold65 (.A(\debounce2_b.button_hist[1] ),
    .X(net87));
 sky130_fd_sc_hd__dlygate4sd3_1 hold66 (.A(\debounce2_a.button_hist[3] ),
    .X(net88));
 sky130_fd_sc_hd__dlygate4sd3_1 hold67 (.A(\debounce0_a.button_hist[3] ),
    .X(net89));
 sky130_fd_sc_hd__dlygate4sd3_1 hold68 (.A(\debounce0_b.button_hist[1] ),
    .X(net90));
 sky130_fd_sc_hd__dlygate4sd3_1 hold69 (.A(\debounce1_a.button_hist[1] ),
    .X(net91));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(_047_),
    .X(net29));
 sky130_fd_sc_hd__dlygate4sd3_1 hold70 (.A(\debounce1_a.button_hist[3] ),
    .X(net92));
 sky130_fd_sc_hd__dlygate4sd3_1 hold71 (.A(\debounce2_a.button_hist[2] ),
    .X(net93));
 sky130_fd_sc_hd__dlygate4sd3_1 hold72 (.A(\debounce1_a.button_hist[0] ),
    .X(net94));
 sky130_fd_sc_hd__dlygate4sd3_1 hold73 (.A(\debounce1_a.button_hist[2] ),
    .X(net95));
 sky130_fd_sc_hd__dlygate4sd3_1 hold74 (.A(\debounce1_b.button_hist[3] ),
    .X(net96));
 sky130_fd_sc_hd__dlygate4sd3_1 hold75 (.A(\debounce0_b.button_hist[2] ),
    .X(net97));
 sky130_fd_sc_hd__dlygate4sd3_1 hold76 (.A(\debounce1_b.button_hist[2] ),
    .X(net98));
 sky130_fd_sc_hd__dlygate4sd3_1 hold77 (.A(\pwm0.count[3] ),
    .X(net99));
 sky130_fd_sc_hd__dlygate4sd3_1 hold78 (.A(\debounce0_a.button_hist[1] ),
    .X(net100));
 sky130_fd_sc_hd__dlygate4sd3_1 hold79 (.A(\encoder0.value[1] ),
    .X(net101));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(\debounce1_a.button_hist[5] ),
    .X(net30));
 sky130_fd_sc_hd__dlygate4sd3_1 hold80 (.A(_065_),
    .X(net102));
 sky130_fd_sc_hd__dlygate4sd3_1 hold81 (.A(\debounce2_a.button_hist[1] ),
    .X(net103));
 sky130_fd_sc_hd__dlygate4sd3_1 hold82 (.A(\encoder2.value[1] ),
    .X(net104));
 sky130_fd_sc_hd__dlygate4sd3_1 hold83 (.A(_085_),
    .X(net105));
 sky130_fd_sc_hd__dlygate4sd3_1 hold84 (.A(\debounce2_a.button_hist[0] ),
    .X(net106));
 sky130_fd_sc_hd__dlygate4sd3_1 hold85 (.A(\encoder1.value[1] ),
    .X(net107));
 sky130_fd_sc_hd__dlygate4sd3_1 hold86 (.A(_075_),
    .X(net108));
 sky130_fd_sc_hd__dlygate4sd3_1 hold87 (.A(\debounce0_b.button_hist[6] ),
    .X(net109));
 sky130_fd_sc_hd__dlygate4sd3_1 hold88 (.A(\debounce0_a.button_hist[0] ),
    .X(net110));
 sky130_fd_sc_hd__dlygate4sd3_1 hold89 (.A(\debounce1_b.button_hist[0] ),
    .X(net111));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(_019_),
    .X(net31));
 sky130_fd_sc_hd__dlygate4sd3_1 hold90 (.A(\debounce2_b.button_hist[6] ),
    .X(net112));
 sky130_fd_sc_hd__dlygate4sd3_1 hold91 (.A(\debounce1_b.button_hist[4] ),
    .X(net113));
 sky130_fd_sc_hd__dlygate4sd3_1 hold92 (.A(\encoder2.value[7] ),
    .X(net114));
 sky130_fd_sc_hd__dlygate4sd3_1 hold93 (.A(_091_),
    .X(net115));
 sky130_fd_sc_hd__dlygate4sd3_1 hold94 (.A(\debounce1_a.button_hist[4] ),
    .X(net116));
 sky130_fd_sc_hd__dlygate4sd3_1 hold95 (.A(\debounce0_a.button_hist[4] ),
    .X(net117));
 sky130_fd_sc_hd__dlygate4sd3_1 hold96 (.A(\debounce0_b.button_hist[0] ),
    .X(net118));
 sky130_fd_sc_hd__dlygate4sd3_1 hold97 (.A(\encoder1.value[7] ),
    .X(net119));
 sky130_fd_sc_hd__dlygate4sd3_1 hold98 (.A(_081_),
    .X(net120));
 sky130_fd_sc_hd__dlygate4sd3_1 hold99 (.A(\debounce0_b.button_hist[4] ),
    .X(net121));
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(enc0_a),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(enc0_b),
    .X(net2));
 sky130_fd_sc_hd__buf_1 input3 (.A(enc1_a),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(enc1_b),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(enc2_a),
    .X(net5));
 sky130_fd_sc_hd__buf_1 input6 (.A(enc2_b),
    .X(net6));
 sky130_fd_sc_hd__buf_1 input7 (.A(net172),
    .X(net7));
 sky130_fd_sc_hd__buf_12 output10 (.A(net10),
    .X(pwm2_out));
 sky130_fd_sc_hd__buf_12 output11 (.A(net11),
    .X(sync));
 sky130_fd_sc_hd__buf_12 output8 (.A(net8),
    .X(pwm0_out));
 sky130_fd_sc_hd__buf_12 output9 (.A(net9),
    .X(pwm1_out));
 sky130_fd_sc_hd__conb_1 rgb_mixer_13 (.LO(net13));
 sky130_fd_sc_hd__conb_1 rgb_mixer_14 (.LO(net14));
 sky130_fd_sc_hd__conb_1 rgb_mixer_15 (.LO(net15));
 sky130_fd_sc_hd__conb_1 rgb_mixer_16 (.LO(net16));
 sky130_fd_sc_hd__conb_1 rgb_mixer_17 (.HI(net17));
 sky130_fd_sc_hd__conb_1 rgb_mixer_18 (.HI(net18));
 sky130_fd_sc_hd__conb_1 rgb_mixer_19 (.HI(net19));
 sky130_fd_sc_hd__conb_1 rgb_mixer_20 (.HI(net20));
 sky130_fd_sc_hd__conb_1 rgb_mixer_21 (.HI(net21));
 sky130_fd_sc_hd__conb_1 rgb_mixer_22 (.HI(net22));
 assign io_oeb_high[0] = net17;
 assign io_oeb_high[1] = net18;
 assign io_oeb_high[2] = net19;
 assign io_oeb_high[3] = net20;
 assign io_oeb_high[4] = net21;
 assign io_oeb_high[5] = net22;
 assign io_oeb_low[0] = net13;
 assign io_oeb_low[1] = net14;
 assign io_oeb_low[2] = net15;
 assign io_oeb_low[3] = net16;
endmodule

