magic
tech sky130A
magscale 1 2
timestamp 1696494444
<< viali >>
rect 17785 39593 17819 39627
rect 14657 39457 14691 39491
rect 16405 39457 16439 39491
rect 17877 39457 17911 39491
rect 22477 39457 22511 39491
rect 34529 39457 34563 39491
rect 1409 39389 1443 39423
rect 1777 39389 1811 39423
rect 2421 39389 2455 39423
rect 2513 39389 2547 39423
rect 3065 39389 3099 39423
rect 8677 39389 8711 39423
rect 14473 39389 14507 39423
rect 15117 39389 15151 39423
rect 15485 39389 15519 39423
rect 15669 39389 15703 39423
rect 15761 39389 15795 39423
rect 16865 39389 16899 39423
rect 17509 39389 17543 39423
rect 17601 39389 17635 39423
rect 18061 39389 18095 39423
rect 18245 39389 18279 39423
rect 20729 39389 20763 39423
rect 21281 39389 21315 39423
rect 22201 39389 22235 39423
rect 17785 39321 17819 39355
rect 1593 39253 1627 39287
rect 8493 39253 8527 39287
rect 14289 39253 14323 39287
rect 14933 39253 14967 39287
rect 15301 39253 15335 39287
rect 17049 39253 17083 39287
rect 17325 39253 17359 39287
rect 20545 39253 20579 39287
rect 21465 39253 21499 39287
rect 2053 39049 2087 39083
rect 14013 39049 14047 39083
rect 15485 39049 15519 39083
rect 21557 39049 21591 39083
rect 14372 38981 14406 39015
rect 17386 38981 17420 39015
rect 20444 38981 20478 39015
rect 22946 38981 22980 39015
rect 1409 38913 1443 38947
rect 13829 38913 13863 38947
rect 15577 38913 15611 38947
rect 16681 38913 16715 38947
rect 16865 38913 16899 38947
rect 23305 38913 23339 38947
rect 14105 38845 14139 38879
rect 15945 38845 15979 38879
rect 16497 38845 16531 38879
rect 17049 38845 17083 38879
rect 17141 38845 17175 38879
rect 20177 38845 20211 38879
rect 23213 38845 23247 38879
rect 15761 38709 15795 38743
rect 18521 38709 18555 38743
rect 21833 38709 21867 38743
rect 23949 38709 23983 38743
rect 18153 38505 18187 38539
rect 22753 38505 22787 38539
rect 23213 38505 23247 38539
rect 21005 38437 21039 38471
rect 15853 38369 15887 38403
rect 18981 38369 19015 38403
rect 21281 38369 21315 38403
rect 21925 38369 21959 38403
rect 23121 38369 23155 38403
rect 23581 38369 23615 38403
rect 4905 38301 4939 38335
rect 8401 38301 8435 38335
rect 8493 38301 8527 38335
rect 13737 38301 13771 38335
rect 14197 38301 14231 38335
rect 17601 38301 17635 38335
rect 19625 38301 19659 38335
rect 22017 38301 22051 38335
rect 22937 38301 22971 38335
rect 23397 38301 23431 38335
rect 14442 38233 14476 38267
rect 16098 38233 16132 38267
rect 19892 38233 19926 38267
rect 5457 38165 5491 38199
rect 8677 38165 8711 38199
rect 13921 38165 13955 38199
rect 15577 38165 15611 38199
rect 17233 38165 17267 38199
rect 18429 38165 18463 38199
rect 22661 38165 22695 38199
rect 14657 37961 14691 37995
rect 17693 37961 17727 37995
rect 17969 37961 18003 37995
rect 20729 37961 20763 37995
rect 22109 37961 22143 37995
rect 14994 37893 15028 37927
rect 17785 37893 17819 37927
rect 21833 37893 21867 37927
rect 22017 37893 22051 37927
rect 8861 37825 8895 37859
rect 10333 37825 10367 37859
rect 10425 37825 10459 37859
rect 10609 37825 10643 37859
rect 10701 37825 10735 37859
rect 10885 37825 10919 37859
rect 11161 37825 11195 37859
rect 11713 37825 11747 37859
rect 13093 37825 13127 37859
rect 14473 37825 14507 37859
rect 17509 37825 17543 37859
rect 19082 37825 19116 37859
rect 19625 37825 19659 37859
rect 19717 37825 19751 37859
rect 20453 37825 20487 37859
rect 20637 37825 20671 37859
rect 20913 37825 20947 37859
rect 21373 37825 21407 37859
rect 21465 37825 21499 37859
rect 21649 37825 21683 37859
rect 22201 37825 22235 37859
rect 11069 37757 11103 37791
rect 11897 37757 11931 37791
rect 14749 37757 14783 37791
rect 17417 37757 17451 37791
rect 17877 37757 17911 37791
rect 19349 37757 19383 37791
rect 20269 37757 20303 37791
rect 22569 37757 22603 37791
rect 23213 37757 23247 37791
rect 11345 37689 11379 37723
rect 16129 37689 16163 37723
rect 7389 37621 7423 37655
rect 9045 37621 9079 37655
rect 10149 37621 10183 37655
rect 10885 37621 10919 37655
rect 11529 37621 11563 37655
rect 12449 37621 12483 37655
rect 12909 37621 12943 37655
rect 17233 37621 17267 37655
rect 19441 37621 19475 37655
rect 21189 37621 21223 37655
rect 21649 37621 21683 37655
rect 22385 37621 22419 37655
rect 10977 37417 11011 37451
rect 14105 37417 14139 37451
rect 15025 37417 15059 37451
rect 17325 37417 17359 37451
rect 17509 37417 17543 37451
rect 18337 37417 18371 37451
rect 19073 37417 19107 37451
rect 17785 37349 17819 37383
rect 7297 37281 7331 37315
rect 16129 37281 16163 37315
rect 17417 37281 17451 37315
rect 22385 37281 22419 37315
rect 6929 37213 6963 37247
rect 9597 37213 9631 37247
rect 11069 37213 11103 37247
rect 12541 37213 12575 37247
rect 14289 37213 14323 37247
rect 14381 37213 14415 37247
rect 15209 37213 15243 37247
rect 15393 37213 15427 37247
rect 15485 37213 15519 37247
rect 16865 37213 16899 37247
rect 17233 37213 17267 37247
rect 17693 37213 17727 37247
rect 18153 37213 18187 37247
rect 18521 37213 18555 37247
rect 20637 37213 20671 37247
rect 20729 37213 20763 37247
rect 20913 37213 20947 37247
rect 22201 37213 22235 37247
rect 22569 37213 22603 37247
rect 22753 37213 22787 37247
rect 22845 37213 22879 37247
rect 9864 37145 9898 37179
rect 11336 37145 11370 37179
rect 12808 37145 12842 37179
rect 18061 37145 18095 37179
rect 20370 37145 20404 37179
rect 8723 37077 8757 37111
rect 12449 37077 12483 37111
rect 13921 37077 13955 37111
rect 16221 37077 16255 37111
rect 16957 37077 16991 37111
rect 17969 37077 18003 37111
rect 19257 37077 19291 37111
rect 21097 37077 21131 37111
rect 21649 37077 21683 37111
rect 23029 37077 23063 37111
rect 8033 36873 8067 36907
rect 12817 36873 12851 36907
rect 13921 36873 13955 36907
rect 15761 36873 15795 36907
rect 18061 36873 18095 36907
rect 21925 36873 21959 36907
rect 23397 36873 23431 36907
rect 9036 36805 9070 36839
rect 18245 36805 18279 36839
rect 23038 36805 23072 36839
rect 7481 36737 7515 36771
rect 8769 36737 8803 36771
rect 10425 36737 10459 36771
rect 12449 36737 12483 36771
rect 12909 36737 12943 36771
rect 13001 36737 13035 36771
rect 15577 36737 15611 36771
rect 16681 36737 16715 36771
rect 16937 36737 16971 36771
rect 19993 36737 20027 36771
rect 20269 36737 20303 36771
rect 21189 36737 21223 36771
rect 21373 36737 21407 36771
rect 21557 36737 21591 36771
rect 23305 36737 23339 36771
rect 24510 36737 24544 36771
rect 24777 36737 24811 36771
rect 8585 36669 8619 36703
rect 10609 36669 10643 36703
rect 10793 36669 10827 36703
rect 12541 36669 12575 36703
rect 12633 36669 12667 36703
rect 13277 36669 13311 36703
rect 14013 36669 14047 36703
rect 15945 36669 15979 36703
rect 16497 36669 16531 36703
rect 20545 36669 20579 36703
rect 10149 36601 10183 36635
rect 7665 36533 7699 36567
rect 10241 36533 10275 36567
rect 11345 36533 11379 36567
rect 11805 36533 11839 36567
rect 13185 36533 13219 36567
rect 14657 36533 14691 36567
rect 20085 36533 20119 36567
rect 21097 36533 21131 36567
rect 7941 36329 7975 36363
rect 10977 36329 11011 36363
rect 12265 36329 12299 36363
rect 13093 36329 13127 36363
rect 16773 36329 16807 36363
rect 19073 36329 19107 36363
rect 12357 36261 12391 36295
rect 15485 36261 15519 36295
rect 19257 36261 19291 36295
rect 20729 36261 20763 36295
rect 9137 36193 9171 36227
rect 10793 36193 10827 36227
rect 11529 36193 11563 36227
rect 11713 36193 11747 36227
rect 12725 36193 12759 36227
rect 13277 36193 13311 36227
rect 15853 36193 15887 36227
rect 18061 36193 18095 36227
rect 20821 36193 20855 36227
rect 1409 36125 1443 36159
rect 7849 36125 7883 36159
rect 10149 36125 10183 36159
rect 11897 36125 11931 36159
rect 11989 36125 12023 36159
rect 12541 36125 12575 36159
rect 12909 36125 12943 36159
rect 13185 36125 13219 36159
rect 13369 36125 13403 36159
rect 14105 36125 14139 36159
rect 14372 36125 14406 36159
rect 16037 36125 16071 36159
rect 16405 36125 16439 36159
rect 16497 36125 16531 36159
rect 17049 36125 17083 36159
rect 17141 36125 17175 36159
rect 17233 36125 17267 36159
rect 17417 36125 17451 36159
rect 17693 36125 17727 36159
rect 17785 36125 17819 36159
rect 18705 36125 18739 36159
rect 18889 36125 18923 36159
rect 19901 36125 19935 36159
rect 20085 36125 20119 36159
rect 20269 36125 20303 36159
rect 20361 36125 20395 36159
rect 20453 36125 20487 36159
rect 23765 36125 23799 36159
rect 10241 36057 10275 36091
rect 12081 36057 12115 36091
rect 17969 36057 18003 36091
rect 21088 36057 21122 36091
rect 23520 36057 23554 36091
rect 9781 35989 9815 36023
rect 9965 35989 9999 36023
rect 13645 35989 13679 36023
rect 16221 35989 16255 36023
rect 16681 35989 16715 36023
rect 22201 35989 22235 36023
rect 22385 35989 22419 36023
rect 8953 35785 8987 35819
rect 10977 35785 11011 35819
rect 13277 35785 13311 35819
rect 19073 35785 19107 35819
rect 20545 35785 20579 35819
rect 21373 35785 21407 35819
rect 21833 35785 21867 35819
rect 23857 35785 23891 35819
rect 24317 35785 24351 35819
rect 9413 35717 9447 35751
rect 12173 35717 12207 35751
rect 16773 35717 16807 35751
rect 19432 35717 19466 35751
rect 8769 35649 8803 35683
rect 9853 35649 9887 35683
rect 11161 35649 11195 35683
rect 11897 35649 11931 35683
rect 12357 35649 12391 35683
rect 12633 35649 12667 35683
rect 12817 35649 12851 35683
rect 12909 35649 12943 35683
rect 13001 35649 13035 35683
rect 14473 35649 14507 35683
rect 14565 35649 14599 35683
rect 15108 35649 15142 35683
rect 17417 35649 17451 35683
rect 17693 35649 17727 35683
rect 17949 35649 17983 35683
rect 19165 35649 19199 35683
rect 20637 35649 20671 35683
rect 21557 35649 21591 35683
rect 22109 35649 22143 35683
rect 22201 35649 22235 35683
rect 22385 35649 22419 35683
rect 22569 35649 22603 35683
rect 23581 35649 23615 35683
rect 23765 35649 23799 35683
rect 24041 35649 24075 35683
rect 24133 35649 24167 35683
rect 9597 35581 9631 35615
rect 12541 35581 12575 35615
rect 13921 35581 13955 35615
rect 14841 35581 14875 35615
rect 22661 35581 22695 35615
rect 23305 35581 23339 35615
rect 23397 35581 23431 35615
rect 11805 35513 11839 35547
rect 17049 35513 17083 35547
rect 17601 35513 17635 35547
rect 22293 35513 22327 35547
rect 9321 35445 9355 35479
rect 11345 35445 11379 35479
rect 13369 35445 13403 35479
rect 14749 35445 14783 35479
rect 16221 35445 16255 35479
rect 17233 35445 17267 35479
rect 21281 35445 21315 35479
rect 10885 35241 10919 35275
rect 12449 35241 12483 35275
rect 19073 35241 19107 35275
rect 20269 35241 20303 35275
rect 21741 35241 21775 35275
rect 23857 35241 23891 35275
rect 10793 35173 10827 35207
rect 14105 35173 14139 35207
rect 15945 35173 15979 35207
rect 17049 35173 17083 35207
rect 19717 35173 19751 35207
rect 9413 35105 9447 35139
rect 12081 35105 12115 35139
rect 14565 35105 14599 35139
rect 16037 35105 16071 35139
rect 17141 35105 17175 35139
rect 18613 35105 18647 35139
rect 22017 35105 22051 35139
rect 22293 35105 22327 35139
rect 22385 35105 22419 35139
rect 9680 35037 9714 35071
rect 11069 35037 11103 35071
rect 11253 35037 11287 35071
rect 11345 35037 11379 35071
rect 11621 35037 11655 35071
rect 12265 35037 12299 35071
rect 13921 35037 13955 35071
rect 14289 35037 14323 35071
rect 16221 35037 16255 35071
rect 16405 35037 16439 35071
rect 16773 35037 16807 35071
rect 16865 35037 16899 35071
rect 17785 35037 17819 35071
rect 18429 35037 18463 35071
rect 18521 35037 18555 35071
rect 18797 35037 18831 35071
rect 18889 35037 18923 35071
rect 19901 35037 19935 35071
rect 21649 35037 21683 35071
rect 21925 35037 21959 35071
rect 22569 35037 22603 35071
rect 23581 35037 23615 35071
rect 23673 35037 23707 35071
rect 34529 35037 34563 35071
rect 13676 34969 13710 35003
rect 14832 34969 14866 35003
rect 21382 34969 21416 35003
rect 11529 34901 11563 34935
rect 11805 34901 11839 34935
rect 12541 34901 12575 34935
rect 16589 34901 16623 34935
rect 22201 34901 22235 34935
rect 22753 34901 22787 34935
rect 34345 34901 34379 34935
rect 9505 34697 9539 34731
rect 10149 34697 10183 34731
rect 11345 34697 11379 34731
rect 13369 34697 13403 34731
rect 15025 34697 15059 34731
rect 16037 34697 16071 34731
rect 16405 34697 16439 34731
rect 17233 34697 17267 34731
rect 17601 34697 17635 34731
rect 20637 34697 20671 34731
rect 23397 34697 23431 34731
rect 13553 34629 13587 34663
rect 18714 34629 18748 34663
rect 22385 34629 22419 34663
rect 9137 34561 9171 34595
rect 9229 34561 9263 34595
rect 9689 34561 9723 34595
rect 9965 34561 9999 34595
rect 10977 34561 11011 34595
rect 11161 34561 11195 34595
rect 11621 34561 11655 34595
rect 12256 34561 12290 34595
rect 14381 34561 14415 34595
rect 15209 34561 15243 34595
rect 16221 34561 16255 34595
rect 16313 34561 16347 34595
rect 16497 34561 16531 34595
rect 18981 34561 19015 34595
rect 19257 34561 19291 34595
rect 19524 34561 19558 34595
rect 20729 34561 20763 34595
rect 22201 34561 22235 34595
rect 24510 34561 24544 34595
rect 25421 34561 25455 34595
rect 9781 34493 9815 34527
rect 10241 34493 10275 34527
rect 10793 34493 10827 34527
rect 11989 34493 12023 34527
rect 15853 34493 15887 34527
rect 16773 34493 16807 34527
rect 22017 34493 22051 34527
rect 22477 34493 22511 34527
rect 23029 34493 23063 34527
rect 24777 34493 24811 34527
rect 13829 34425 13863 34459
rect 17141 34425 17175 34459
rect 8953 34357 8987 34391
rect 11805 34357 11839 34391
rect 14289 34357 14323 34391
rect 15301 34357 15335 34391
rect 21373 34357 21407 34391
rect 24869 34357 24903 34391
rect 8953 34153 8987 34187
rect 9689 34153 9723 34187
rect 13737 34153 13771 34187
rect 14105 34153 14139 34187
rect 17693 34153 17727 34187
rect 18705 34153 18739 34187
rect 13001 34085 13035 34119
rect 13277 34085 13311 34119
rect 13553 34085 13587 34119
rect 9505 34017 9539 34051
rect 9781 34017 9815 34051
rect 13461 34017 13495 34051
rect 24777 34017 24811 34051
rect 8493 33949 8527 33983
rect 8585 33949 8619 33983
rect 9965 33949 9999 33983
rect 12449 33949 12483 33983
rect 12541 33949 12575 33983
rect 13185 33949 13219 33983
rect 14749 33949 14783 33983
rect 15016 33949 15050 33983
rect 16865 33949 16899 33983
rect 17969 33949 18003 33983
rect 18061 33949 18095 33983
rect 18153 33949 18187 33983
rect 18337 33949 18371 33983
rect 19809 33949 19843 33983
rect 20453 33949 20487 33983
rect 20729 33949 20763 33983
rect 20913 33949 20947 33983
rect 22385 33949 22419 33983
rect 22477 33949 22511 33983
rect 24133 33949 24167 33983
rect 24409 33949 24443 33983
rect 24593 33949 24627 33983
rect 9689 33881 9723 33915
rect 10425 33881 10459 33915
rect 12817 33881 12851 33915
rect 13461 33881 13495 33915
rect 13921 33881 13955 33915
rect 14289 33881 14323 33915
rect 14473 33881 14507 33915
rect 18797 33881 18831 33915
rect 22140 33881 22174 33915
rect 22744 33881 22778 33915
rect 8309 33813 8343 33847
rect 8769 33813 8803 33847
rect 10149 33813 10183 33847
rect 11897 33813 11931 33847
rect 12265 33813 12299 33847
rect 13721 33813 13755 33847
rect 16129 33813 16163 33847
rect 16681 33813 16715 33847
rect 20545 33813 20579 33847
rect 21005 33813 21039 33847
rect 23857 33813 23891 33847
rect 23949 33813 23983 33847
rect 8953 33609 8987 33643
rect 11161 33609 11195 33643
rect 15485 33609 15519 33643
rect 17785 33609 17819 33643
rect 22661 33609 22695 33643
rect 24593 33609 24627 33643
rect 7656 33541 7690 33575
rect 10824 33541 10858 33575
rect 17049 33541 17083 33575
rect 19555 33541 19589 33575
rect 20361 33541 20395 33575
rect 23796 33541 23830 33575
rect 11345 33473 11379 33507
rect 12642 33473 12676 33507
rect 12909 33473 12943 33507
rect 14565 33473 14599 33507
rect 14749 33473 14783 33507
rect 14841 33473 14875 33507
rect 15025 33473 15059 33507
rect 15117 33473 15151 33507
rect 15209 33473 15243 33507
rect 15577 33473 15611 33507
rect 15945 33473 15979 33507
rect 16129 33473 16163 33507
rect 16681 33473 16715 33507
rect 16865 33473 16899 33507
rect 16957 33473 16991 33507
rect 17141 33473 17175 33507
rect 18061 33473 18095 33507
rect 18981 33473 19015 33507
rect 19257 33473 19291 33507
rect 20177 33473 20211 33507
rect 20453 33473 20487 33507
rect 20637 33473 20671 33507
rect 20913 33473 20947 33507
rect 21833 33473 21867 33507
rect 24041 33473 24075 33507
rect 24225 33473 24259 33507
rect 24317 33473 24351 33507
rect 24501 33473 24535 33507
rect 24777 33473 24811 33507
rect 7389 33405 7423 33439
rect 9597 33405 9631 33439
rect 11069 33405 11103 33439
rect 13645 33405 13679 33439
rect 14473 33405 14507 33439
rect 14657 33405 14691 33439
rect 15853 33405 15887 33439
rect 17785 33405 17819 33439
rect 19441 33405 19475 33439
rect 19717 33405 19751 33439
rect 20085 33405 20119 33439
rect 9689 33337 9723 33371
rect 15669 33337 15703 33371
rect 16037 33337 16071 33371
rect 19165 33337 19199 33371
rect 19349 33337 19383 33371
rect 19625 33337 19659 33371
rect 20821 33337 20855 33371
rect 22477 33337 22511 33371
rect 8769 33269 8803 33303
rect 11529 33269 11563 33303
rect 13093 33269 13127 33303
rect 13829 33269 13863 33303
rect 15761 33269 15795 33303
rect 16865 33269 16899 33303
rect 17969 33269 18003 33303
rect 20453 33269 20487 33303
rect 8033 33065 8067 33099
rect 10333 33065 10367 33099
rect 12265 33065 12299 33099
rect 15025 33065 15059 33099
rect 16129 33065 16163 33099
rect 17049 33065 17083 33099
rect 19257 33065 19291 33099
rect 20545 33065 20579 33099
rect 21097 33065 21131 33099
rect 22293 33065 22327 33099
rect 24685 33065 24719 33099
rect 13921 32997 13955 33031
rect 18153 32997 18187 33031
rect 22201 32997 22235 33031
rect 7665 32929 7699 32963
rect 8125 32929 8159 32963
rect 14749 32929 14783 32963
rect 15393 32929 15427 32963
rect 17233 32929 17267 32963
rect 18889 32929 18923 32963
rect 21833 32929 21867 32963
rect 23397 32929 23431 32963
rect 7849 32861 7883 32895
rect 8769 32861 8803 32895
rect 8953 32861 8987 32895
rect 9220 32861 9254 32895
rect 10517 32861 10551 32895
rect 11345 32861 11379 32895
rect 11621 32861 11655 32895
rect 12541 32861 12575 32895
rect 12808 32861 12842 32895
rect 14105 32861 14139 32895
rect 14657 32861 14691 32895
rect 15301 32861 15335 32895
rect 15945 32861 15979 32895
rect 16313 32861 16347 32895
rect 17325 32861 17359 32895
rect 17693 32861 17727 32895
rect 17785 32861 17819 32895
rect 17877 32861 17911 32895
rect 17969 32861 18003 32895
rect 18337 32861 18371 32895
rect 19441 32861 19475 32895
rect 19533 32861 19567 32895
rect 19717 32861 19751 32895
rect 19901 32861 19935 32895
rect 20361 32861 20395 32895
rect 20637 32861 20671 32895
rect 21189 32861 21223 32895
rect 21373 32861 21407 32895
rect 22017 32861 22051 32895
rect 22477 32861 22511 32895
rect 23121 32861 23155 32895
rect 23213 32861 23247 32895
rect 24041 32861 24075 32895
rect 24593 32861 24627 32895
rect 25329 32861 25363 32895
rect 15761 32793 15795 32827
rect 20729 32793 20763 32827
rect 20913 32793 20947 32827
rect 21281 32793 21315 32827
rect 11161 32725 11195 32759
rect 11529 32725 11563 32759
rect 14657 32725 14691 32759
rect 16405 32725 16439 32759
rect 20085 32725 20119 32759
rect 20177 32725 20211 32759
rect 23489 32725 23523 32759
rect 24409 32725 24443 32759
rect 7665 32521 7699 32555
rect 10241 32521 10275 32555
rect 13369 32521 13403 32555
rect 14197 32521 14231 32555
rect 14841 32521 14875 32555
rect 15761 32521 15795 32555
rect 18337 32521 18371 32555
rect 19901 32521 19935 32555
rect 23673 32521 23707 32555
rect 23857 32521 23891 32555
rect 25421 32521 25455 32555
rect 25513 32521 25547 32555
rect 9045 32453 9079 32487
rect 9781 32453 9815 32487
rect 10333 32453 10367 32487
rect 14473 32453 14507 32487
rect 17509 32453 17543 32487
rect 23305 32453 23339 32487
rect 24308 32453 24342 32487
rect 7389 32385 7423 32419
rect 7849 32385 7883 32419
rect 7941 32385 7975 32419
rect 8033 32385 8067 32419
rect 9321 32385 9355 32419
rect 9413 32385 9447 32419
rect 9505 32385 9539 32419
rect 9689 32385 9723 32419
rect 9965 32385 9999 32419
rect 10057 32385 10091 32419
rect 10425 32385 10459 32419
rect 10793 32385 10827 32419
rect 10885 32385 10919 32419
rect 11253 32385 11287 32419
rect 12642 32385 12676 32419
rect 13645 32385 13679 32419
rect 13737 32385 13771 32419
rect 13829 32385 13863 32419
rect 14013 32385 14047 32419
rect 14105 32385 14139 32419
rect 14381 32385 14415 32419
rect 14657 32385 14691 32419
rect 14749 32385 14783 32419
rect 14841 32385 14875 32419
rect 15025 32385 15059 32419
rect 15577 32385 15611 32419
rect 15669 32385 15703 32419
rect 15945 32385 15979 32419
rect 16037 32385 16071 32419
rect 16221 32385 16255 32419
rect 16681 32385 16715 32419
rect 16773 32385 16807 32419
rect 16957 32385 16991 32419
rect 17233 32385 17267 32419
rect 17325 32385 17359 32419
rect 17877 32385 17911 32419
rect 18705 32385 18739 32419
rect 18981 32385 19015 32419
rect 19073 32385 19107 32419
rect 19349 32385 19383 32419
rect 19533 32385 19567 32419
rect 19671 32385 19705 32419
rect 19809 32385 19843 32419
rect 20269 32385 20303 32419
rect 20545 32385 20579 32419
rect 22845 32385 22879 32419
rect 22937 32385 22971 32419
rect 23029 32385 23063 32419
rect 23213 32385 23247 32419
rect 23581 32385 23615 32419
rect 24041 32385 24075 32419
rect 8401 32317 8435 32351
rect 11069 32317 11103 32351
rect 12909 32317 12943 32351
rect 15393 32317 15427 32351
rect 16129 32317 16163 32351
rect 17509 32317 17543 32351
rect 17785 32317 17819 32351
rect 18245 32317 18279 32351
rect 18613 32317 18647 32351
rect 19257 32317 19291 32351
rect 20177 32317 20211 32351
rect 21097 32317 21131 32351
rect 21925 32317 21959 32351
rect 22569 32317 22603 32351
rect 23489 32317 23523 32351
rect 23949 32317 23983 32351
rect 26065 32317 26099 32351
rect 7573 32249 7607 32283
rect 8217 32249 8251 32283
rect 11529 32249 11563 32283
rect 15485 32249 15519 32283
rect 19165 32249 19199 32283
rect 8953 32181 8987 32215
rect 10517 32181 10551 32215
rect 10977 32181 11011 32215
rect 14381 32181 14415 32215
rect 14473 32181 14507 32215
rect 17141 32181 17175 32215
rect 17601 32181 17635 32215
rect 19441 32181 19475 32215
rect 22477 32181 22511 32215
rect 8769 31977 8803 32011
rect 12265 31977 12299 32011
rect 15853 31977 15887 32011
rect 21373 31977 21407 32011
rect 22937 31977 22971 32011
rect 23397 31977 23431 32011
rect 23489 31977 23523 32011
rect 24225 31977 24259 32011
rect 25789 31977 25823 32011
rect 10333 31909 10367 31943
rect 14565 31909 14599 31943
rect 17233 31909 17267 31943
rect 17969 31909 18003 31943
rect 21465 31909 21499 31943
rect 23305 31909 23339 31943
rect 23765 31909 23799 31943
rect 7389 31841 7423 31875
rect 12909 31841 12943 31875
rect 13829 31841 13863 31875
rect 16221 31841 16255 31875
rect 18521 31841 18555 31875
rect 19809 31841 19843 31875
rect 22845 31841 22879 31875
rect 24409 31841 24443 31875
rect 8953 31773 8987 31807
rect 9220 31773 9254 31807
rect 10885 31773 10919 31807
rect 14381 31773 14415 31807
rect 16129 31773 16163 31807
rect 16681 31773 16715 31807
rect 16865 31773 16899 31807
rect 17049 31773 17083 31807
rect 17509 31773 17543 31807
rect 17693 31773 17727 31807
rect 17785 31773 17819 31807
rect 18705 31773 18739 31807
rect 18889 31773 18923 31807
rect 18981 31773 19015 31807
rect 19533 31773 19567 31807
rect 19717 31773 19751 31807
rect 19901 31773 19935 31807
rect 20085 31773 20119 31807
rect 20269 31773 20303 31807
rect 20361 31773 20395 31807
rect 21189 31773 21223 31807
rect 23213 31773 23247 31807
rect 23673 31773 23707 31807
rect 23949 31773 23983 31807
rect 24041 31773 24075 31807
rect 24225 31773 24259 31807
rect 7656 31705 7690 31739
rect 11152 31705 11186 31739
rect 16957 31705 16991 31739
rect 22578 31705 22612 31739
rect 24654 31705 24688 31739
rect 12357 31637 12391 31671
rect 13277 31637 13311 31671
rect 17601 31637 17635 31671
rect 21005 31637 21039 31671
rect 8033 31433 8067 31467
rect 9505 31433 9539 31467
rect 14197 31433 14231 31467
rect 17141 31433 17175 31467
rect 19901 31433 19935 31467
rect 23213 31433 23247 31467
rect 23857 31433 23891 31467
rect 23949 31433 23983 31467
rect 24225 31433 24259 31467
rect 24317 31433 24351 31467
rect 12992 31365 13026 31399
rect 15485 31365 15519 31399
rect 21014 31365 21048 31399
rect 22100 31365 22134 31399
rect 8217 31297 8251 31331
rect 8309 31297 8343 31331
rect 8493 31297 8527 31331
rect 8677 31297 8711 31331
rect 8769 31297 8803 31331
rect 9689 31297 9723 31331
rect 10241 31297 10275 31331
rect 11529 31297 11563 31331
rect 11713 31297 11747 31331
rect 11805 31297 11839 31331
rect 11897 31297 11931 31331
rect 12357 31297 12391 31331
rect 12449 31297 12483 31331
rect 14381 31297 14415 31331
rect 14657 31297 14691 31331
rect 14841 31297 14875 31331
rect 15301 31297 15335 31331
rect 15761 31297 15795 31331
rect 15853 31297 15887 31331
rect 16037 31297 16071 31331
rect 17325 31297 17359 31331
rect 17601 31297 17635 31331
rect 17785 31297 17819 31331
rect 17877 31297 17911 31331
rect 17969 31297 18003 31331
rect 18153 31297 18187 31331
rect 21281 31297 21315 31331
rect 21833 31297 21867 31331
rect 23673 31297 23707 31331
rect 24133 31297 24167 31331
rect 24869 31297 24903 31331
rect 9413 31229 9447 31263
rect 9873 31229 9907 31263
rect 10517 31229 10551 31263
rect 12725 31229 12759 31263
rect 14565 31229 14599 31263
rect 18337 31229 18371 31263
rect 18429 31229 18463 31263
rect 24501 31229 24535 31263
rect 10057 31093 10091 31127
rect 11161 31093 11195 31127
rect 12173 31093 12207 31127
rect 12633 31093 12667 31127
rect 14105 31093 14139 31127
rect 15117 31093 15151 31127
rect 15669 31093 15703 31127
rect 16037 31093 16071 31127
rect 19073 31093 19107 31127
rect 25513 31093 25547 31127
rect 8217 30889 8251 30923
rect 10333 30889 10367 30923
rect 13829 30889 13863 30923
rect 17233 30889 17267 30923
rect 17693 30889 17727 30923
rect 20729 30889 20763 30923
rect 22661 30889 22695 30923
rect 24593 30889 24627 30923
rect 22109 30821 22143 30855
rect 12173 30753 12207 30787
rect 19073 30753 19107 30787
rect 23029 30753 23063 30787
rect 24961 30753 24995 30787
rect 6837 30685 6871 30719
rect 8953 30685 8987 30719
rect 12817 30685 12851 30719
rect 14289 30685 14323 30719
rect 14381 30685 14415 30719
rect 14657 30685 14691 30719
rect 14749 30685 14783 30719
rect 15117 30685 15151 30719
rect 15853 30685 15887 30719
rect 17601 30685 17635 30719
rect 18817 30685 18851 30719
rect 19349 30685 19383 30719
rect 19625 30685 19659 30719
rect 19717 30685 19751 30719
rect 19993 30685 20027 30719
rect 20177 30685 20211 30719
rect 20269 30685 20303 30719
rect 20361 30685 20395 30719
rect 20545 30685 20579 30719
rect 22845 30685 22879 30719
rect 23305 30685 23339 30719
rect 24777 30685 24811 30719
rect 7082 30617 7116 30651
rect 9220 30617 9254 30651
rect 10425 30617 10459 30651
rect 13553 30617 13587 30651
rect 14565 30617 14599 30651
rect 16098 30617 16132 30651
rect 19533 30617 19567 30651
rect 20821 30617 20855 30651
rect 12265 30549 12299 30583
rect 14105 30549 14139 30583
rect 14933 30549 14967 30583
rect 15761 30549 15795 30583
rect 17509 30549 17543 30583
rect 19901 30549 19935 30583
rect 23949 30549 23983 30583
rect 14841 30345 14875 30379
rect 19717 30345 19751 30379
rect 20545 30345 20579 30379
rect 24685 30345 24719 30379
rect 9505 30277 9539 30311
rect 9864 30277 9898 30311
rect 12164 30277 12198 30311
rect 18245 30277 18279 30311
rect 18337 30277 18371 30311
rect 22109 30277 22143 30311
rect 6561 30209 6595 30243
rect 8125 30209 8159 30243
rect 9321 30209 9355 30243
rect 11529 30209 11563 30243
rect 11897 30209 11931 30243
rect 13737 30209 13771 30243
rect 15117 30209 15151 30243
rect 15209 30209 15243 30243
rect 15301 30209 15335 30243
rect 15485 30209 15519 30243
rect 15577 30209 15611 30243
rect 16773 30209 16807 30243
rect 16957 30209 16991 30243
rect 17049 30209 17083 30243
rect 17233 30209 17267 30243
rect 17325 30209 17359 30243
rect 17417 30209 17451 30243
rect 17601 30209 17635 30243
rect 17785 30209 17819 30243
rect 17969 30209 18003 30243
rect 18117 30209 18151 30243
rect 18475 30209 18509 30243
rect 18705 30209 18739 30243
rect 18889 30209 18923 30243
rect 18981 30209 19015 30243
rect 19165 30209 19199 30243
rect 19257 30209 19291 30243
rect 19533 30209 19567 30243
rect 19993 30209 20027 30243
rect 20085 30209 20119 30243
rect 20269 30209 20303 30243
rect 20637 30209 20671 30243
rect 21833 30209 21867 30243
rect 23305 30209 23339 30243
rect 23572 30209 23606 30243
rect 9137 30141 9171 30175
rect 9597 30141 9631 30175
rect 14013 30141 14047 30175
rect 14105 30141 14139 30175
rect 19349 30141 19383 30175
rect 6745 30073 6779 30107
rect 13553 30073 13587 30107
rect 18613 30073 18647 30107
rect 22385 30073 22419 30107
rect 7941 30005 7975 30039
rect 10977 30005 11011 30039
rect 11713 30005 11747 30039
rect 13277 30005 13311 30039
rect 13921 30005 13955 30039
rect 14749 30005 14783 30039
rect 15761 30005 15795 30039
rect 16957 30005 16991 30039
rect 18889 30005 18923 30039
rect 20269 30005 20303 30039
rect 22017 30005 22051 30039
rect 22569 30005 22603 30039
rect 6285 29801 6319 29835
rect 10517 29801 10551 29835
rect 15485 29801 15519 29835
rect 16129 29801 16163 29835
rect 18429 29801 18463 29835
rect 18981 29801 19015 29835
rect 19257 29801 19291 29835
rect 19441 29801 19475 29835
rect 20729 29801 20763 29835
rect 23397 29801 23431 29835
rect 23857 29801 23891 29835
rect 21741 29733 21775 29767
rect 5917 29665 5951 29699
rect 14105 29665 14139 29699
rect 6101 29597 6135 29631
rect 7389 29597 7423 29631
rect 7656 29597 7690 29631
rect 9505 29597 9539 29631
rect 10149 29597 10183 29631
rect 10241 29597 10275 29631
rect 10425 29597 10459 29631
rect 10701 29597 10735 29631
rect 11917 29597 11951 29631
rect 12173 29597 12207 29631
rect 12265 29597 12299 29631
rect 13093 29597 13127 29631
rect 14372 29597 14406 29631
rect 15577 29597 15611 29631
rect 15761 29597 15795 29631
rect 15853 29597 15887 29631
rect 15945 29597 15979 29631
rect 18521 29597 18555 29631
rect 18705 29597 18739 29631
rect 19073 29597 19107 29631
rect 20453 29597 20487 29631
rect 20637 29597 20671 29631
rect 20913 29597 20947 29631
rect 21097 29597 21131 29631
rect 21373 29597 21407 29631
rect 21925 29597 21959 29631
rect 23581 29597 23615 29631
rect 23765 29597 23799 29631
rect 24041 29597 24075 29631
rect 13461 29529 13495 29563
rect 17969 29529 18003 29563
rect 18061 29529 18095 29563
rect 18245 29529 18279 29563
rect 19625 29529 19659 29563
rect 22170 29529 22204 29563
rect 8769 29461 8803 29495
rect 8953 29461 8987 29495
rect 10793 29461 10827 29495
rect 12909 29461 12943 29495
rect 16681 29461 16715 29495
rect 18613 29461 18647 29495
rect 19415 29461 19449 29495
rect 19901 29461 19935 29495
rect 21281 29461 21315 29495
rect 21833 29461 21867 29495
rect 23305 29461 23339 29495
rect 1593 29257 1627 29291
rect 8033 29257 8067 29291
rect 9413 29257 9447 29291
rect 9873 29257 9907 29291
rect 11345 29257 11379 29291
rect 13921 29257 13955 29291
rect 14197 29257 14231 29291
rect 14473 29257 14507 29291
rect 16497 29257 16531 29291
rect 17969 29257 18003 29291
rect 19165 29257 19199 29291
rect 21005 29257 21039 29291
rect 24133 29257 24167 29291
rect 9597 29189 9631 29223
rect 10885 29189 10919 29223
rect 12265 29189 12299 29223
rect 14657 29189 14691 29223
rect 14857 29189 14891 29223
rect 15945 29189 15979 29223
rect 17233 29189 17267 29223
rect 17449 29189 17483 29223
rect 1409 29121 1443 29155
rect 6009 29121 6043 29155
rect 6561 29121 6595 29155
rect 6817 29121 6851 29155
rect 8217 29121 8251 29155
rect 8401 29121 8435 29155
rect 9505 29121 9539 29155
rect 10057 29121 10091 29155
rect 10149 29121 10183 29155
rect 10609 29121 10643 29155
rect 11161 29121 11195 29155
rect 13093 29121 13127 29155
rect 13185 29121 13219 29155
rect 14013 29121 14047 29155
rect 14289 29121 14323 29155
rect 14381 29121 14415 29155
rect 15117 29121 15151 29155
rect 16037 29121 16071 29155
rect 16313 29121 16347 29155
rect 16865 29121 16899 29155
rect 17049 29121 17083 29155
rect 17693 29121 17727 29155
rect 18337 29121 18371 29155
rect 18797 29121 18831 29155
rect 19349 29121 19383 29155
rect 19441 29121 19475 29155
rect 19625 29121 19659 29155
rect 19892 29121 19926 29155
rect 21097 29121 21131 29155
rect 21833 29121 21867 29155
rect 22089 29121 22123 29155
rect 23489 29121 23523 29155
rect 23765 29121 23799 29155
rect 23949 29121 23983 29155
rect 24225 29121 24259 29155
rect 24409 29121 24443 29155
rect 5825 29053 5859 29087
rect 9045 29053 9079 29087
rect 9229 29053 9263 29087
rect 10977 29053 11011 29087
rect 12081 29053 12115 29087
rect 16129 29053 16163 29087
rect 17141 29053 17175 29087
rect 17969 29053 18003 29087
rect 18061 29053 18095 29087
rect 19073 29053 19107 29087
rect 23673 29053 23707 29087
rect 7941 28985 7975 29019
rect 9781 28985 9815 29019
rect 10333 28985 10367 29019
rect 12541 28985 12575 29019
rect 15761 28985 15795 29019
rect 17785 28985 17819 29019
rect 18153 28985 18187 29019
rect 18521 28985 18555 29019
rect 18981 28985 19015 29019
rect 21281 28985 21315 29019
rect 23213 28985 23247 29019
rect 6193 28917 6227 28951
rect 8493 28917 8527 28951
rect 10425 28917 10459 28951
rect 10517 28917 10551 28951
rect 11529 28917 11563 28951
rect 12725 28917 12759 28951
rect 12909 28917 12943 28951
rect 14841 28917 14875 28951
rect 15025 28917 15059 28951
rect 16681 28917 16715 28951
rect 17417 28917 17451 28951
rect 17601 28917 17635 28951
rect 18613 28917 18647 28951
rect 23305 28917 23339 28951
rect 24225 28917 24259 28951
rect 6561 28713 6595 28747
rect 8309 28713 8343 28747
rect 8769 28713 8803 28747
rect 10793 28713 10827 28747
rect 13185 28713 13219 28747
rect 14289 28713 14323 28747
rect 15945 28713 15979 28747
rect 17601 28713 17635 28747
rect 19441 28713 19475 28747
rect 20177 28713 20211 28747
rect 20545 28713 20579 28747
rect 22753 28713 22787 28747
rect 23029 28713 23063 28747
rect 10885 28645 10919 28679
rect 16681 28645 16715 28679
rect 7757 28577 7791 28611
rect 8677 28577 8711 28611
rect 9597 28577 9631 28611
rect 11805 28577 11839 28611
rect 13369 28577 13403 28611
rect 15669 28577 15703 28611
rect 18245 28577 18279 28611
rect 18981 28577 19015 28611
rect 20085 28577 20119 28611
rect 20729 28577 20763 28611
rect 21281 28577 21315 28611
rect 6377 28509 6411 28543
rect 7573 28509 7607 28543
rect 8033 28509 8067 28543
rect 8217 28509 8251 28543
rect 8493 28509 8527 28543
rect 9781 28509 9815 28543
rect 10149 28509 10183 28543
rect 10241 28509 10275 28543
rect 10517 28509 10551 28543
rect 10609 28509 10643 28543
rect 11437 28509 11471 28543
rect 13277 28509 13311 28543
rect 13553 28509 13587 28543
rect 13645 28509 13679 28543
rect 15761 28509 15795 28543
rect 15945 28509 15979 28543
rect 16037 28509 16071 28543
rect 16773 28509 16807 28543
rect 20361 28509 20395 28543
rect 20637 28509 20671 28543
rect 22477 28509 22511 28543
rect 22569 28509 22603 28543
rect 22845 28509 22879 28543
rect 22937 28509 22971 28543
rect 23213 28509 23247 28543
rect 23305 28509 23339 28543
rect 8769 28441 8803 28475
rect 12050 28441 12084 28475
rect 15402 28441 15436 28475
rect 7389 28373 7423 28407
rect 7849 28373 7883 28407
rect 9045 28373 9079 28407
rect 9965 28373 9999 28407
rect 10425 28373 10459 28407
rect 13829 28373 13863 28407
rect 17417 28373 17451 28407
rect 18429 28373 18463 28407
rect 22293 28373 22327 28407
rect 23489 28373 23523 28407
rect 7481 28169 7515 28203
rect 9045 28169 9079 28203
rect 11253 28169 11287 28203
rect 11529 28169 11563 28203
rect 12633 28169 12667 28203
rect 13461 28169 13495 28203
rect 15485 28169 15519 28203
rect 18061 28169 18095 28203
rect 19717 28169 19751 28203
rect 7818 28101 7852 28135
rect 10118 28101 10152 28135
rect 12173 28101 12207 28135
rect 21265 28101 21299 28135
rect 21465 28101 21499 28135
rect 22201 28101 22235 28135
rect 7021 28033 7055 28067
rect 7297 28033 7331 28067
rect 9597 28033 9631 28067
rect 11713 28033 11747 28067
rect 11805 28033 11839 28067
rect 12725 28033 12759 28067
rect 13001 28033 13035 28067
rect 13093 28033 13127 28067
rect 13369 28033 13403 28067
rect 13553 28033 13587 28067
rect 13921 28033 13955 28067
rect 14188 28033 14222 28067
rect 16221 28033 16255 28067
rect 16313 28033 16347 28067
rect 16948 28033 16982 28067
rect 18337 28033 18371 28067
rect 18593 28033 18627 28067
rect 20361 28033 20395 28067
rect 22017 28033 22051 28067
rect 7573 27965 7607 27999
rect 9873 27965 9907 27999
rect 12817 27965 12851 27999
rect 16129 27965 16163 27999
rect 16497 27965 16531 27999
rect 16681 27965 16715 27999
rect 8953 27897 8987 27931
rect 12449 27897 12483 27931
rect 16221 27897 16255 27931
rect 7205 27829 7239 27863
rect 13277 27829 13311 27863
rect 15301 27829 15335 27863
rect 19809 27829 19843 27863
rect 21097 27829 21131 27863
rect 21281 27829 21315 27863
rect 21833 27829 21867 27863
rect 8769 27625 8803 27659
rect 10609 27625 10643 27659
rect 14197 27625 14231 27659
rect 15945 27625 15979 27659
rect 16037 27625 16071 27659
rect 19257 27557 19291 27591
rect 13829 27489 13863 27523
rect 14749 27489 14783 27523
rect 20361 27489 20395 27523
rect 21005 27489 21039 27523
rect 21741 27489 21775 27523
rect 7389 27421 7423 27455
rect 9229 27421 9263 27455
rect 12173 27421 12207 27455
rect 12357 27421 12391 27455
rect 12909 27421 12943 27455
rect 13737 27421 13771 27455
rect 13921 27421 13955 27455
rect 15393 27421 15427 27455
rect 15669 27421 15703 27455
rect 15945 27421 15979 27455
rect 17150 27421 17184 27455
rect 17417 27421 17451 27455
rect 17693 27421 17727 27455
rect 17960 27421 17994 27455
rect 19809 27421 19843 27455
rect 21281 27421 21315 27455
rect 21373 27421 21407 27455
rect 21486 27418 21520 27452
rect 21649 27421 21683 27455
rect 22937 27421 22971 27455
rect 23121 27421 23155 27455
rect 23305 27421 23339 27455
rect 25053 27421 25087 27455
rect 34529 27421 34563 27455
rect 7634 27353 7668 27387
rect 9496 27353 9530 27387
rect 12265 27285 12299 27319
rect 13553 27285 13587 27319
rect 15577 27285 15611 27319
rect 15761 27285 15795 27319
rect 19073 27285 19107 27319
rect 20913 27285 20947 27319
rect 22385 27285 22419 27319
rect 22937 27285 22971 27319
rect 23949 27285 23983 27319
rect 24869 27285 24903 27319
rect 9413 27081 9447 27115
rect 12541 27081 12575 27115
rect 19901 27081 19935 27115
rect 21465 27081 21499 27115
rect 22385 27081 22419 27115
rect 23121 27081 23155 27115
rect 13838 27013 13872 27047
rect 16865 27013 16899 27047
rect 21014 27013 21048 27047
rect 23480 27013 23514 27047
rect 9045 26945 9079 26979
rect 9229 26945 9263 26979
rect 11529 26945 11563 26979
rect 11989 26945 12023 26979
rect 12173 26945 12207 26979
rect 12357 26945 12391 26979
rect 14105 26945 14139 26979
rect 14841 26945 14875 26979
rect 15117 26945 15151 26979
rect 15209 26945 15243 26979
rect 15393 26945 15427 26979
rect 15761 26945 15795 26979
rect 16773 26945 16807 26979
rect 17049 26945 17083 26979
rect 18797 26945 18831 26979
rect 19809 26945 19843 26979
rect 21281 26945 21315 26979
rect 21376 26967 21410 27001
rect 21649 26945 21683 26979
rect 22095 26945 22129 26979
rect 22477 26945 22511 26979
rect 22661 26945 22695 26979
rect 22753 26945 22787 26979
rect 22845 26945 22879 26979
rect 15485 26877 15519 26911
rect 16405 26877 16439 26911
rect 17141 26877 17175 26911
rect 18429 26877 18463 26911
rect 19441 26877 19475 26911
rect 22017 26877 22051 26911
rect 23213 26877 23247 26911
rect 11713 26809 11747 26843
rect 17877 26809 17911 26843
rect 11621 26741 11655 26775
rect 11851 26741 11885 26775
rect 12725 26741 12759 26775
rect 14657 26741 14691 26775
rect 14933 26741 14967 26775
rect 15393 26741 15427 26775
rect 15577 26741 15611 26775
rect 15669 26741 15703 26775
rect 15853 26741 15887 26775
rect 17049 26741 17083 26775
rect 17785 26741 17819 26775
rect 19717 26741 19751 26775
rect 21649 26741 21683 26775
rect 24593 26741 24627 26775
rect 12725 26537 12759 26571
rect 13553 26537 13587 26571
rect 17141 26537 17175 26571
rect 20545 26537 20579 26571
rect 22753 26537 22787 26571
rect 23397 26537 23431 26571
rect 14749 26469 14783 26503
rect 19073 26469 19107 26503
rect 19349 26469 19383 26503
rect 11713 26401 11747 26435
rect 12541 26401 12575 26435
rect 13737 26401 13771 26435
rect 16129 26401 16163 26435
rect 17693 26401 17727 26435
rect 20729 26401 20763 26435
rect 21465 26401 21499 26435
rect 22937 26401 22971 26435
rect 23121 26401 23155 26435
rect 9781 26333 9815 26367
rect 11437 26333 11471 26367
rect 11621 26333 11655 26367
rect 11805 26333 11839 26367
rect 11989 26333 12023 26367
rect 12265 26333 12299 26367
rect 12449 26333 12483 26367
rect 13001 26333 13035 26367
rect 13093 26333 13127 26367
rect 13185 26333 13219 26367
rect 13369 26333 13403 26367
rect 13461 26333 13495 26367
rect 14289 26333 14323 26367
rect 15862 26333 15896 26367
rect 16405 26333 16439 26367
rect 17141 26333 17175 26367
rect 17233 26333 17267 26367
rect 17949 26333 17983 26367
rect 19257 26333 19291 26367
rect 19533 26333 19567 26367
rect 19625 26333 19659 26367
rect 19901 26333 19935 26367
rect 19993 26333 20027 26367
rect 20177 26333 20211 26367
rect 20453 26333 20487 26367
rect 21373 26333 21407 26367
rect 22017 26333 22051 26367
rect 22201 26333 22235 26367
rect 22385 26333 22419 26367
rect 22661 26333 22695 26367
rect 23029 26333 23063 26367
rect 23213 26333 23247 26367
rect 23305 26333 23339 26367
rect 23489 26333 23523 26367
rect 10048 26265 10082 26299
rect 12081 26265 12115 26299
rect 13737 26265 13771 26299
rect 17417 26265 17451 26299
rect 20729 26265 20763 26299
rect 20821 26265 20855 26299
rect 21097 26265 21131 26299
rect 22569 26265 22603 26299
rect 11161 26197 11195 26231
rect 11253 26197 11287 26231
rect 14473 26197 14507 26231
rect 17049 26197 17083 26231
rect 19809 26197 19843 26231
rect 20361 26197 20395 26231
rect 21925 26197 21959 26231
rect 22937 26197 22971 26231
rect 8309 25993 8343 26027
rect 23029 25993 23063 26027
rect 10701 25925 10735 25959
rect 12909 25925 12943 25959
rect 15485 25925 15519 25959
rect 15669 25925 15703 25959
rect 19993 25925 20027 25959
rect 23949 25925 23983 25959
rect 9597 25857 9631 25891
rect 11253 25857 11287 25891
rect 11529 25857 11563 25891
rect 12449 25857 12483 25891
rect 12725 25857 12759 25891
rect 13093 25857 13127 25891
rect 13553 25857 13587 25891
rect 14289 25857 14323 25891
rect 14749 25857 14783 25891
rect 14933 25857 14967 25891
rect 15025 25857 15059 25891
rect 15117 25857 15151 25891
rect 15761 25857 15795 25891
rect 16681 25857 16715 25891
rect 16948 25857 16982 25891
rect 18245 25857 18279 25891
rect 20269 25857 20303 25891
rect 20453 25857 20487 25891
rect 20821 25857 20855 25891
rect 21097 25857 21131 25891
rect 21649 25863 21683 25897
rect 22073 25857 22107 25891
rect 22293 25857 22327 25891
rect 22385 25857 22419 25891
rect 22845 25857 22879 25891
rect 23121 25857 23155 25891
rect 24133 25857 24167 25891
rect 24225 25857 24259 25891
rect 12541 25789 12575 25823
rect 13277 25789 13311 25823
rect 14381 25789 14415 25823
rect 15853 25789 15887 25823
rect 20545 25789 20579 25823
rect 20729 25789 20763 25823
rect 21373 25789 21407 25823
rect 23765 25789 23799 25823
rect 23949 25789 23983 25823
rect 12265 25721 12299 25755
rect 12633 25721 12667 25755
rect 15485 25721 15519 25755
rect 18061 25721 18095 25755
rect 21005 25721 21039 25755
rect 21465 25721 21499 25755
rect 22201 25721 22235 25755
rect 11713 25653 11747 25687
rect 13645 25653 13679 25687
rect 14565 25653 14599 25687
rect 15393 25653 15427 25687
rect 16497 25653 16531 25687
rect 20085 25653 20119 25687
rect 21557 25653 21591 25687
rect 22569 25653 22603 25687
rect 22661 25653 22695 25687
rect 23213 25653 23247 25687
rect 11069 25449 11103 25483
rect 12909 25449 12943 25483
rect 13369 25449 13403 25483
rect 13737 25449 13771 25483
rect 14841 25449 14875 25483
rect 15577 25449 15611 25483
rect 18797 25449 18831 25483
rect 20821 25449 20855 25483
rect 22293 25449 22327 25483
rect 10517 25381 10551 25415
rect 12633 25381 12667 25415
rect 17601 25381 17635 25415
rect 20361 25381 20395 25415
rect 10701 25313 10735 25347
rect 11621 25313 11655 25347
rect 12817 25313 12851 25347
rect 13001 25313 13035 25347
rect 13921 25313 13955 25347
rect 16221 25313 16255 25347
rect 17693 25313 17727 25347
rect 21925 25313 21959 25347
rect 22845 25313 22879 25347
rect 10333 25245 10367 25279
rect 10517 25245 10551 25279
rect 10793 25245 10827 25279
rect 11437 25245 11471 25279
rect 11713 25245 11747 25279
rect 12173 25245 12207 25279
rect 12265 25245 12299 25279
rect 12449 25245 12483 25279
rect 12725 25245 12759 25279
rect 13369 25245 13403 25279
rect 13553 25245 13587 25279
rect 13645 25245 13679 25279
rect 14657 25245 14691 25279
rect 14749 25245 14783 25279
rect 14933 25245 14967 25279
rect 15485 25245 15519 25279
rect 15669 25245 15703 25279
rect 16488 25245 16522 25279
rect 17969 25245 18003 25279
rect 19436 25245 19470 25279
rect 19625 25245 19659 25279
rect 19753 25245 19787 25279
rect 19901 25245 19935 25279
rect 20637 25245 20671 25279
rect 20729 25245 20763 25279
rect 20913 25245 20947 25279
rect 22017 25245 22051 25279
rect 23112 25245 23146 25279
rect 25053 25245 25087 25279
rect 11805 25177 11839 25211
rect 11989 25177 12023 25211
rect 14289 25177 14323 25211
rect 14473 25177 14507 25211
rect 18981 25177 19015 25211
rect 19533 25177 19567 25211
rect 20361 25177 20395 25211
rect 11253 25109 11287 25143
rect 13921 25109 13955 25143
rect 18613 25109 18647 25143
rect 18771 25109 18805 25143
rect 19257 25109 19291 25143
rect 20545 25109 20579 25143
rect 24225 25109 24259 25143
rect 24869 25109 24903 25143
rect 12173 24905 12207 24939
rect 13461 24905 13495 24939
rect 14289 24905 14323 24939
rect 17417 24905 17451 24939
rect 19257 24905 19291 24939
rect 21833 24905 21867 24939
rect 15117 24837 15151 24871
rect 19441 24837 19475 24871
rect 9781 24769 9815 24803
rect 9965 24769 9999 24803
rect 10241 24769 10275 24803
rect 10333 24769 10367 24803
rect 10609 24769 10643 24803
rect 10885 24769 10919 24803
rect 10977 24769 11011 24803
rect 11345 24769 11379 24803
rect 11621 24769 11655 24803
rect 12081 24769 12115 24803
rect 12357 24769 12391 24803
rect 13001 24769 13035 24803
rect 13645 24769 13679 24803
rect 13737 24769 13771 24803
rect 13921 24769 13955 24803
rect 14105 24769 14139 24803
rect 14289 24769 14323 24803
rect 14565 24769 14599 24803
rect 14749 24769 14783 24803
rect 14841 24769 14875 24803
rect 15301 24769 15335 24803
rect 15577 24769 15611 24803
rect 16681 24769 16715 24803
rect 17601 24769 17635 24803
rect 17693 24769 17727 24803
rect 17877 24769 17911 24803
rect 17969 24769 18003 24803
rect 18153 24769 18187 24803
rect 19349 24769 19383 24803
rect 19625 24769 19659 24803
rect 19993 24769 20027 24803
rect 20260 24769 20294 24803
rect 22661 24769 22695 24803
rect 22845 24769 22879 24803
rect 22937 24769 22971 24803
rect 23029 24769 23063 24803
rect 10701 24701 10735 24735
rect 12541 24701 12575 24735
rect 13093 24701 13127 24735
rect 15485 24701 15519 24735
rect 15853 24701 15887 24735
rect 17233 24701 17267 24735
rect 22385 24701 22419 24735
rect 23305 24701 23339 24735
rect 9965 24633 9999 24667
rect 13369 24633 13403 24667
rect 13829 24633 13863 24667
rect 14565 24633 14599 24667
rect 17693 24633 17727 24667
rect 21373 24633 21407 24667
rect 10057 24565 10091 24599
rect 10517 24565 10551 24599
rect 11713 24565 11747 24599
rect 11805 24565 11839 24599
rect 11943 24565 11977 24599
rect 15669 24565 15703 24599
rect 15761 24565 15795 24599
rect 18153 24565 18187 24599
rect 19809 24565 19843 24599
rect 13829 24361 13863 24395
rect 18797 24361 18831 24395
rect 20361 24361 20395 24395
rect 21465 24361 21499 24395
rect 10333 24293 10367 24327
rect 10701 24293 10735 24327
rect 13737 24293 13771 24327
rect 18889 24293 18923 24327
rect 22753 24293 22787 24327
rect 11805 24225 11839 24259
rect 13921 24225 13955 24259
rect 14933 24225 14967 24259
rect 15577 24225 15611 24259
rect 18705 24225 18739 24259
rect 19901 24225 19935 24259
rect 21557 24225 21591 24259
rect 22937 24225 22971 24259
rect 8953 24157 8987 24191
rect 10517 24157 10551 24191
rect 12725 24157 12759 24191
rect 13461 24157 13495 24191
rect 13645 24157 13679 24191
rect 14289 24157 14323 24191
rect 14565 24157 14599 24191
rect 15485 24157 15519 24191
rect 17325 24157 17359 24191
rect 17969 24157 18003 24191
rect 18429 24157 18463 24191
rect 18613 24157 18647 24191
rect 18981 24157 19015 24191
rect 21005 24157 21039 24191
rect 21097 24157 21131 24191
rect 21281 24157 21315 24191
rect 22201 24157 22235 24191
rect 22385 24157 22419 24191
rect 22569 24157 22603 24191
rect 22661 24157 22695 24191
rect 23213 24157 23247 24191
rect 25053 24157 25087 24191
rect 9220 24089 9254 24123
rect 14105 24089 14139 24123
rect 14473 24089 14507 24123
rect 17080 24089 17114 24123
rect 17417 24089 17451 24123
rect 11253 24021 11287 24055
rect 12173 24021 12207 24055
rect 12909 24021 12943 24055
rect 15209 24021 15243 24055
rect 15945 24021 15979 24055
rect 18245 24021 18279 24055
rect 19349 24021 19383 24055
rect 22937 24021 22971 24055
rect 23857 24021 23891 24055
rect 24869 24021 24903 24055
rect 9781 23817 9815 23851
rect 10609 23817 10643 23851
rect 12265 23817 12299 23851
rect 12817 23817 12851 23851
rect 14289 23817 14323 23851
rect 15117 23817 15151 23851
rect 15501 23817 15535 23851
rect 15669 23817 15703 23851
rect 16405 23817 16439 23851
rect 19625 23817 19659 23851
rect 22293 23817 22327 23851
rect 23029 23817 23063 23851
rect 15301 23749 15335 23783
rect 18490 23749 18524 23783
rect 20085 23749 20119 23783
rect 23388 23749 23422 23783
rect 9689 23681 9723 23715
rect 9873 23681 9907 23715
rect 10241 23681 10275 23715
rect 11529 23681 11563 23715
rect 11713 23681 11747 23715
rect 11805 23681 11839 23715
rect 12081 23681 12115 23715
rect 13093 23681 13127 23715
rect 13185 23681 13219 23715
rect 13277 23681 13311 23715
rect 13461 23681 13495 23715
rect 14197 23681 14231 23715
rect 14473 23681 14507 23715
rect 14565 23681 14599 23715
rect 14657 23681 14691 23715
rect 14749 23681 14783 23715
rect 14933 23681 14967 23715
rect 15025 23681 15059 23715
rect 15209 23681 15243 23715
rect 15761 23681 15795 23715
rect 15945 23681 15979 23715
rect 16037 23681 16071 23715
rect 16129 23681 16163 23715
rect 17040 23681 17074 23715
rect 19901 23681 19935 23715
rect 19993 23681 20027 23715
rect 20269 23681 20303 23715
rect 22109 23681 22143 23715
rect 22385 23681 22419 23715
rect 22569 23681 22603 23715
rect 22661 23681 22695 23715
rect 22753 23681 22787 23715
rect 10149 23613 10183 23647
rect 11253 23613 11287 23647
rect 11897 23613 11931 23647
rect 14289 23613 14323 23647
rect 16773 23613 16807 23647
rect 18245 23613 18279 23647
rect 21833 23613 21867 23647
rect 23121 23613 23155 23647
rect 10701 23545 10735 23579
rect 13553 23545 13587 23579
rect 21925 23545 21959 23579
rect 14933 23477 14967 23511
rect 15476 23477 15510 23511
rect 18153 23477 18187 23511
rect 19717 23477 19751 23511
rect 24501 23477 24535 23511
rect 10609 23273 10643 23307
rect 11069 23273 11103 23307
rect 13921 23273 13955 23307
rect 14473 23273 14507 23307
rect 17325 23273 17359 23307
rect 19441 23273 19475 23307
rect 19625 23273 19659 23307
rect 22477 23273 22511 23307
rect 22615 23273 22649 23307
rect 17141 23205 17175 23239
rect 21557 23205 21591 23239
rect 14381 23137 14415 23171
rect 15761 23137 15795 23171
rect 16773 23137 16807 23171
rect 17877 23137 17911 23171
rect 18245 23137 18279 23171
rect 21189 23137 21223 23171
rect 21925 23137 21959 23171
rect 10701 23069 10735 23103
rect 12182 23069 12216 23103
rect 12449 23069 12483 23103
rect 12541 23069 12575 23103
rect 14657 23069 14691 23103
rect 14841 23069 14875 23103
rect 14933 23069 14967 23103
rect 16313 23069 16347 23103
rect 16957 23069 16991 23103
rect 17233 23069 17267 23103
rect 18889 23069 18923 23103
rect 19073 23069 19107 23103
rect 20545 23069 20579 23103
rect 21373 23069 21407 23103
rect 21833 23069 21867 23103
rect 22017 23069 22051 23103
rect 22109 23069 22143 23103
rect 22293 23069 22327 23103
rect 22753 23069 22787 23103
rect 22937 23069 22971 23103
rect 25053 23069 25087 23103
rect 12808 23001 12842 23035
rect 18797 23001 18831 23035
rect 19257 23001 19291 23035
rect 19457 23001 19491 23035
rect 23673 23001 23707 23035
rect 23857 23001 23891 23035
rect 15577 22933 15611 22967
rect 18981 22933 19015 22967
rect 20453 22933 20487 22967
rect 21649 22933 21683 22967
rect 22385 22933 22419 22967
rect 23581 22933 23615 22967
rect 24041 22933 24075 22967
rect 24869 22933 24903 22967
rect 16129 22729 16163 22763
rect 17417 22729 17451 22763
rect 21557 22729 21591 22763
rect 22753 22729 22787 22763
rect 24409 22729 24443 22763
rect 15016 22661 15050 22695
rect 16221 22661 16255 22695
rect 23112 22661 23146 22695
rect 9873 22593 9907 22627
rect 10057 22593 10091 22627
rect 10149 22593 10183 22627
rect 11253 22593 11287 22627
rect 12633 22593 12667 22627
rect 13369 22593 13403 22627
rect 13737 22593 13771 22627
rect 14105 22593 14139 22627
rect 14381 22593 14415 22627
rect 14657 22593 14691 22627
rect 16497 22593 16531 22627
rect 16865 22593 16899 22627
rect 17601 22593 17635 22627
rect 19441 22593 19475 22627
rect 19625 22593 19659 22627
rect 19717 22593 19751 22627
rect 19993 22593 20027 22627
rect 20453 22593 20487 22627
rect 20545 22593 20579 22627
rect 20913 22593 20947 22627
rect 21465 22593 21499 22627
rect 21649 22593 21683 22627
rect 22017 22593 22051 22627
rect 22201 22593 22235 22627
rect 22293 22593 22327 22627
rect 22569 22593 22603 22627
rect 24317 22593 24351 22627
rect 24501 22593 24535 22627
rect 10793 22525 10827 22559
rect 13461 22525 13495 22559
rect 14749 22525 14783 22559
rect 16221 22525 16255 22559
rect 17141 22525 17175 22559
rect 17877 22525 17911 22559
rect 18521 22525 18555 22559
rect 19349 22525 19383 22559
rect 19809 22525 19843 22559
rect 20821 22525 20855 22559
rect 22385 22525 22419 22559
rect 22845 22525 22879 22559
rect 21281 22457 21315 22491
rect 9873 22389 9907 22423
rect 10241 22389 10275 22423
rect 11161 22389 11195 22423
rect 12541 22389 12575 22423
rect 13277 22389 13311 22423
rect 13553 22389 13587 22423
rect 13645 22389 13679 22423
rect 14013 22389 14047 22423
rect 14289 22389 14323 22423
rect 14565 22389 14599 22423
rect 16405 22389 16439 22423
rect 17785 22389 17819 22423
rect 17969 22389 18003 22423
rect 18705 22389 18739 22423
rect 20177 22389 20211 22423
rect 24225 22389 24259 22423
rect 19441 22185 19475 22219
rect 20821 22185 20855 22219
rect 23397 22185 23431 22219
rect 23489 22185 23523 22219
rect 10333 22117 10367 22151
rect 13921 22117 13955 22151
rect 15577 22117 15611 22151
rect 19073 22117 19107 22151
rect 8953 22049 8987 22083
rect 10425 22049 10459 22083
rect 12357 22049 12391 22083
rect 14933 22049 14967 22083
rect 16129 22049 16163 22083
rect 16957 22049 16991 22083
rect 23305 22049 23339 22083
rect 2697 21981 2731 22015
rect 10793 21981 10827 22015
rect 10977 21981 11011 22015
rect 11253 21981 11287 22015
rect 11529 21981 11563 22015
rect 11621 21981 11655 22015
rect 12081 21981 12115 22015
rect 12265 21981 12299 22015
rect 12449 21981 12483 22015
rect 12633 21981 12667 22015
rect 13185 21981 13219 22015
rect 13645 21981 13679 22015
rect 13921 21981 13955 22015
rect 14243 21981 14277 22015
rect 14381 21981 14415 22015
rect 14473 21981 14507 22015
rect 14656 21981 14690 22015
rect 14749 21981 14783 22015
rect 14841 21981 14875 22015
rect 15117 21981 15151 22015
rect 15209 21981 15243 22015
rect 15761 21981 15795 22015
rect 15945 21981 15979 22015
rect 16037 21981 16071 22015
rect 17693 21981 17727 22015
rect 17960 21981 17994 22015
rect 19896 21981 19930 22015
rect 20268 21981 20302 22015
rect 20361 21981 20395 22015
rect 20729 21981 20763 22015
rect 21005 21981 21039 22015
rect 21097 21981 21131 22015
rect 23581 21981 23615 22015
rect 1593 21913 1627 21947
rect 9220 21913 9254 21947
rect 10885 21913 10919 21947
rect 13369 21913 13403 21947
rect 19625 21913 19659 21947
rect 19993 21913 20027 21947
rect 20085 21913 20119 21947
rect 11897 21845 11931 21879
rect 13001 21845 13035 21879
rect 13737 21845 13771 21879
rect 14105 21845 14139 21879
rect 15393 21845 15427 21879
rect 16773 21845 16807 21879
rect 17601 21845 17635 21879
rect 19257 21845 19291 21879
rect 19420 21845 19454 21879
rect 19717 21845 19751 21879
rect 21281 21845 21315 21879
rect 9505 21641 9539 21675
rect 10425 21641 10459 21675
rect 11529 21641 11563 21675
rect 12449 21641 12483 21675
rect 15117 21641 15151 21675
rect 16681 21641 16715 21675
rect 18429 21641 18463 21675
rect 22569 21641 22603 21675
rect 12725 21573 12759 21607
rect 12817 21573 12851 21607
rect 17224 21573 17258 21607
rect 8953 21505 8987 21539
rect 9229 21505 9263 21539
rect 10609 21505 10643 21539
rect 10793 21505 10827 21539
rect 10977 21505 11011 21539
rect 11161 21505 11195 21539
rect 11708 21505 11742 21539
rect 11805 21505 11839 21539
rect 11897 21505 11931 21539
rect 12080 21505 12114 21539
rect 12173 21505 12207 21539
rect 12633 21505 12667 21539
rect 13001 21505 13035 21539
rect 13277 21505 13311 21539
rect 13559 21505 13593 21539
rect 13737 21505 13771 21539
rect 14933 21505 14967 21539
rect 15209 21505 15243 21539
rect 15393 21505 15427 21539
rect 16865 21505 16899 21539
rect 19165 21505 19199 21539
rect 19349 21505 19383 21539
rect 19901 21505 19935 21539
rect 20085 21505 20119 21539
rect 20453 21505 20487 21539
rect 21373 21505 21407 21539
rect 21833 21505 21867 21539
rect 22385 21505 22419 21539
rect 22477 21505 22511 21539
rect 22661 21505 22695 21539
rect 9413 21437 9447 21471
rect 10057 21437 10091 21471
rect 10885 21437 10919 21471
rect 13461 21437 13495 21471
rect 13829 21437 13863 21471
rect 14381 21437 14415 21471
rect 15945 21437 15979 21471
rect 16957 21437 16991 21471
rect 19073 21437 19107 21471
rect 19533 21437 19567 21471
rect 20177 21437 20211 21471
rect 20269 21437 20303 21471
rect 22293 21437 22327 21471
rect 23489 21437 23523 21471
rect 18337 21369 18371 21403
rect 9045 21301 9079 21335
rect 13093 21301 13127 21335
rect 13553 21301 13587 21335
rect 14749 21301 14783 21335
rect 15669 21301 15703 21335
rect 16497 21301 16531 21335
rect 20637 21301 20671 21335
rect 20821 21301 20855 21335
rect 22017 21301 22051 21335
rect 22937 21301 22971 21335
rect 8677 21097 8711 21131
rect 12633 21097 12667 21131
rect 13553 21097 13587 21131
rect 13737 21097 13771 21131
rect 14657 21097 14691 21131
rect 15025 21097 15059 21131
rect 15301 21097 15335 21131
rect 15669 21097 15703 21131
rect 23765 21097 23799 21131
rect 14473 21029 14507 21063
rect 18705 21029 18739 21063
rect 19901 21029 19935 21063
rect 8309 20961 8343 20995
rect 8953 20961 8987 20995
rect 10333 20961 10367 20995
rect 12725 20961 12759 20995
rect 13461 20961 13495 20995
rect 14565 20961 14599 20995
rect 21925 20961 21959 20995
rect 8493 20893 8527 20927
rect 8769 20893 8803 20927
rect 10425 20893 10459 20927
rect 12449 20893 12483 20927
rect 12817 20893 12851 20927
rect 14197 20893 14231 20927
rect 14841 20893 14875 20927
rect 16782 20893 16816 20927
rect 17049 20893 17083 20927
rect 17877 20893 17911 20927
rect 18061 20893 18095 20927
rect 18705 20893 18739 20927
rect 18981 20893 19015 20927
rect 20085 20893 20119 20927
rect 20637 20893 20671 20927
rect 20729 20893 20763 20927
rect 21557 20893 21591 20927
rect 21741 20893 21775 20927
rect 21833 20893 21867 20927
rect 22109 20893 22143 20927
rect 22385 20893 22419 20927
rect 13921 20825 13955 20859
rect 14289 20825 14323 20859
rect 14473 20825 14507 20859
rect 15285 20825 15319 20859
rect 15485 20825 15519 20859
rect 22652 20825 22686 20859
rect 9597 20757 9631 20791
rect 9689 20757 9723 20791
rect 11713 20757 11747 20791
rect 12265 20757 12299 20791
rect 13721 20757 13755 20791
rect 15117 20757 15151 20791
rect 17969 20757 18003 20791
rect 18889 20757 18923 20791
rect 22293 20757 22327 20791
rect 9137 20553 9171 20587
rect 10701 20553 10735 20587
rect 14197 20553 14231 20587
rect 15117 20553 15151 20587
rect 21005 20553 21039 20587
rect 9566 20485 9600 20519
rect 11989 20485 12023 20519
rect 16252 20485 16286 20519
rect 16681 20485 16715 20519
rect 19993 20485 20027 20519
rect 23121 20485 23155 20519
rect 23581 20485 23615 20519
rect 11759 20451 11793 20485
rect 9045 20417 9079 20451
rect 9229 20417 9263 20451
rect 10977 20417 11011 20451
rect 11161 20417 11195 20451
rect 12173 20417 12207 20451
rect 12817 20417 12851 20451
rect 13084 20417 13118 20451
rect 20085 20417 20119 20451
rect 20269 20417 20303 20451
rect 20361 20417 20395 20451
rect 20545 20417 20579 20451
rect 20821 20401 20855 20435
rect 22017 20417 22051 20451
rect 22477 20417 22511 20451
rect 23213 20417 23247 20451
rect 23673 20417 23707 20451
rect 9321 20349 9355 20383
rect 11253 20349 11287 20383
rect 14381 20349 14415 20383
rect 16497 20349 16531 20383
rect 17233 20349 17267 20383
rect 21925 20349 21959 20383
rect 22385 20281 22419 20315
rect 23489 20281 23523 20315
rect 10793 20213 10827 20247
rect 11621 20213 11655 20247
rect 11805 20213 11839 20247
rect 12725 20213 12759 20247
rect 15025 20213 15059 20247
rect 18521 20213 18555 20247
rect 20269 20213 20303 20247
rect 20545 20213 20579 20247
rect 23351 20213 23385 20247
rect 9781 20009 9815 20043
rect 13277 20009 13311 20043
rect 15669 20009 15703 20043
rect 16405 20009 16439 20043
rect 19073 20009 19107 20043
rect 20821 20009 20855 20043
rect 20913 20009 20947 20043
rect 21741 20009 21775 20043
rect 22109 20009 22143 20043
rect 22661 20009 22695 20043
rect 11529 19941 11563 19975
rect 15577 19941 15611 19975
rect 10149 19873 10183 19907
rect 13001 19873 13035 19907
rect 14197 19873 14231 19907
rect 16221 19873 16255 19907
rect 9597 19805 9631 19839
rect 9781 19805 9815 19839
rect 12734 19805 12768 19839
rect 13093 19805 13127 19839
rect 13277 19805 13311 19839
rect 14464 19805 14498 19839
rect 16405 19805 16439 19839
rect 16589 19805 16623 19839
rect 17693 19805 17727 19839
rect 19441 19805 19475 19839
rect 21097 19805 21131 19839
rect 21189 19805 21223 19839
rect 21557 19805 21591 19839
rect 21925 19805 21959 19839
rect 22201 19805 22235 19839
rect 22477 19805 22511 19839
rect 33149 19805 33183 19839
rect 10416 19737 10450 19771
rect 17960 19737 17994 19771
rect 19708 19737 19742 19771
rect 22293 19737 22327 19771
rect 34345 19737 34379 19771
rect 11621 19669 11655 19703
rect 10609 19465 10643 19499
rect 12265 19465 12299 19499
rect 14289 19465 14323 19499
rect 18429 19465 18463 19499
rect 18981 19465 19015 19499
rect 21649 19465 21683 19499
rect 11529 19397 11563 19431
rect 14565 19397 14599 19431
rect 12081 19329 12115 19363
rect 12449 19329 12483 19363
rect 12541 19329 12575 19363
rect 14289 19329 14323 19363
rect 15761 19329 15795 19363
rect 18613 19329 18647 19363
rect 18797 19329 18831 19363
rect 18889 19329 18923 19363
rect 19625 19329 19659 19363
rect 20821 19329 20855 19363
rect 21281 19329 21315 19363
rect 21465 19329 21499 19363
rect 11161 19261 11195 19295
rect 14381 19261 14415 19295
rect 15485 19261 15519 19295
rect 20729 19261 20763 19295
rect 1593 14569 1627 14603
rect 1409 14365 1443 14399
rect 34529 13277 34563 13311
rect 34345 13141 34379 13175
rect 1409 7157 1443 7191
rect 34529 5593 34563 5627
rect 20729 2465 20763 2499
rect 13645 2397 13679 2431
rect 20269 2397 20303 2431
rect 1409 2261 1443 2295
rect 6561 2261 6595 2295
rect 27169 2261 27203 2295
rect 34253 2261 34287 2295
<< metal1 >>
rect 1104 39738 34868 39760
rect 1104 39686 5170 39738
rect 5222 39686 5234 39738
rect 5286 39686 5298 39738
rect 5350 39686 5362 39738
rect 5414 39686 5426 39738
rect 5478 39686 13611 39738
rect 13663 39686 13675 39738
rect 13727 39686 13739 39738
rect 13791 39686 13803 39738
rect 13855 39686 13867 39738
rect 13919 39686 22052 39738
rect 22104 39686 22116 39738
rect 22168 39686 22180 39738
rect 22232 39686 22244 39738
rect 22296 39686 22308 39738
rect 22360 39686 30493 39738
rect 30545 39686 30557 39738
rect 30609 39686 30621 39738
rect 30673 39686 30685 39738
rect 30737 39686 30749 39738
rect 30801 39686 34868 39738
rect 1104 39664 34868 39686
rect 17773 39627 17831 39633
rect 17773 39624 17785 39627
rect 16408 39596 17785 39624
rect 16408 39500 16436 39596
rect 17773 39593 17785 39596
rect 17819 39624 17831 39627
rect 18322 39624 18328 39636
rect 17819 39596 18328 39624
rect 17819 39593 17831 39596
rect 17773 39587 17831 39593
rect 18322 39584 18328 39596
rect 18380 39584 18386 39636
rect 22830 39556 22836 39568
rect 21284 39528 22836 39556
rect 14645 39491 14703 39497
rect 14645 39457 14657 39491
rect 14691 39488 14703 39491
rect 14691 39460 15424 39488
rect 14691 39457 14703 39460
rect 14645 39451 14703 39457
rect 1397 39423 1455 39429
rect 1397 39389 1409 39423
rect 1443 39420 1455 39423
rect 1765 39423 1823 39429
rect 1765 39420 1777 39423
rect 1443 39392 1777 39420
rect 1443 39389 1455 39392
rect 1397 39383 1455 39389
rect 1765 39389 1777 39392
rect 1811 39389 1823 39423
rect 1765 39383 1823 39389
rect 2409 39423 2467 39429
rect 2409 39389 2421 39423
rect 2455 39420 2467 39423
rect 2501 39423 2559 39429
rect 2501 39420 2513 39423
rect 2455 39392 2513 39420
rect 2455 39389 2467 39392
rect 2409 39383 2467 39389
rect 2501 39389 2513 39392
rect 2547 39389 2559 39423
rect 2501 39383 2559 39389
rect 3050 39380 3056 39432
rect 3108 39380 3114 39432
rect 8386 39380 8392 39432
rect 8444 39420 8450 39432
rect 8665 39423 8723 39429
rect 8665 39420 8677 39423
rect 8444 39392 8677 39420
rect 8444 39380 8450 39392
rect 8665 39389 8677 39392
rect 8711 39389 8723 39423
rect 8665 39383 8723 39389
rect 14461 39423 14519 39429
rect 14461 39389 14473 39423
rect 14507 39389 14519 39423
rect 14461 39383 14519 39389
rect 14476 39352 14504 39383
rect 14826 39380 14832 39432
rect 14884 39420 14890 39432
rect 15105 39423 15163 39429
rect 15105 39420 15117 39423
rect 14884 39392 15117 39420
rect 14884 39380 14890 39392
rect 15105 39389 15117 39392
rect 15151 39389 15163 39423
rect 15105 39383 15163 39389
rect 15396 39420 15424 39460
rect 16390 39448 16396 39500
rect 16448 39448 16454 39500
rect 17865 39491 17923 39497
rect 17865 39488 17877 39491
rect 16868 39460 17877 39488
rect 16868 39429 16896 39460
rect 17865 39457 17877 39460
rect 17911 39457 17923 39491
rect 17865 39451 17923 39457
rect 15473 39423 15531 39429
rect 15473 39420 15485 39423
rect 15396 39392 15485 39420
rect 14476 39324 14964 39352
rect 1581 39287 1639 39293
rect 1581 39253 1593 39287
rect 1627 39284 1639 39287
rect 4890 39284 4896 39296
rect 1627 39256 4896 39284
rect 1627 39253 1639 39256
rect 1581 39247 1639 39253
rect 4890 39244 4896 39256
rect 4948 39244 4954 39296
rect 8478 39244 8484 39296
rect 8536 39244 8542 39296
rect 13906 39244 13912 39296
rect 13964 39284 13970 39296
rect 14936 39293 14964 39324
rect 15396 39296 15424 39392
rect 15473 39389 15485 39392
rect 15519 39389 15531 39423
rect 15473 39383 15531 39389
rect 15657 39423 15715 39429
rect 15657 39389 15669 39423
rect 15703 39420 15715 39423
rect 15749 39423 15807 39429
rect 15749 39420 15761 39423
rect 15703 39392 15761 39420
rect 15703 39389 15715 39392
rect 15657 39383 15715 39389
rect 15749 39389 15761 39392
rect 15795 39389 15807 39423
rect 15749 39383 15807 39389
rect 16853 39423 16911 39429
rect 16853 39389 16865 39423
rect 16899 39389 16911 39423
rect 16853 39383 16911 39389
rect 17494 39380 17500 39432
rect 17552 39380 17558 39432
rect 17586 39380 17592 39432
rect 17644 39380 17650 39432
rect 18049 39423 18107 39429
rect 18049 39389 18061 39423
rect 18095 39389 18107 39423
rect 18049 39383 18107 39389
rect 16114 39312 16120 39364
rect 16172 39352 16178 39364
rect 17773 39355 17831 39361
rect 17773 39352 17785 39355
rect 16172 39324 17785 39352
rect 16172 39312 16178 39324
rect 17773 39321 17785 39324
rect 17819 39321 17831 39355
rect 18064 39352 18092 39383
rect 18230 39380 18236 39432
rect 18288 39380 18294 39432
rect 21284 39429 21312 39528
rect 22830 39516 22836 39528
rect 22888 39516 22894 39568
rect 21910 39448 21916 39500
rect 21968 39488 21974 39500
rect 22465 39491 22523 39497
rect 22465 39488 22477 39491
rect 21968 39460 22477 39488
rect 21968 39448 21974 39460
rect 22465 39457 22477 39460
rect 22511 39457 22523 39491
rect 22465 39451 22523 39457
rect 34517 39491 34575 39497
rect 34517 39457 34529 39491
rect 34563 39488 34575 39491
rect 35434 39488 35440 39500
rect 34563 39460 35440 39488
rect 34563 39457 34575 39460
rect 34517 39451 34575 39457
rect 35434 39448 35440 39460
rect 35492 39448 35498 39500
rect 20717 39423 20775 39429
rect 20717 39389 20729 39423
rect 20763 39389 20775 39423
rect 20717 39383 20775 39389
rect 21269 39423 21327 39429
rect 21269 39389 21281 39423
rect 21315 39389 21327 39423
rect 21269 39383 21327 39389
rect 22189 39423 22247 39429
rect 22189 39389 22201 39423
rect 22235 39420 22247 39423
rect 23106 39420 23112 39432
rect 22235 39392 23112 39420
rect 22235 39389 22247 39392
rect 22189 39383 22247 39389
rect 19150 39352 19156 39364
rect 18064 39324 19156 39352
rect 17773 39315 17831 39321
rect 19150 39312 19156 39324
rect 19208 39312 19214 39364
rect 20732 39352 20760 39383
rect 23106 39380 23112 39392
rect 23164 39380 23170 39432
rect 22738 39352 22744 39364
rect 20732 39324 22744 39352
rect 22738 39312 22744 39324
rect 22796 39312 22802 39364
rect 14277 39287 14335 39293
rect 14277 39284 14289 39287
rect 13964 39256 14289 39284
rect 13964 39244 13970 39256
rect 14277 39253 14289 39256
rect 14323 39253 14335 39287
rect 14277 39247 14335 39253
rect 14921 39287 14979 39293
rect 14921 39253 14933 39287
rect 14967 39253 14979 39287
rect 14921 39247 14979 39253
rect 15286 39244 15292 39296
rect 15344 39244 15350 39296
rect 15378 39244 15384 39296
rect 15436 39244 15442 39296
rect 17034 39244 17040 39296
rect 17092 39244 17098 39296
rect 17310 39244 17316 39296
rect 17368 39244 17374 39296
rect 20530 39244 20536 39296
rect 20588 39244 20594 39296
rect 21450 39244 21456 39296
rect 21508 39244 21514 39296
rect 1104 39194 35027 39216
rect 1104 39142 9390 39194
rect 9442 39142 9454 39194
rect 9506 39142 9518 39194
rect 9570 39142 9582 39194
rect 9634 39142 9646 39194
rect 9698 39142 17831 39194
rect 17883 39142 17895 39194
rect 17947 39142 17959 39194
rect 18011 39142 18023 39194
rect 18075 39142 18087 39194
rect 18139 39142 26272 39194
rect 26324 39142 26336 39194
rect 26388 39142 26400 39194
rect 26452 39142 26464 39194
rect 26516 39142 26528 39194
rect 26580 39142 34713 39194
rect 34765 39142 34777 39194
rect 34829 39142 34841 39194
rect 34893 39142 34905 39194
rect 34957 39142 34969 39194
rect 35021 39142 35027 39194
rect 1104 39120 35027 39142
rect 2041 39083 2099 39089
rect 2041 39049 2053 39083
rect 2087 39080 2099 39083
rect 3050 39080 3056 39092
rect 2087 39052 3056 39080
rect 2087 39049 2099 39052
rect 2041 39043 2099 39049
rect 3050 39040 3056 39052
rect 3108 39040 3114 39092
rect 13906 39040 13912 39092
rect 13964 39040 13970 39092
rect 14001 39083 14059 39089
rect 14001 39049 14013 39083
rect 14047 39049 14059 39083
rect 14001 39043 14059 39049
rect 15473 39083 15531 39089
rect 15473 39049 15485 39083
rect 15519 39080 15531 39083
rect 16390 39080 16396 39092
rect 15519 39052 16396 39080
rect 15519 39049 15531 39052
rect 15473 39043 15531 39049
rect 1302 38904 1308 38956
rect 1360 38944 1366 38956
rect 1397 38947 1455 38953
rect 1397 38944 1409 38947
rect 1360 38916 1409 38944
rect 1360 38904 1366 38916
rect 1397 38913 1409 38916
rect 1443 38913 1455 38947
rect 1397 38907 1455 38913
rect 13817 38947 13875 38953
rect 13817 38913 13829 38947
rect 13863 38944 13875 38947
rect 13924 38944 13952 39040
rect 14016 39012 14044 39043
rect 16390 39040 16396 39052
rect 16448 39040 16454 39092
rect 17034 39040 17040 39092
rect 17092 39040 17098 39092
rect 20530 39040 20536 39092
rect 20588 39040 20594 39092
rect 21450 39040 21456 39092
rect 21508 39040 21514 39092
rect 21545 39083 21603 39089
rect 21545 39049 21557 39083
rect 21591 39080 21603 39083
rect 21634 39080 21640 39092
rect 21591 39052 21640 39080
rect 21591 39049 21603 39052
rect 21545 39043 21603 39049
rect 21634 39040 21640 39052
rect 21692 39080 21698 39092
rect 21692 39052 23336 39080
rect 21692 39040 21698 39052
rect 14360 39015 14418 39021
rect 14360 39012 14372 39015
rect 14016 38984 14372 39012
rect 14360 38981 14372 38984
rect 14406 38981 14418 39015
rect 17052 39012 17080 39040
rect 17374 39015 17432 39021
rect 17374 39012 17386 39015
rect 14360 38975 14418 38981
rect 15396 38984 16896 39012
rect 17052 38984 17386 39012
rect 15396 38956 15424 38984
rect 13863 38916 13952 38944
rect 13863 38913 13875 38916
rect 13817 38907 13875 38913
rect 15378 38904 15384 38956
rect 15436 38904 15442 38956
rect 16868 38953 16896 38984
rect 17374 38981 17386 38984
rect 17420 38981 17432 39015
rect 17374 38975 17432 38981
rect 20432 39015 20490 39021
rect 20432 38981 20444 39015
rect 20478 39012 20490 39015
rect 20548 39012 20576 39040
rect 20478 38984 20576 39012
rect 21468 39012 21496 39040
rect 22934 39015 22992 39021
rect 22934 39012 22946 39015
rect 21468 38984 22946 39012
rect 20478 38981 20490 38984
rect 20432 38975 20490 38981
rect 22934 38981 22946 38984
rect 22980 38981 22992 39015
rect 22934 38975 22992 38981
rect 23308 38953 23336 39052
rect 15565 38947 15623 38953
rect 15565 38913 15577 38947
rect 15611 38944 15623 38947
rect 16669 38947 16727 38953
rect 16669 38944 16681 38947
rect 15611 38916 16681 38944
rect 15611 38913 15623 38916
rect 15565 38907 15623 38913
rect 16669 38913 16681 38916
rect 16715 38913 16727 38947
rect 16669 38907 16727 38913
rect 16853 38947 16911 38953
rect 16853 38913 16865 38947
rect 16899 38913 16911 38947
rect 16853 38907 16911 38913
rect 23293 38947 23351 38953
rect 23293 38913 23305 38947
rect 23339 38913 23351 38947
rect 23293 38907 23351 38913
rect 14090 38836 14096 38888
rect 14148 38836 14154 38888
rect 15933 38879 15991 38885
rect 15933 38845 15945 38879
rect 15979 38876 15991 38879
rect 16114 38876 16120 38888
rect 15979 38848 16120 38876
rect 15979 38845 15991 38848
rect 15933 38839 15991 38845
rect 16114 38836 16120 38848
rect 16172 38836 16178 38888
rect 16485 38879 16543 38885
rect 16485 38845 16497 38879
rect 16531 38876 16543 38879
rect 17037 38879 17095 38885
rect 17037 38876 17049 38879
rect 16531 38848 17049 38876
rect 16531 38845 16543 38848
rect 16485 38839 16543 38845
rect 17037 38845 17049 38848
rect 17083 38845 17095 38879
rect 17037 38839 17095 38845
rect 17129 38879 17187 38885
rect 17129 38845 17141 38879
rect 17175 38845 17187 38879
rect 17129 38839 17187 38845
rect 17144 38808 17172 38839
rect 19334 38836 19340 38888
rect 19392 38876 19398 38888
rect 20165 38879 20223 38885
rect 20165 38876 20177 38879
rect 19392 38848 20177 38876
rect 19392 38836 19398 38848
rect 20165 38845 20177 38848
rect 20211 38845 20223 38879
rect 20165 38839 20223 38845
rect 23198 38836 23204 38888
rect 23256 38836 23262 38888
rect 17052 38780 17172 38808
rect 17052 38752 17080 38780
rect 15746 38700 15752 38752
rect 15804 38700 15810 38752
rect 17034 38700 17040 38752
rect 17092 38700 17098 38752
rect 18506 38700 18512 38752
rect 18564 38700 18570 38752
rect 21818 38700 21824 38752
rect 21876 38700 21882 38752
rect 23934 38700 23940 38752
rect 23992 38700 23998 38752
rect 1104 38650 34868 38672
rect 1104 38598 5170 38650
rect 5222 38598 5234 38650
rect 5286 38598 5298 38650
rect 5350 38598 5362 38650
rect 5414 38598 5426 38650
rect 5478 38598 13611 38650
rect 13663 38598 13675 38650
rect 13727 38598 13739 38650
rect 13791 38598 13803 38650
rect 13855 38598 13867 38650
rect 13919 38598 22052 38650
rect 22104 38598 22116 38650
rect 22168 38598 22180 38650
rect 22232 38598 22244 38650
rect 22296 38598 22308 38650
rect 22360 38598 30493 38650
rect 30545 38598 30557 38650
rect 30609 38598 30621 38650
rect 30673 38598 30685 38650
rect 30737 38598 30749 38650
rect 30801 38598 34868 38650
rect 1104 38576 34868 38598
rect 15286 38536 15292 38548
rect 13740 38508 15292 38536
rect 4890 38292 4896 38344
rect 4948 38332 4954 38344
rect 7466 38332 7472 38344
rect 4948 38304 7472 38332
rect 4948 38292 4954 38304
rect 7466 38292 7472 38304
rect 7524 38292 7530 38344
rect 8386 38292 8392 38344
rect 8444 38292 8450 38344
rect 8478 38292 8484 38344
rect 8536 38292 8542 38344
rect 13740 38341 13768 38508
rect 15286 38496 15292 38508
rect 15344 38496 15350 38548
rect 18141 38539 18199 38545
rect 18141 38505 18153 38539
rect 18187 38536 18199 38539
rect 18230 38536 18236 38548
rect 18187 38508 18236 38536
rect 18187 38505 18199 38508
rect 18141 38499 18199 38505
rect 18230 38496 18236 38508
rect 18288 38496 18294 38548
rect 22738 38496 22744 38548
rect 22796 38496 22802 38548
rect 22830 38496 22836 38548
rect 22888 38536 22894 38548
rect 23201 38539 23259 38545
rect 23201 38536 23213 38539
rect 22888 38508 23213 38536
rect 22888 38496 22894 38508
rect 23201 38505 23213 38508
rect 23247 38505 23259 38539
rect 23201 38499 23259 38505
rect 20993 38471 21051 38477
rect 20993 38437 21005 38471
rect 21039 38468 21051 38471
rect 21039 38440 21312 38468
rect 21039 38437 21051 38440
rect 20993 38431 21051 38437
rect 21284 38412 21312 38440
rect 15841 38403 15899 38409
rect 15841 38369 15853 38403
rect 15887 38369 15899 38403
rect 15841 38363 15899 38369
rect 13725 38335 13783 38341
rect 13725 38301 13737 38335
rect 13771 38301 13783 38335
rect 13725 38295 13783 38301
rect 14090 38292 14096 38344
rect 14148 38332 14154 38344
rect 14185 38335 14243 38341
rect 14185 38332 14197 38335
rect 14148 38304 14197 38332
rect 14148 38292 14154 38304
rect 14185 38301 14197 38304
rect 14231 38301 14243 38335
rect 14185 38295 14243 38301
rect 15746 38292 15752 38344
rect 15804 38292 15810 38344
rect 15856 38332 15884 38363
rect 18506 38360 18512 38412
rect 18564 38400 18570 38412
rect 18969 38403 19027 38409
rect 18969 38400 18981 38403
rect 18564 38372 18981 38400
rect 18564 38360 18570 38372
rect 18969 38369 18981 38372
rect 19015 38369 19027 38403
rect 18969 38363 19027 38369
rect 21266 38360 21272 38412
rect 21324 38360 21330 38412
rect 21818 38360 21824 38412
rect 21876 38360 21882 38412
rect 21913 38403 21971 38409
rect 21913 38369 21925 38403
rect 21959 38400 21971 38403
rect 23109 38403 23167 38409
rect 23109 38400 23121 38403
rect 21959 38372 23121 38400
rect 21959 38369 21971 38372
rect 21913 38363 21971 38369
rect 23109 38369 23121 38372
rect 23155 38369 23167 38403
rect 23109 38363 23167 38369
rect 23569 38403 23627 38409
rect 23569 38369 23581 38403
rect 23615 38400 23627 38403
rect 23934 38400 23940 38412
rect 23615 38372 23940 38400
rect 23615 38369 23627 38372
rect 23569 38363 23627 38369
rect 23934 38360 23940 38372
rect 23992 38360 23998 38412
rect 17034 38332 17040 38344
rect 15856 38304 17040 38332
rect 17034 38292 17040 38304
rect 17092 38292 17098 38344
rect 17586 38292 17592 38344
rect 17644 38332 17650 38344
rect 18230 38332 18236 38344
rect 17644 38304 18236 38332
rect 17644 38292 17650 38304
rect 18230 38292 18236 38304
rect 18288 38292 18294 38344
rect 19334 38292 19340 38344
rect 19392 38332 19398 38344
rect 19613 38335 19671 38341
rect 19613 38332 19625 38335
rect 19392 38304 19625 38332
rect 19392 38292 19398 38304
rect 19613 38301 19625 38304
rect 19659 38301 19671 38335
rect 21836 38332 21864 38360
rect 22005 38335 22063 38341
rect 22005 38332 22017 38335
rect 21836 38304 22017 38332
rect 19613 38295 19671 38301
rect 22005 38301 22017 38304
rect 22051 38301 22063 38335
rect 22925 38335 22983 38341
rect 22925 38332 22937 38335
rect 22005 38295 22063 38301
rect 22572 38304 22937 38332
rect 14430 38267 14488 38273
rect 14430 38264 14442 38267
rect 13924 38236 14442 38264
rect 5445 38199 5503 38205
rect 5445 38165 5457 38199
rect 5491 38196 5503 38199
rect 6914 38196 6920 38208
rect 5491 38168 6920 38196
rect 5491 38165 5503 38168
rect 5445 38159 5503 38165
rect 6914 38156 6920 38168
rect 6972 38156 6978 38208
rect 8662 38156 8668 38208
rect 8720 38156 8726 38208
rect 13924 38205 13952 38236
rect 14430 38233 14442 38236
rect 14476 38233 14488 38267
rect 15764 38264 15792 38292
rect 16086 38267 16144 38273
rect 16086 38264 16098 38267
rect 15764 38236 16098 38264
rect 14430 38227 14488 38233
rect 16086 38233 16098 38236
rect 16132 38233 16144 38267
rect 16086 38227 16144 38233
rect 13909 38199 13967 38205
rect 13909 38165 13921 38199
rect 13955 38165 13967 38199
rect 13909 38159 13967 38165
rect 15562 38156 15568 38208
rect 15620 38156 15626 38208
rect 17221 38199 17279 38205
rect 17221 38165 17233 38199
rect 17267 38196 17279 38199
rect 17604 38196 17632 38292
rect 19880 38267 19938 38273
rect 19880 38233 19892 38267
rect 19926 38264 19938 38267
rect 20714 38264 20720 38276
rect 19926 38236 20720 38264
rect 19926 38233 19938 38236
rect 19880 38227 19938 38233
rect 20714 38224 20720 38236
rect 20772 38224 20778 38276
rect 22572 38208 22600 38304
rect 22925 38301 22937 38304
rect 22971 38332 22983 38335
rect 23385 38335 23443 38341
rect 23385 38332 23397 38335
rect 22971 38304 23397 38332
rect 22971 38301 22983 38304
rect 22925 38295 22983 38301
rect 23385 38301 23397 38304
rect 23431 38301 23443 38335
rect 23385 38295 23443 38301
rect 17267 38168 17632 38196
rect 17267 38165 17279 38168
rect 17221 38159 17279 38165
rect 18414 38156 18420 38208
rect 18472 38156 18478 38208
rect 22554 38156 22560 38208
rect 22612 38156 22618 38208
rect 22646 38156 22652 38208
rect 22704 38156 22710 38208
rect 1104 38106 35027 38128
rect 1104 38054 9390 38106
rect 9442 38054 9454 38106
rect 9506 38054 9518 38106
rect 9570 38054 9582 38106
rect 9634 38054 9646 38106
rect 9698 38054 17831 38106
rect 17883 38054 17895 38106
rect 17947 38054 17959 38106
rect 18011 38054 18023 38106
rect 18075 38054 18087 38106
rect 18139 38054 26272 38106
rect 26324 38054 26336 38106
rect 26388 38054 26400 38106
rect 26452 38054 26464 38106
rect 26516 38054 26528 38106
rect 26580 38054 34713 38106
rect 34765 38054 34777 38106
rect 34829 38054 34841 38106
rect 34893 38054 34905 38106
rect 34957 38054 34969 38106
rect 35021 38054 35027 38106
rect 1104 38032 35027 38054
rect 8662 37952 8668 38004
rect 8720 37952 8726 38004
rect 14645 37995 14703 38001
rect 14645 37961 14657 37995
rect 14691 37961 14703 37995
rect 14645 37955 14703 37961
rect 8680 37856 8708 37952
rect 14660 37924 14688 37955
rect 17678 37952 17684 38004
rect 17736 37992 17742 38004
rect 17957 37995 18015 38001
rect 17957 37992 17969 37995
rect 17736 37964 17969 37992
rect 17736 37952 17742 37964
rect 17957 37961 17969 37964
rect 18003 37961 18015 37995
rect 17957 37955 18015 37961
rect 20714 37952 20720 38004
rect 20772 37952 20778 38004
rect 21266 37952 21272 38004
rect 21324 37952 21330 38004
rect 21542 37952 21548 38004
rect 21600 37992 21606 38004
rect 21910 37992 21916 38004
rect 21600 37964 21916 37992
rect 21600 37952 21606 37964
rect 21910 37952 21916 37964
rect 21968 37992 21974 38004
rect 22097 37995 22155 38001
rect 22097 37992 22109 37995
rect 21968 37964 22109 37992
rect 21968 37952 21974 37964
rect 22097 37961 22109 37964
rect 22143 37961 22155 37995
rect 22097 37955 22155 37961
rect 14982 37927 15040 37933
rect 14982 37924 14994 37927
rect 9876 37896 14596 37924
rect 14660 37896 14994 37924
rect 8849 37859 8907 37865
rect 8849 37856 8861 37859
rect 8680 37828 8861 37856
rect 8849 37825 8861 37828
rect 8895 37825 8907 37859
rect 8849 37819 8907 37825
rect 5994 37748 6000 37800
rect 6052 37788 6058 37800
rect 8386 37788 8392 37800
rect 6052 37760 8392 37788
rect 6052 37748 6058 37760
rect 8386 37748 8392 37760
rect 8444 37788 8450 37800
rect 9876 37788 9904 37896
rect 10321 37859 10379 37865
rect 10321 37825 10333 37859
rect 10367 37856 10379 37859
rect 10413 37859 10471 37865
rect 10413 37856 10425 37859
rect 10367 37828 10425 37856
rect 10367 37825 10379 37828
rect 10321 37819 10379 37825
rect 10413 37825 10425 37828
rect 10459 37825 10471 37859
rect 10413 37819 10471 37825
rect 10502 37816 10508 37868
rect 10560 37856 10566 37868
rect 10597 37859 10655 37865
rect 10597 37856 10609 37859
rect 10560 37828 10609 37856
rect 10560 37816 10566 37828
rect 10597 37825 10609 37828
rect 10643 37825 10655 37859
rect 10597 37819 10655 37825
rect 10686 37816 10692 37868
rect 10744 37816 10750 37868
rect 10778 37816 10784 37868
rect 10836 37856 10842 37868
rect 10873 37859 10931 37865
rect 10873 37856 10885 37859
rect 10836 37828 10885 37856
rect 10836 37816 10842 37828
rect 10873 37825 10885 37828
rect 10919 37825 10931 37859
rect 10873 37819 10931 37825
rect 11146 37816 11152 37868
rect 11204 37816 11210 37868
rect 11698 37816 11704 37868
rect 11756 37816 11762 37868
rect 13081 37859 13139 37865
rect 13081 37825 13093 37859
rect 13127 37856 13139 37859
rect 13998 37856 14004 37868
rect 13127 37828 14004 37856
rect 13127 37825 13139 37828
rect 13081 37819 13139 37825
rect 13998 37816 14004 37828
rect 14056 37816 14062 37868
rect 14458 37816 14464 37868
rect 14516 37816 14522 37868
rect 14568 37856 14596 37896
rect 14982 37893 14994 37896
rect 15028 37893 15040 37927
rect 15378 37924 15384 37936
rect 14982 37887 15040 37893
rect 15120 37896 15384 37924
rect 15120 37856 15148 37896
rect 15378 37884 15384 37896
rect 15436 37884 15442 37936
rect 17773 37927 17831 37933
rect 17773 37893 17785 37927
rect 17819 37924 17831 37927
rect 18046 37924 18052 37936
rect 17819 37896 18052 37924
rect 17819 37893 17831 37896
rect 17773 37887 17831 37893
rect 18046 37884 18052 37896
rect 18104 37884 18110 37936
rect 19150 37884 19156 37936
rect 19208 37884 19214 37936
rect 19242 37884 19248 37936
rect 19300 37924 19306 37936
rect 21284 37924 21312 37952
rect 21821 37927 21879 37933
rect 21821 37924 21833 37927
rect 19300 37896 19748 37924
rect 19300 37884 19306 37896
rect 14568 37828 15148 37856
rect 17497 37859 17555 37865
rect 17497 37825 17509 37859
rect 17543 37856 17555 37859
rect 17586 37856 17592 37868
rect 17543 37828 17592 37856
rect 17543 37825 17555 37828
rect 17497 37819 17555 37825
rect 17586 37816 17592 37828
rect 17644 37856 17650 37868
rect 18506 37856 18512 37868
rect 17644 37828 18512 37856
rect 17644 37816 17650 37828
rect 18506 37816 18512 37828
rect 18564 37816 18570 37868
rect 18598 37816 18604 37868
rect 18656 37856 18662 37868
rect 19070 37859 19128 37865
rect 19070 37856 19082 37859
rect 18656 37828 19082 37856
rect 18656 37816 18662 37828
rect 19070 37825 19082 37828
rect 19116 37825 19128 37859
rect 19168 37856 19196 37884
rect 19720 37865 19748 37896
rect 21284 37896 21833 37924
rect 19613 37859 19671 37865
rect 19613 37856 19625 37859
rect 19168 37828 19625 37856
rect 19070 37819 19128 37825
rect 19613 37825 19625 37828
rect 19659 37825 19671 37859
rect 19613 37819 19671 37825
rect 19705 37859 19763 37865
rect 19705 37825 19717 37859
rect 19751 37825 19763 37859
rect 20441 37859 20499 37865
rect 20441 37856 20453 37859
rect 19705 37819 19763 37825
rect 19812 37828 20453 37856
rect 8444 37760 9904 37788
rect 8444 37748 8450 37760
rect 11054 37748 11060 37800
rect 11112 37788 11118 37800
rect 11885 37791 11943 37797
rect 11885 37788 11897 37791
rect 11112 37760 11897 37788
rect 11112 37748 11118 37760
rect 11885 37757 11897 37760
rect 11931 37788 11943 37791
rect 11974 37788 11980 37800
rect 11931 37760 11980 37788
rect 11931 37757 11943 37760
rect 11885 37751 11943 37757
rect 11974 37748 11980 37760
rect 12032 37748 12038 37800
rect 14090 37748 14096 37800
rect 14148 37788 14154 37800
rect 14737 37791 14795 37797
rect 14737 37788 14749 37791
rect 14148 37760 14749 37788
rect 14148 37748 14154 37760
rect 14737 37757 14749 37760
rect 14783 37757 14795 37791
rect 14737 37751 14795 37757
rect 17402 37748 17408 37800
rect 17460 37748 17466 37800
rect 17862 37748 17868 37800
rect 17920 37748 17926 37800
rect 19334 37748 19340 37800
rect 19392 37748 19398 37800
rect 19628 37788 19656 37819
rect 19812 37788 19840 37828
rect 20441 37825 20453 37828
rect 20487 37856 20499 37859
rect 20530 37856 20536 37868
rect 20487 37828 20536 37856
rect 20487 37825 20499 37828
rect 20441 37819 20499 37825
rect 20530 37816 20536 37828
rect 20588 37816 20594 37868
rect 20625 37859 20683 37865
rect 20625 37825 20637 37859
rect 20671 37856 20683 37859
rect 20901 37859 20959 37865
rect 20901 37856 20913 37859
rect 20671 37828 20913 37856
rect 20671 37825 20683 37828
rect 20625 37819 20683 37825
rect 20901 37825 20913 37828
rect 20947 37825 20959 37859
rect 21284 37856 21312 37896
rect 21821 37893 21833 37896
rect 21867 37893 21879 37927
rect 21821 37887 21879 37893
rect 22005 37927 22063 37933
rect 22005 37893 22017 37927
rect 22051 37924 22063 37927
rect 22051 37896 22692 37924
rect 22051 37893 22063 37896
rect 22005 37887 22063 37893
rect 21361 37859 21419 37865
rect 21361 37856 21373 37859
rect 21284 37828 21373 37856
rect 20901 37819 20959 37825
rect 21361 37825 21373 37828
rect 21407 37825 21419 37859
rect 21361 37819 21419 37825
rect 21453 37859 21511 37865
rect 21453 37825 21465 37859
rect 21499 37856 21511 37859
rect 21542 37856 21548 37868
rect 21499 37828 21548 37856
rect 21499 37825 21511 37828
rect 21453 37819 21511 37825
rect 21542 37816 21548 37828
rect 21600 37816 21606 37868
rect 21634 37816 21640 37868
rect 21692 37856 21698 37868
rect 22189 37859 22247 37865
rect 22189 37856 22201 37859
rect 21692 37828 22201 37856
rect 21692 37816 21698 37828
rect 22189 37825 22201 37828
rect 22235 37825 22247 37859
rect 22189 37819 22247 37825
rect 19628 37760 19840 37788
rect 20257 37791 20315 37797
rect 20257 37757 20269 37791
rect 20303 37757 20315 37791
rect 22557 37791 22615 37797
rect 22557 37788 22569 37791
rect 20257 37751 20315 37757
rect 21560 37760 22569 37788
rect 11333 37723 11391 37729
rect 11333 37689 11345 37723
rect 11379 37720 11391 37723
rect 12986 37720 12992 37732
rect 11379 37692 12992 37720
rect 11379 37689 11391 37692
rect 11333 37683 11391 37689
rect 12986 37680 12992 37692
rect 13044 37680 13050 37732
rect 16114 37680 16120 37732
rect 16172 37720 16178 37732
rect 16172 37692 17356 37720
rect 16172 37680 16178 37692
rect 7282 37612 7288 37664
rect 7340 37652 7346 37664
rect 7377 37655 7435 37661
rect 7377 37652 7389 37655
rect 7340 37624 7389 37652
rect 7340 37612 7346 37624
rect 7377 37621 7389 37624
rect 7423 37621 7435 37655
rect 7377 37615 7435 37621
rect 9030 37612 9036 37664
rect 9088 37612 9094 37664
rect 10134 37612 10140 37664
rect 10192 37612 10198 37664
rect 10870 37612 10876 37664
rect 10928 37612 10934 37664
rect 11514 37612 11520 37664
rect 11572 37612 11578 37664
rect 12437 37655 12495 37661
rect 12437 37621 12449 37655
rect 12483 37652 12495 37655
rect 12618 37652 12624 37664
rect 12483 37624 12624 37652
rect 12483 37621 12495 37624
rect 12437 37615 12495 37621
rect 12618 37612 12624 37624
rect 12676 37612 12682 37664
rect 12894 37612 12900 37664
rect 12952 37612 12958 37664
rect 17218 37612 17224 37664
rect 17276 37612 17282 37664
rect 17328 37652 17356 37692
rect 17494 37680 17500 37732
rect 17552 37720 17558 37732
rect 17770 37720 17776 37732
rect 17552 37692 17776 37720
rect 17552 37680 17558 37692
rect 17770 37680 17776 37692
rect 17828 37680 17834 37732
rect 20272 37720 20300 37751
rect 21560 37720 21588 37760
rect 22557 37757 22569 37760
rect 22603 37757 22615 37791
rect 22557 37751 22615 37757
rect 22664 37720 22692 37896
rect 23201 37791 23259 37797
rect 23201 37757 23213 37791
rect 23247 37788 23259 37791
rect 23382 37788 23388 37800
rect 23247 37760 23388 37788
rect 23247 37757 23259 37760
rect 23201 37751 23259 37757
rect 23216 37720 23244 37751
rect 23382 37748 23388 37760
rect 23440 37748 23446 37800
rect 20272 37692 21588 37720
rect 22066 37692 23244 37720
rect 18138 37652 18144 37664
rect 17328 37624 18144 37652
rect 18138 37612 18144 37624
rect 18196 37612 18202 37664
rect 19426 37612 19432 37664
rect 19484 37612 19490 37664
rect 21174 37612 21180 37664
rect 21232 37612 21238 37664
rect 21637 37655 21695 37661
rect 21637 37621 21649 37655
rect 21683 37652 21695 37655
rect 22066 37652 22094 37692
rect 21683 37624 22094 37652
rect 21683 37621 21695 37624
rect 21637 37615 21695 37621
rect 22370 37612 22376 37664
rect 22428 37612 22434 37664
rect 1104 37562 34868 37584
rect 1104 37510 5170 37562
rect 5222 37510 5234 37562
rect 5286 37510 5298 37562
rect 5350 37510 5362 37562
rect 5414 37510 5426 37562
rect 5478 37510 13611 37562
rect 13663 37510 13675 37562
rect 13727 37510 13739 37562
rect 13791 37510 13803 37562
rect 13855 37510 13867 37562
rect 13919 37510 22052 37562
rect 22104 37510 22116 37562
rect 22168 37510 22180 37562
rect 22232 37510 22244 37562
rect 22296 37510 22308 37562
rect 22360 37510 30493 37562
rect 30545 37510 30557 37562
rect 30609 37510 30621 37562
rect 30673 37510 30685 37562
rect 30737 37510 30749 37562
rect 30801 37510 34868 37562
rect 1104 37488 34868 37510
rect 10965 37451 11023 37457
rect 10965 37417 10977 37451
rect 11011 37448 11023 37451
rect 11054 37448 11060 37460
rect 11011 37420 11060 37448
rect 11011 37417 11023 37420
rect 10965 37411 11023 37417
rect 11054 37408 11060 37420
rect 11112 37408 11118 37460
rect 13998 37408 14004 37460
rect 14056 37448 14062 37460
rect 14093 37451 14151 37457
rect 14093 37448 14105 37451
rect 14056 37420 14105 37448
rect 14056 37408 14062 37420
rect 14093 37417 14105 37420
rect 14139 37417 14151 37451
rect 14093 37411 14151 37417
rect 14458 37408 14464 37460
rect 14516 37448 14522 37460
rect 15013 37451 15071 37457
rect 15013 37448 15025 37451
rect 14516 37420 15025 37448
rect 14516 37408 14522 37420
rect 15013 37417 15025 37420
rect 15059 37417 15071 37451
rect 15013 37411 15071 37417
rect 17310 37408 17316 37460
rect 17368 37408 17374 37460
rect 17497 37451 17555 37457
rect 17497 37417 17509 37451
rect 17543 37448 17555 37451
rect 17678 37448 17684 37460
rect 17543 37420 17684 37448
rect 17543 37417 17555 37420
rect 17497 37411 17555 37417
rect 17678 37408 17684 37420
rect 17736 37408 17742 37460
rect 17862 37408 17868 37460
rect 17920 37448 17926 37460
rect 18325 37451 18383 37457
rect 18325 37448 18337 37451
rect 17920 37420 18337 37448
rect 17920 37408 17926 37420
rect 18325 37417 18337 37420
rect 18371 37417 18383 37451
rect 18325 37411 18383 37417
rect 19061 37451 19119 37457
rect 19061 37417 19073 37451
rect 19107 37448 19119 37451
rect 19242 37448 19248 37460
rect 19107 37420 19248 37448
rect 19107 37417 19119 37420
rect 19061 37411 19119 37417
rect 19242 37408 19248 37420
rect 19300 37408 19306 37460
rect 21174 37408 21180 37460
rect 21232 37448 21238 37460
rect 22462 37448 22468 37460
rect 21232 37420 22468 37448
rect 21232 37408 21238 37420
rect 22462 37408 22468 37420
rect 22520 37408 22526 37460
rect 22646 37408 22652 37460
rect 22704 37408 22710 37460
rect 15562 37340 15568 37392
rect 15620 37380 15626 37392
rect 17770 37380 17776 37392
rect 15620 37352 17776 37380
rect 15620 37340 15626 37352
rect 7282 37272 7288 37324
rect 7340 37272 7346 37324
rect 16132 37321 16160 37352
rect 17770 37340 17776 37352
rect 17828 37340 17834 37392
rect 16117 37315 16175 37321
rect 16117 37281 16129 37315
rect 16163 37281 16175 37315
rect 16117 37275 16175 37281
rect 17405 37315 17463 37321
rect 17405 37281 17417 37315
rect 17451 37312 17463 37315
rect 18046 37312 18052 37324
rect 17451 37284 18052 37312
rect 17451 37281 17463 37284
rect 17405 37275 17463 37281
rect 18046 37272 18052 37284
rect 18104 37312 18110 37324
rect 22373 37315 22431 37321
rect 18104 37284 18552 37312
rect 18104 37272 18110 37284
rect 6917 37247 6975 37253
rect 6917 37213 6929 37247
rect 6963 37244 6975 37247
rect 8846 37244 8852 37256
rect 6963 37216 7052 37244
rect 6963 37213 6975 37216
rect 6917 37207 6975 37213
rect 7024 37108 7052 37216
rect 8404 37216 8852 37244
rect 8018 37136 8024 37188
rect 8076 37136 8082 37188
rect 8404 37108 8432 37216
rect 8846 37204 8852 37216
rect 8904 37244 8910 37256
rect 9585 37247 9643 37253
rect 9585 37244 9597 37247
rect 8904 37216 9597 37244
rect 8904 37204 8910 37216
rect 9585 37213 9597 37216
rect 9631 37244 9643 37247
rect 11057 37247 11115 37253
rect 11057 37244 11069 37247
rect 9631 37216 11069 37244
rect 9631 37213 9643 37216
rect 9585 37207 9643 37213
rect 11057 37213 11069 37216
rect 11103 37244 11115 37247
rect 12529 37247 12587 37253
rect 12529 37244 12541 37247
rect 11103 37216 12541 37244
rect 11103 37213 11115 37216
rect 11057 37207 11115 37213
rect 12529 37213 12541 37216
rect 12575 37244 12587 37247
rect 14090 37244 14096 37256
rect 12575 37216 14096 37244
rect 12575 37213 12587 37216
rect 12529 37207 12587 37213
rect 14090 37204 14096 37216
rect 14148 37204 14154 37256
rect 14277 37247 14335 37253
rect 14277 37213 14289 37247
rect 14323 37213 14335 37247
rect 14277 37207 14335 37213
rect 9852 37179 9910 37185
rect 9852 37145 9864 37179
rect 9898 37176 9910 37179
rect 10134 37176 10140 37188
rect 9898 37148 10140 37176
rect 9898 37145 9910 37148
rect 9852 37139 9910 37145
rect 10134 37136 10140 37148
rect 10192 37136 10198 37188
rect 11324 37179 11382 37185
rect 11324 37145 11336 37179
rect 11370 37176 11382 37179
rect 11514 37176 11520 37188
rect 11370 37148 11520 37176
rect 11370 37145 11382 37148
rect 11324 37139 11382 37145
rect 11514 37136 11520 37148
rect 11572 37136 11578 37188
rect 12796 37179 12854 37185
rect 12796 37145 12808 37179
rect 12842 37176 12854 37179
rect 12894 37176 12900 37188
rect 12842 37148 12900 37176
rect 12842 37145 12854 37148
rect 12796 37139 12854 37145
rect 12894 37136 12900 37148
rect 12952 37136 12958 37188
rect 13078 37136 13084 37188
rect 13136 37176 13142 37188
rect 14292 37176 14320 37207
rect 14366 37204 14372 37256
rect 14424 37204 14430 37256
rect 15197 37247 15255 37253
rect 15197 37213 15209 37247
rect 15243 37213 15255 37247
rect 15197 37207 15255 37213
rect 15381 37247 15439 37253
rect 15381 37213 15393 37247
rect 15427 37244 15439 37247
rect 15473 37247 15531 37253
rect 15473 37244 15485 37247
rect 15427 37216 15485 37244
rect 15427 37213 15439 37216
rect 15381 37207 15439 37213
rect 15473 37213 15485 37216
rect 15519 37213 15531 37247
rect 15473 37207 15531 37213
rect 16853 37247 16911 37253
rect 16853 37213 16865 37247
rect 16899 37244 16911 37247
rect 17221 37247 17279 37253
rect 17221 37244 17233 37247
rect 16899 37216 17233 37244
rect 16899 37213 16911 37216
rect 16853 37207 16911 37213
rect 17221 37213 17233 37216
rect 17267 37244 17279 37247
rect 17310 37244 17316 37256
rect 17267 37216 17316 37244
rect 17267 37213 17279 37216
rect 17221 37207 17279 37213
rect 13136 37148 14320 37176
rect 15212 37176 15240 37207
rect 17310 37204 17316 37216
rect 17368 37204 17374 37256
rect 17586 37204 17592 37256
rect 17644 37244 17650 37256
rect 17681 37247 17739 37253
rect 17681 37244 17693 37247
rect 17644 37216 17693 37244
rect 17644 37204 17650 37216
rect 17681 37213 17693 37216
rect 17727 37213 17739 37247
rect 17681 37207 17739 37213
rect 18138 37204 18144 37256
rect 18196 37204 18202 37256
rect 18524 37253 18552 37284
rect 22373 37281 22385 37315
rect 22419 37312 22431 37315
rect 22664 37312 22692 37408
rect 22419 37284 22692 37312
rect 22419 37281 22431 37284
rect 22373 37275 22431 37281
rect 18509 37247 18567 37253
rect 18509 37213 18521 37247
rect 18555 37244 18567 37247
rect 18555 37216 18644 37244
rect 18555 37213 18567 37216
rect 18509 37207 18567 37213
rect 18049 37179 18107 37185
rect 15212 37148 15424 37176
rect 13136 37136 13142 37148
rect 15396 37120 15424 37148
rect 18049 37145 18061 37179
rect 18095 37176 18107 37179
rect 18230 37176 18236 37188
rect 18095 37148 18236 37176
rect 18095 37145 18107 37148
rect 18049 37139 18107 37145
rect 18230 37136 18236 37148
rect 18288 37136 18294 37188
rect 7024 37080 8432 37108
rect 8711 37111 8769 37117
rect 8711 37077 8723 37111
rect 8757 37108 8769 37111
rect 9122 37108 9128 37120
rect 8757 37080 9128 37108
rect 8757 37077 8769 37080
rect 8711 37071 8769 37077
rect 9122 37068 9128 37080
rect 9180 37068 9186 37120
rect 12434 37068 12440 37120
rect 12492 37068 12498 37120
rect 13262 37068 13268 37120
rect 13320 37108 13326 37120
rect 13909 37111 13967 37117
rect 13909 37108 13921 37111
rect 13320 37080 13921 37108
rect 13320 37068 13326 37080
rect 13909 37077 13921 37080
rect 13955 37077 13967 37111
rect 13909 37071 13967 37077
rect 15378 37068 15384 37120
rect 15436 37068 15442 37120
rect 16209 37111 16267 37117
rect 16209 37077 16221 37111
rect 16255 37108 16267 37111
rect 16298 37108 16304 37120
rect 16255 37080 16304 37108
rect 16255 37077 16267 37080
rect 16209 37071 16267 37077
rect 16298 37068 16304 37080
rect 16356 37068 16362 37120
rect 16942 37068 16948 37120
rect 17000 37068 17006 37120
rect 17034 37068 17040 37120
rect 17092 37108 17098 37120
rect 17678 37108 17684 37120
rect 17092 37080 17684 37108
rect 17092 37068 17098 37080
rect 17678 37068 17684 37080
rect 17736 37068 17742 37120
rect 17957 37111 18015 37117
rect 17957 37077 17969 37111
rect 18003 37108 18015 37111
rect 18322 37108 18328 37120
rect 18003 37080 18328 37108
rect 18003 37077 18015 37080
rect 17957 37071 18015 37077
rect 18322 37068 18328 37080
rect 18380 37068 18386 37120
rect 18616 37108 18644 37216
rect 19334 37204 19340 37256
rect 19392 37244 19398 37256
rect 20622 37244 20628 37256
rect 19392 37216 20628 37244
rect 19392 37204 19398 37216
rect 20622 37204 20628 37216
rect 20680 37204 20686 37256
rect 20714 37204 20720 37256
rect 20772 37204 20778 37256
rect 20901 37247 20959 37253
rect 20901 37213 20913 37247
rect 20947 37213 20959 37247
rect 20901 37207 20959 37213
rect 19058 37136 19064 37188
rect 19116 37176 19122 37188
rect 20358 37179 20416 37185
rect 20358 37176 20370 37179
rect 19116 37148 20370 37176
rect 19116 37136 19122 37148
rect 20358 37145 20370 37148
rect 20404 37145 20416 37179
rect 20358 37139 20416 37145
rect 20530 37136 20536 37188
rect 20588 37176 20594 37188
rect 20916 37176 20944 37207
rect 21910 37204 21916 37256
rect 21968 37244 21974 37256
rect 22189 37247 22247 37253
rect 22189 37244 22201 37247
rect 21968 37216 22201 37244
rect 21968 37204 21974 37216
rect 22189 37213 22201 37216
rect 22235 37213 22247 37247
rect 22189 37207 22247 37213
rect 22554 37204 22560 37256
rect 22612 37204 22618 37256
rect 22741 37247 22799 37253
rect 22741 37213 22753 37247
rect 22787 37244 22799 37247
rect 22833 37247 22891 37253
rect 22833 37244 22845 37247
rect 22787 37216 22845 37244
rect 22787 37213 22799 37216
rect 22741 37207 22799 37213
rect 22833 37213 22845 37216
rect 22879 37213 22891 37247
rect 22833 37207 22891 37213
rect 22572 37176 22600 37204
rect 20588 37148 22600 37176
rect 20588 37136 20594 37148
rect 19245 37111 19303 37117
rect 19245 37108 19257 37111
rect 18616 37080 19257 37108
rect 19245 37077 19257 37080
rect 19291 37077 19303 37111
rect 19245 37071 19303 37077
rect 21082 37068 21088 37120
rect 21140 37068 21146 37120
rect 21634 37068 21640 37120
rect 21692 37068 21698 37120
rect 23014 37068 23020 37120
rect 23072 37068 23078 37120
rect 1104 37018 35027 37040
rect 1104 36966 9390 37018
rect 9442 36966 9454 37018
rect 9506 36966 9518 37018
rect 9570 36966 9582 37018
rect 9634 36966 9646 37018
rect 9698 36966 17831 37018
rect 17883 36966 17895 37018
rect 17947 36966 17959 37018
rect 18011 36966 18023 37018
rect 18075 36966 18087 37018
rect 18139 36966 26272 37018
rect 26324 36966 26336 37018
rect 26388 36966 26400 37018
rect 26452 36966 26464 37018
rect 26516 36966 26528 37018
rect 26580 36966 34713 37018
rect 34765 36966 34777 37018
rect 34829 36966 34841 37018
rect 34893 36966 34905 37018
rect 34957 36966 34969 37018
rect 35021 36966 35027 37018
rect 1104 36944 35027 36966
rect 8018 36864 8024 36916
rect 8076 36864 8082 36916
rect 12434 36864 12440 36916
rect 12492 36864 12498 36916
rect 12805 36907 12863 36913
rect 12805 36873 12817 36907
rect 12851 36904 12863 36907
rect 13262 36904 13268 36916
rect 12851 36876 13268 36904
rect 12851 36873 12863 36876
rect 12805 36867 12863 36873
rect 13262 36864 13268 36876
rect 13320 36864 13326 36916
rect 13909 36907 13967 36913
rect 13909 36873 13921 36907
rect 13955 36904 13967 36907
rect 14366 36904 14372 36916
rect 13955 36876 14372 36904
rect 13955 36873 13967 36876
rect 13909 36867 13967 36873
rect 14366 36864 14372 36876
rect 14424 36864 14430 36916
rect 15749 36907 15807 36913
rect 15749 36873 15761 36907
rect 15795 36904 15807 36907
rect 15795 36876 17264 36904
rect 15795 36873 15807 36876
rect 15749 36867 15807 36873
rect 9030 36845 9036 36848
rect 9024 36836 9036 36845
rect 8991 36808 9036 36836
rect 9024 36799 9036 36808
rect 9030 36796 9036 36799
rect 9088 36796 9094 36848
rect 7466 36728 7472 36780
rect 7524 36728 7530 36780
rect 8757 36771 8815 36777
rect 8757 36737 8769 36771
rect 8803 36768 8815 36771
rect 8846 36768 8852 36780
rect 8803 36740 8852 36768
rect 8803 36737 8815 36740
rect 8757 36731 8815 36737
rect 8846 36728 8852 36740
rect 8904 36728 8910 36780
rect 10042 36728 10048 36780
rect 10100 36768 10106 36780
rect 12452 36777 12480 36864
rect 17034 36836 17040 36848
rect 16684 36808 17040 36836
rect 10413 36771 10471 36777
rect 10413 36768 10425 36771
rect 10100 36740 10425 36768
rect 10100 36728 10106 36740
rect 10413 36737 10425 36740
rect 10459 36737 10471 36771
rect 10413 36731 10471 36737
rect 12437 36771 12495 36777
rect 12437 36737 12449 36771
rect 12483 36768 12495 36771
rect 12894 36768 12900 36780
rect 12483 36740 12900 36768
rect 12483 36737 12495 36740
rect 12437 36731 12495 36737
rect 12894 36728 12900 36740
rect 12952 36728 12958 36780
rect 16684 36777 16712 36808
rect 17034 36796 17040 36808
rect 17092 36796 17098 36848
rect 17236 36836 17264 36876
rect 17310 36864 17316 36916
rect 17368 36904 17374 36916
rect 18049 36907 18107 36913
rect 18049 36904 18061 36907
rect 17368 36876 18061 36904
rect 17368 36864 17374 36876
rect 18049 36873 18061 36876
rect 18095 36873 18107 36907
rect 18049 36867 18107 36873
rect 20530 36864 20536 36916
rect 20588 36864 20594 36916
rect 21634 36864 21640 36916
rect 21692 36864 21698 36916
rect 21910 36864 21916 36916
rect 21968 36864 21974 36916
rect 23382 36864 23388 36916
rect 23440 36864 23446 36916
rect 17236 36808 17448 36836
rect 12989 36771 13047 36777
rect 12989 36737 13001 36771
rect 13035 36768 13047 36771
rect 15565 36771 15623 36777
rect 13035 36740 13400 36768
rect 13035 36737 13047 36740
rect 12989 36731 13047 36737
rect 8570 36660 8576 36712
rect 8628 36660 8634 36712
rect 10594 36660 10600 36712
rect 10652 36660 10658 36712
rect 10781 36703 10839 36709
rect 10781 36669 10793 36703
rect 10827 36700 10839 36703
rect 10870 36700 10876 36712
rect 10827 36672 10876 36700
rect 10827 36669 10839 36672
rect 10781 36663 10839 36669
rect 10137 36635 10195 36641
rect 10137 36601 10149 36635
rect 10183 36632 10195 36635
rect 10796 36632 10824 36663
rect 10870 36660 10876 36672
rect 10928 36660 10934 36712
rect 12526 36660 12532 36712
rect 12584 36660 12590 36712
rect 12621 36703 12679 36709
rect 12621 36669 12633 36703
rect 12667 36700 12679 36703
rect 12710 36700 12716 36712
rect 12667 36672 12716 36700
rect 12667 36669 12679 36672
rect 12621 36663 12679 36669
rect 12710 36660 12716 36672
rect 12768 36660 12774 36712
rect 13265 36703 13323 36709
rect 13265 36669 13277 36703
rect 13311 36669 13323 36703
rect 13265 36663 13323 36669
rect 10183 36604 10824 36632
rect 12728 36632 12756 36660
rect 13280 36632 13308 36663
rect 12728 36604 13308 36632
rect 10183 36601 10195 36604
rect 10137 36595 10195 36601
rect 13372 36576 13400 36740
rect 15565 36737 15577 36771
rect 15611 36768 15623 36771
rect 16669 36771 16727 36777
rect 15611 36740 16436 36768
rect 15611 36737 15623 36740
rect 15565 36731 15623 36737
rect 13446 36660 13452 36712
rect 13504 36700 13510 36712
rect 14001 36703 14059 36709
rect 14001 36700 14013 36703
rect 13504 36672 14013 36700
rect 13504 36660 13510 36672
rect 14001 36669 14013 36672
rect 14047 36669 14059 36703
rect 14001 36663 14059 36669
rect 15930 36660 15936 36712
rect 15988 36660 15994 36712
rect 7650 36524 7656 36576
rect 7708 36524 7714 36576
rect 10226 36524 10232 36576
rect 10284 36524 10290 36576
rect 11238 36524 11244 36576
rect 11296 36564 11302 36576
rect 11333 36567 11391 36573
rect 11333 36564 11345 36567
rect 11296 36536 11345 36564
rect 11296 36524 11302 36536
rect 11333 36533 11345 36536
rect 11379 36533 11391 36567
rect 11333 36527 11391 36533
rect 11793 36567 11851 36573
rect 11793 36533 11805 36567
rect 11839 36564 11851 36567
rect 12434 36564 12440 36576
rect 11839 36536 12440 36564
rect 11839 36533 11851 36536
rect 11793 36527 11851 36533
rect 12434 36524 12440 36536
rect 12492 36524 12498 36576
rect 13170 36524 13176 36576
rect 13228 36524 13234 36576
rect 13354 36524 13360 36576
rect 13412 36524 13418 36576
rect 14642 36524 14648 36576
rect 14700 36524 14706 36576
rect 16408 36564 16436 36740
rect 16669 36737 16681 36771
rect 16715 36737 16727 36771
rect 16925 36771 16983 36777
rect 16925 36768 16937 36771
rect 16669 36731 16727 36737
rect 16776 36740 16937 36768
rect 16485 36703 16543 36709
rect 16485 36669 16497 36703
rect 16531 36700 16543 36703
rect 16776 36700 16804 36740
rect 16925 36737 16937 36740
rect 16971 36737 16983 36771
rect 17420 36768 17448 36808
rect 17678 36796 17684 36848
rect 17736 36836 17742 36848
rect 18233 36839 18291 36845
rect 18233 36836 18245 36839
rect 17736 36808 18245 36836
rect 17736 36796 17742 36808
rect 18233 36805 18245 36808
rect 18279 36836 18291 36839
rect 19334 36836 19340 36848
rect 18279 36808 19340 36836
rect 18279 36805 18291 36808
rect 18233 36799 18291 36805
rect 19334 36796 19340 36808
rect 19392 36796 19398 36848
rect 20548 36836 20576 36864
rect 20548 36808 21404 36836
rect 18598 36768 18604 36780
rect 17420 36740 18604 36768
rect 16925 36731 16983 36737
rect 18598 36728 18604 36740
rect 18656 36728 18662 36780
rect 19978 36728 19984 36780
rect 20036 36728 20042 36780
rect 21376 36777 21404 36808
rect 20257 36771 20315 36777
rect 20257 36737 20269 36771
rect 20303 36768 20315 36771
rect 21177 36771 21235 36777
rect 21177 36768 21189 36771
rect 20303 36740 21189 36768
rect 20303 36737 20315 36740
rect 20257 36731 20315 36737
rect 21177 36737 21189 36740
rect 21223 36737 21235 36771
rect 21177 36731 21235 36737
rect 21361 36771 21419 36777
rect 21361 36737 21373 36771
rect 21407 36737 21419 36771
rect 21361 36731 21419 36737
rect 21545 36771 21603 36777
rect 21545 36737 21557 36771
rect 21591 36768 21603 36771
rect 21652 36768 21680 36864
rect 23014 36796 23020 36848
rect 23072 36845 23078 36848
rect 23072 36799 23084 36845
rect 23308 36808 24808 36836
rect 23072 36796 23078 36799
rect 21591 36740 21680 36768
rect 21591 36737 21603 36740
rect 21545 36731 21603 36737
rect 23198 36728 23204 36780
rect 23256 36768 23262 36780
rect 23308 36777 23336 36808
rect 23293 36771 23351 36777
rect 23293 36768 23305 36771
rect 23256 36740 23305 36768
rect 23256 36728 23262 36740
rect 23293 36737 23305 36740
rect 23339 36737 23351 36771
rect 23293 36731 23351 36737
rect 24486 36728 24492 36780
rect 24544 36777 24550 36780
rect 24780 36777 24808 36808
rect 24544 36731 24556 36777
rect 24765 36771 24823 36777
rect 24765 36737 24777 36771
rect 24811 36737 24823 36771
rect 24765 36731 24823 36737
rect 24544 36728 24550 36731
rect 16531 36672 16804 36700
rect 16531 36669 16543 36672
rect 16485 36663 16543 36669
rect 19426 36660 19432 36712
rect 19484 36660 19490 36712
rect 20530 36660 20536 36712
rect 20588 36660 20594 36712
rect 19444 36564 19472 36660
rect 16408 36536 19472 36564
rect 20070 36524 20076 36576
rect 20128 36524 20134 36576
rect 20714 36524 20720 36576
rect 20772 36564 20778 36576
rect 21085 36567 21143 36573
rect 21085 36564 21097 36567
rect 20772 36536 21097 36564
rect 20772 36524 20778 36536
rect 21085 36533 21097 36536
rect 21131 36533 21143 36567
rect 21085 36527 21143 36533
rect 1104 36474 34868 36496
rect 1104 36422 5170 36474
rect 5222 36422 5234 36474
rect 5286 36422 5298 36474
rect 5350 36422 5362 36474
rect 5414 36422 5426 36474
rect 5478 36422 13611 36474
rect 13663 36422 13675 36474
rect 13727 36422 13739 36474
rect 13791 36422 13803 36474
rect 13855 36422 13867 36474
rect 13919 36422 22052 36474
rect 22104 36422 22116 36474
rect 22168 36422 22180 36474
rect 22232 36422 22244 36474
rect 22296 36422 22308 36474
rect 22360 36422 30493 36474
rect 30545 36422 30557 36474
rect 30609 36422 30621 36474
rect 30673 36422 30685 36474
rect 30737 36422 30749 36474
rect 30801 36422 34868 36474
rect 1104 36400 34868 36422
rect 7929 36363 7987 36369
rect 7929 36329 7941 36363
rect 7975 36360 7987 36363
rect 8570 36360 8576 36372
rect 7975 36332 8576 36360
rect 7975 36329 7987 36332
rect 7929 36323 7987 36329
rect 8570 36320 8576 36332
rect 8628 36320 8634 36372
rect 9122 36320 9128 36372
rect 9180 36320 9186 36372
rect 10226 36320 10232 36372
rect 10284 36320 10290 36372
rect 10594 36320 10600 36372
rect 10652 36360 10658 36372
rect 10965 36363 11023 36369
rect 10965 36360 10977 36363
rect 10652 36332 10977 36360
rect 10652 36320 10658 36332
rect 10965 36329 10977 36332
rect 11011 36329 11023 36363
rect 10965 36323 11023 36329
rect 11698 36320 11704 36372
rect 11756 36320 11762 36372
rect 12253 36363 12311 36369
rect 12253 36329 12265 36363
rect 12299 36360 12311 36363
rect 12526 36360 12532 36372
rect 12299 36332 12532 36360
rect 12299 36329 12311 36332
rect 12253 36323 12311 36329
rect 12526 36320 12532 36332
rect 12584 36320 12590 36372
rect 12894 36320 12900 36372
rect 12952 36320 12958 36372
rect 12986 36320 12992 36372
rect 13044 36320 13050 36372
rect 13081 36363 13139 36369
rect 13081 36329 13093 36363
rect 13127 36360 13139 36363
rect 13262 36360 13268 36372
rect 13127 36332 13268 36360
rect 13127 36329 13139 36332
rect 13081 36323 13139 36329
rect 13262 36320 13268 36332
rect 13320 36320 13326 36372
rect 13354 36320 13360 36372
rect 13412 36360 13418 36372
rect 13412 36332 15516 36360
rect 13412 36320 13418 36332
rect 9140 36233 9168 36320
rect 9125 36227 9183 36233
rect 9125 36193 9137 36227
rect 9171 36193 9183 36227
rect 9125 36187 9183 36193
rect 934 36116 940 36168
rect 992 36156 998 36168
rect 1397 36159 1455 36165
rect 1397 36156 1409 36159
rect 992 36128 1409 36156
rect 992 36116 998 36128
rect 1397 36125 1409 36128
rect 1443 36125 1455 36159
rect 1397 36119 1455 36125
rect 6914 36116 6920 36168
rect 6972 36156 6978 36168
rect 7837 36159 7895 36165
rect 7837 36156 7849 36159
rect 6972 36128 7849 36156
rect 6972 36116 6978 36128
rect 7837 36125 7849 36128
rect 7883 36125 7895 36159
rect 7837 36119 7895 36125
rect 10137 36159 10195 36165
rect 10137 36125 10149 36159
rect 10183 36156 10195 36159
rect 10244 36156 10272 36320
rect 11716 36292 11744 36320
rect 12345 36295 12403 36301
rect 12345 36292 12357 36295
rect 11716 36264 12357 36292
rect 12345 36261 12357 36264
rect 12391 36261 12403 36295
rect 12345 36255 12403 36261
rect 10778 36184 10784 36236
rect 10836 36184 10842 36236
rect 11146 36184 11152 36236
rect 11204 36224 11210 36236
rect 11517 36227 11575 36233
rect 11517 36224 11529 36227
rect 11204 36196 11529 36224
rect 11204 36184 11210 36196
rect 11517 36193 11529 36196
rect 11563 36224 11575 36227
rect 11701 36227 11759 36233
rect 11701 36224 11713 36227
rect 11563 36196 11713 36224
rect 11563 36193 11575 36196
rect 11517 36187 11575 36193
rect 11701 36193 11713 36196
rect 11747 36193 11759 36227
rect 11701 36187 11759 36193
rect 12618 36184 12624 36236
rect 12676 36224 12682 36236
rect 12713 36227 12771 36233
rect 12713 36224 12725 36227
rect 12676 36196 12725 36224
rect 12676 36184 12682 36196
rect 12713 36193 12725 36196
rect 12759 36193 12771 36227
rect 12713 36187 12771 36193
rect 10183 36128 10272 36156
rect 10183 36125 10195 36128
rect 10137 36119 10195 36125
rect 10229 36091 10287 36097
rect 10229 36057 10241 36091
rect 10275 36088 10287 36091
rect 10686 36088 10692 36100
rect 10275 36060 10692 36088
rect 10275 36057 10287 36060
rect 10229 36051 10287 36057
rect 10686 36048 10692 36060
rect 10744 36048 10750 36100
rect 10796 36088 10824 36184
rect 10870 36116 10876 36168
rect 10928 36156 10934 36168
rect 11885 36159 11943 36165
rect 11885 36156 11897 36159
rect 10928 36128 11897 36156
rect 10928 36116 10934 36128
rect 11885 36125 11897 36128
rect 11931 36125 11943 36159
rect 11885 36119 11943 36125
rect 11974 36116 11980 36168
rect 12032 36116 12038 36168
rect 12912 36165 12940 36320
rect 13004 36224 13032 36320
rect 13265 36227 13323 36233
rect 13265 36224 13277 36227
rect 13004 36196 13277 36224
rect 13265 36193 13277 36196
rect 13311 36193 13323 36227
rect 13265 36187 13323 36193
rect 13372 36165 13400 36320
rect 15488 36304 15516 36332
rect 15930 36320 15936 36372
rect 15988 36360 15994 36372
rect 16761 36363 16819 36369
rect 16761 36360 16773 36363
rect 15988 36332 16773 36360
rect 15988 36320 15994 36332
rect 16761 36329 16773 36332
rect 16807 36329 16819 36363
rect 16761 36323 16819 36329
rect 16868 36332 17264 36360
rect 15470 36252 15476 36304
rect 15528 36252 15534 36304
rect 15841 36227 15899 36233
rect 15841 36193 15853 36227
rect 15887 36224 15899 36227
rect 16758 36224 16764 36236
rect 15887 36196 16764 36224
rect 15887 36193 15899 36196
rect 15841 36187 15899 36193
rect 16758 36184 16764 36196
rect 16816 36184 16822 36236
rect 12529 36159 12587 36165
rect 12529 36125 12541 36159
rect 12575 36125 12587 36159
rect 12529 36119 12587 36125
rect 12897 36159 12955 36165
rect 12897 36125 12909 36159
rect 12943 36125 12955 36159
rect 12897 36119 12955 36125
rect 13173 36159 13231 36165
rect 13173 36125 13185 36159
rect 13219 36125 13231 36159
rect 13173 36119 13231 36125
rect 13357 36159 13415 36165
rect 13357 36125 13369 36159
rect 13403 36125 13415 36159
rect 13357 36119 13415 36125
rect 12069 36091 12127 36097
rect 12069 36088 12081 36091
rect 10796 36060 12081 36088
rect 12069 36057 12081 36060
rect 12115 36057 12127 36091
rect 12069 36051 12127 36057
rect 12544 36032 12572 36119
rect 12710 36048 12716 36100
rect 12768 36088 12774 36100
rect 13188 36088 13216 36119
rect 14090 36116 14096 36168
rect 14148 36116 14154 36168
rect 14360 36159 14418 36165
rect 14360 36125 14372 36159
rect 14406 36156 14418 36159
rect 14642 36156 14648 36168
rect 14406 36128 14648 36156
rect 14406 36125 14418 36128
rect 14360 36119 14418 36125
rect 14642 36116 14648 36128
rect 14700 36116 14706 36168
rect 16025 36159 16083 36165
rect 16025 36125 16037 36159
rect 16071 36156 16083 36159
rect 16393 36159 16451 36165
rect 16071 36128 16344 36156
rect 16071 36125 16083 36128
rect 16025 36119 16083 36125
rect 12768 36060 13216 36088
rect 14108 36088 14136 36116
rect 14108 36060 14596 36088
rect 12768 36048 12774 36060
rect 14568 36032 14596 36060
rect 9766 35980 9772 36032
rect 9824 35980 9830 36032
rect 9950 35980 9956 36032
rect 10008 35980 10014 36032
rect 12526 35980 12532 36032
rect 12584 36020 12590 36032
rect 13078 36020 13084 36032
rect 12584 35992 13084 36020
rect 12584 35980 12590 35992
rect 13078 35980 13084 35992
rect 13136 35980 13142 36032
rect 13630 35980 13636 36032
rect 13688 35980 13694 36032
rect 14550 35980 14556 36032
rect 14608 35980 14614 36032
rect 16206 35980 16212 36032
rect 16264 35980 16270 36032
rect 16316 36020 16344 36128
rect 16393 36125 16405 36159
rect 16439 36125 16451 36159
rect 16393 36119 16451 36125
rect 16485 36159 16543 36165
rect 16485 36125 16497 36159
rect 16531 36156 16543 36159
rect 16868 36156 16896 36332
rect 16942 36184 16948 36236
rect 17000 36224 17006 36236
rect 17236 36224 17264 36332
rect 19058 36320 19064 36372
rect 19116 36320 19122 36372
rect 20824 36332 22094 36360
rect 17310 36252 17316 36304
rect 17368 36292 17374 36304
rect 19245 36295 19303 36301
rect 19245 36292 19257 36295
rect 17368 36264 19257 36292
rect 17368 36252 17374 36264
rect 19245 36261 19257 36264
rect 19291 36261 19303 36295
rect 19245 36255 19303 36261
rect 20438 36252 20444 36304
rect 20496 36292 20502 36304
rect 20717 36295 20775 36301
rect 20717 36292 20729 36295
rect 20496 36264 20729 36292
rect 20496 36252 20502 36264
rect 20717 36261 20729 36264
rect 20763 36261 20775 36295
rect 20717 36255 20775 36261
rect 20824 36236 20852 36332
rect 17000 36196 17172 36224
rect 17236 36196 17816 36224
rect 17000 36184 17006 36196
rect 17144 36165 17172 36196
rect 16531 36128 16896 36156
rect 17037 36159 17095 36165
rect 16531 36125 16543 36128
rect 16485 36119 16543 36125
rect 17037 36125 17049 36159
rect 17083 36125 17095 36159
rect 17037 36119 17095 36125
rect 17129 36159 17187 36165
rect 17129 36125 17141 36159
rect 17175 36125 17187 36159
rect 17129 36119 17187 36125
rect 16408 36088 16436 36119
rect 17052 36088 17080 36119
rect 17218 36116 17224 36168
rect 17276 36116 17282 36168
rect 17405 36159 17463 36165
rect 17405 36125 17417 36159
rect 17451 36156 17463 36159
rect 17494 36156 17500 36168
rect 17451 36128 17500 36156
rect 17451 36125 17463 36128
rect 17405 36119 17463 36125
rect 17494 36116 17500 36128
rect 17552 36116 17558 36168
rect 17788 36165 17816 36196
rect 17862 36184 17868 36236
rect 17920 36224 17926 36236
rect 18049 36227 18107 36233
rect 18049 36224 18061 36227
rect 17920 36196 18061 36224
rect 17920 36184 17926 36196
rect 18049 36193 18061 36196
rect 18095 36193 18107 36227
rect 18598 36224 18604 36236
rect 18049 36187 18107 36193
rect 18248 36196 18604 36224
rect 17681 36159 17739 36165
rect 17681 36125 17693 36159
rect 17727 36125 17739 36159
rect 17681 36119 17739 36125
rect 17773 36159 17831 36165
rect 17773 36125 17785 36159
rect 17819 36156 17831 36159
rect 18248 36156 18276 36196
rect 18598 36184 18604 36196
rect 18656 36224 18662 36236
rect 19150 36224 19156 36236
rect 18656 36196 19156 36224
rect 18656 36184 18662 36196
rect 19150 36184 19156 36196
rect 19208 36184 19214 36236
rect 20622 36184 20628 36236
rect 20680 36224 20686 36236
rect 20806 36224 20812 36236
rect 20680 36196 20812 36224
rect 20680 36184 20686 36196
rect 20806 36184 20812 36196
rect 20864 36184 20870 36236
rect 17819 36128 18276 36156
rect 17819 36125 17831 36128
rect 17773 36119 17831 36125
rect 17696 36088 17724 36119
rect 18690 36116 18696 36168
rect 18748 36116 18754 36168
rect 18877 36159 18935 36165
rect 18877 36125 18889 36159
rect 18923 36125 18935 36159
rect 18877 36119 18935 36125
rect 17862 36088 17868 36100
rect 16408 36060 16804 36088
rect 17052 36060 17868 36088
rect 16482 36020 16488 36032
rect 16316 35992 16488 36020
rect 16482 35980 16488 35992
rect 16540 35980 16546 36032
rect 16666 35980 16672 36032
rect 16724 35980 16730 36032
rect 16776 36020 16804 36060
rect 17862 36048 17868 36060
rect 17920 36048 17926 36100
rect 17957 36091 18015 36097
rect 17957 36057 17969 36091
rect 18003 36088 18015 36091
rect 18892 36088 18920 36119
rect 19886 36116 19892 36168
rect 19944 36116 19950 36168
rect 20073 36159 20131 36165
rect 20073 36125 20085 36159
rect 20119 36156 20131 36159
rect 20257 36159 20315 36165
rect 20119 36128 20208 36156
rect 20119 36125 20131 36128
rect 20073 36119 20131 36125
rect 18003 36060 18920 36088
rect 18003 36057 18015 36060
rect 17957 36051 18015 36057
rect 20180 36032 20208 36128
rect 20257 36125 20269 36159
rect 20303 36125 20315 36159
rect 20257 36119 20315 36125
rect 20349 36159 20407 36165
rect 20349 36125 20361 36159
rect 20395 36125 20407 36159
rect 20349 36119 20407 36125
rect 20441 36159 20499 36165
rect 20441 36125 20453 36159
rect 20487 36156 20499 36159
rect 20714 36156 20720 36168
rect 20487 36128 20720 36156
rect 20487 36125 20499 36128
rect 20441 36119 20499 36125
rect 18414 36020 18420 36032
rect 16776 35992 18420 36020
rect 18414 35980 18420 35992
rect 18472 35980 18478 36032
rect 20162 35980 20168 36032
rect 20220 35980 20226 36032
rect 20272 36020 20300 36119
rect 20364 36088 20392 36119
rect 20714 36116 20720 36128
rect 20772 36116 20778 36168
rect 22066 36156 22094 36332
rect 23198 36156 23204 36168
rect 22066 36128 23204 36156
rect 23198 36116 23204 36128
rect 23256 36156 23262 36168
rect 23753 36159 23811 36165
rect 23753 36156 23765 36159
rect 23256 36128 23765 36156
rect 23256 36116 23262 36128
rect 23753 36125 23765 36128
rect 23799 36125 23811 36159
rect 23753 36119 23811 36125
rect 21076 36091 21134 36097
rect 20364 36060 21045 36088
rect 20898 36020 20904 36032
rect 20272 35992 20904 36020
rect 20898 35980 20904 35992
rect 20956 35980 20962 36032
rect 21017 36020 21045 36060
rect 21076 36057 21088 36091
rect 21122 36088 21134 36091
rect 21358 36088 21364 36100
rect 21122 36060 21364 36088
rect 21122 36057 21134 36060
rect 21076 36051 21134 36057
rect 21358 36048 21364 36060
rect 21416 36048 21422 36100
rect 23508 36091 23566 36097
rect 23508 36057 23520 36091
rect 23554 36088 23566 36091
rect 23842 36088 23848 36100
rect 23554 36060 23848 36088
rect 23554 36057 23566 36060
rect 23508 36051 23566 36057
rect 23842 36048 23848 36060
rect 23900 36048 23906 36100
rect 21818 36020 21824 36032
rect 21017 35992 21824 36020
rect 21818 35980 21824 35992
rect 21876 35980 21882 36032
rect 22186 35980 22192 36032
rect 22244 35980 22250 36032
rect 22278 35980 22284 36032
rect 22336 36020 22342 36032
rect 22373 36023 22431 36029
rect 22373 36020 22385 36023
rect 22336 35992 22385 36020
rect 22336 35980 22342 35992
rect 22373 35989 22385 35992
rect 22419 35989 22431 36023
rect 22373 35983 22431 35989
rect 1104 35930 35027 35952
rect 1104 35878 9390 35930
rect 9442 35878 9454 35930
rect 9506 35878 9518 35930
rect 9570 35878 9582 35930
rect 9634 35878 9646 35930
rect 9698 35878 17831 35930
rect 17883 35878 17895 35930
rect 17947 35878 17959 35930
rect 18011 35878 18023 35930
rect 18075 35878 18087 35930
rect 18139 35878 26272 35930
rect 26324 35878 26336 35930
rect 26388 35878 26400 35930
rect 26452 35878 26464 35930
rect 26516 35878 26528 35930
rect 26580 35878 34713 35930
rect 34765 35878 34777 35930
rect 34829 35878 34841 35930
rect 34893 35878 34905 35930
rect 34957 35878 34969 35930
rect 35021 35878 35027 35930
rect 1104 35856 35027 35878
rect 8941 35819 8999 35825
rect 8941 35785 8953 35819
rect 8987 35785 8999 35819
rect 9766 35816 9772 35828
rect 8941 35779 8999 35785
rect 9416 35788 9772 35816
rect 8754 35640 8760 35692
rect 8812 35640 8818 35692
rect 8846 35640 8852 35692
rect 8904 35640 8910 35692
rect 8956 35680 8984 35779
rect 9416 35757 9444 35788
rect 9766 35776 9772 35788
rect 9824 35776 9830 35828
rect 10965 35819 11023 35825
rect 10965 35785 10977 35819
rect 11011 35816 11023 35819
rect 11146 35816 11152 35828
rect 11011 35788 11152 35816
rect 11011 35785 11023 35788
rect 10965 35779 11023 35785
rect 11146 35776 11152 35788
rect 11204 35776 11210 35828
rect 11790 35776 11796 35828
rect 11848 35816 11854 35828
rect 12526 35816 12532 35828
rect 11848 35788 12532 35816
rect 11848 35776 11854 35788
rect 9401 35751 9459 35757
rect 9401 35717 9413 35751
rect 9447 35717 9459 35751
rect 12161 35751 12219 35757
rect 12161 35748 12173 35751
rect 9401 35711 9459 35717
rect 11164 35720 12173 35748
rect 11164 35689 11192 35720
rect 12161 35717 12173 35720
rect 12207 35717 12219 35751
rect 12161 35711 12219 35717
rect 9841 35683 9899 35689
rect 9841 35680 9853 35683
rect 8956 35652 9853 35680
rect 9841 35649 9853 35652
rect 9887 35649 9899 35683
rect 9841 35643 9899 35649
rect 11149 35683 11207 35689
rect 11149 35649 11161 35683
rect 11195 35649 11207 35683
rect 11882 35680 11888 35692
rect 11149 35643 11207 35649
rect 11256 35652 11888 35680
rect 8864 35612 8892 35640
rect 9306 35612 9312 35624
rect 8864 35584 9312 35612
rect 9306 35572 9312 35584
rect 9364 35612 9370 35624
rect 9585 35615 9643 35621
rect 9585 35612 9597 35615
rect 9364 35584 9597 35612
rect 9364 35572 9370 35584
rect 9585 35581 9597 35584
rect 9631 35581 9643 35615
rect 9585 35575 9643 35581
rect 9309 35479 9367 35485
rect 9309 35445 9321 35479
rect 9355 35476 9367 35479
rect 11256 35476 11284 35652
rect 11882 35640 11888 35652
rect 11940 35640 11946 35692
rect 12360 35689 12388 35788
rect 12526 35776 12532 35788
rect 12584 35776 12590 35828
rect 13170 35816 13176 35828
rect 12820 35788 13176 35816
rect 12820 35689 12848 35788
rect 13170 35776 13176 35788
rect 13228 35776 13234 35828
rect 13265 35819 13323 35825
rect 13265 35785 13277 35819
rect 13311 35816 13323 35819
rect 13446 35816 13452 35828
rect 13311 35788 13452 35816
rect 13311 35785 13323 35788
rect 13265 35779 13323 35785
rect 13446 35776 13452 35788
rect 13504 35776 13510 35828
rect 13630 35776 13636 35828
rect 13688 35776 13694 35828
rect 16666 35776 16672 35828
rect 16724 35776 16730 35828
rect 18690 35776 18696 35828
rect 18748 35816 18754 35828
rect 19061 35819 19119 35825
rect 19061 35816 19073 35819
rect 18748 35788 19073 35816
rect 18748 35776 18754 35788
rect 19061 35785 19073 35788
rect 19107 35785 19119 35819
rect 19061 35779 19119 35785
rect 20438 35776 20444 35828
rect 20496 35776 20502 35828
rect 20530 35776 20536 35828
rect 20588 35776 20594 35828
rect 21082 35776 21088 35828
rect 21140 35776 21146 35828
rect 21358 35776 21364 35828
rect 21416 35776 21422 35828
rect 21818 35776 21824 35828
rect 21876 35776 21882 35828
rect 22462 35776 22468 35828
rect 22520 35776 22526 35828
rect 23842 35776 23848 35828
rect 23900 35776 23906 35828
rect 24305 35819 24363 35825
rect 24305 35785 24317 35819
rect 24351 35816 24363 35819
rect 24486 35816 24492 35828
rect 24351 35788 24492 35816
rect 24351 35785 24363 35788
rect 24305 35779 24363 35785
rect 24486 35776 24492 35788
rect 24544 35776 24550 35828
rect 13648 35748 13676 35776
rect 12912 35720 13676 35748
rect 14476 35720 16344 35748
rect 12912 35689 12940 35720
rect 12345 35683 12403 35689
rect 12345 35649 12357 35683
rect 12391 35649 12403 35683
rect 12345 35643 12403 35649
rect 12621 35683 12679 35689
rect 12621 35649 12633 35683
rect 12667 35649 12679 35683
rect 12621 35643 12679 35649
rect 12805 35683 12863 35689
rect 12805 35649 12817 35683
rect 12851 35649 12863 35683
rect 12805 35643 12863 35649
rect 12897 35683 12955 35689
rect 12897 35649 12909 35683
rect 12943 35649 12955 35683
rect 12897 35643 12955 35649
rect 12434 35572 12440 35624
rect 12492 35612 12498 35624
rect 12529 35615 12587 35621
rect 12529 35612 12541 35615
rect 12492 35584 12541 35612
rect 12492 35572 12498 35584
rect 12529 35581 12541 35584
rect 12575 35581 12587 35615
rect 12636 35612 12664 35643
rect 12986 35640 12992 35692
rect 13044 35640 13050 35692
rect 14090 35680 14096 35692
rect 13096 35652 14096 35680
rect 13096 35612 13124 35652
rect 14090 35640 14096 35652
rect 14148 35640 14154 35692
rect 14476 35689 14504 35720
rect 14461 35683 14519 35689
rect 14461 35649 14473 35683
rect 14507 35649 14519 35683
rect 14461 35643 14519 35649
rect 14553 35683 14611 35689
rect 14553 35649 14565 35683
rect 14599 35649 14611 35683
rect 14553 35643 14611 35649
rect 15096 35683 15154 35689
rect 15096 35649 15108 35683
rect 15142 35680 15154 35683
rect 16022 35680 16028 35692
rect 15142 35652 16028 35680
rect 15142 35649 15154 35652
rect 15096 35643 15154 35649
rect 12636 35584 13124 35612
rect 12529 35575 12587 35581
rect 13354 35572 13360 35624
rect 13412 35612 13418 35624
rect 13909 35615 13967 35621
rect 13909 35612 13921 35615
rect 13412 35584 13921 35612
rect 13412 35572 13418 35584
rect 13909 35581 13921 35584
rect 13955 35581 13967 35615
rect 14568 35612 14596 35643
rect 16022 35640 16028 35652
rect 16080 35640 16086 35692
rect 13909 35575 13967 35581
rect 14016 35584 14596 35612
rect 14829 35615 14887 35621
rect 11606 35504 11612 35556
rect 11664 35544 11670 35556
rect 11793 35547 11851 35553
rect 11793 35544 11805 35547
rect 11664 35516 11805 35544
rect 11664 35504 11670 35516
rect 11793 35513 11805 35516
rect 11839 35513 11851 35547
rect 11793 35507 11851 35513
rect 13078 35504 13084 35556
rect 13136 35544 13142 35556
rect 14016 35544 14044 35584
rect 14829 35581 14841 35615
rect 14875 35581 14887 35615
rect 14829 35575 14887 35581
rect 13136 35516 14044 35544
rect 13136 35504 13142 35516
rect 14550 35504 14556 35556
rect 14608 35544 14614 35556
rect 14844 35544 14872 35575
rect 16316 35556 16344 35720
rect 16684 35680 16712 35776
rect 16758 35708 16764 35760
rect 16816 35748 16822 35760
rect 17310 35748 17316 35760
rect 16816 35720 17316 35748
rect 16816 35708 16822 35720
rect 17310 35708 17316 35720
rect 17368 35708 17374 35760
rect 18966 35748 18972 35760
rect 17696 35720 18972 35748
rect 17696 35692 17724 35720
rect 18966 35708 18972 35720
rect 19024 35748 19030 35760
rect 19420 35751 19478 35757
rect 19024 35720 19196 35748
rect 19024 35708 19030 35720
rect 17405 35683 17463 35689
rect 17405 35680 17417 35683
rect 16684 35652 17417 35680
rect 17405 35649 17417 35652
rect 17451 35649 17463 35683
rect 17405 35643 17463 35649
rect 17678 35640 17684 35692
rect 17736 35640 17742 35692
rect 19168 35689 19196 35720
rect 19420 35717 19432 35751
rect 19466 35748 19478 35751
rect 20070 35748 20076 35760
rect 19466 35720 20076 35748
rect 19466 35717 19478 35720
rect 19420 35711 19478 35717
rect 20070 35708 20076 35720
rect 20128 35708 20134 35760
rect 17937 35683 17995 35689
rect 17937 35680 17949 35683
rect 17788 35652 17949 35680
rect 17788 35612 17816 35652
rect 17937 35649 17949 35652
rect 17983 35649 17995 35683
rect 17937 35643 17995 35649
rect 19153 35683 19211 35689
rect 19153 35649 19165 35683
rect 19199 35649 19211 35683
rect 20456 35680 20484 35776
rect 20625 35683 20683 35689
rect 20625 35680 20637 35683
rect 20456 35652 20637 35680
rect 19153 35643 19211 35649
rect 20625 35649 20637 35652
rect 20671 35649 20683 35683
rect 21100 35680 21128 35776
rect 22480 35748 22508 35776
rect 21836 35720 22140 35748
rect 21545 35683 21603 35689
rect 21545 35680 21557 35683
rect 21100 35652 21557 35680
rect 20625 35643 20683 35649
rect 21545 35649 21557 35652
rect 21591 35649 21603 35683
rect 21545 35643 21603 35649
rect 17604 35584 17816 35612
rect 14608 35516 14872 35544
rect 14608 35504 14614 35516
rect 16298 35504 16304 35556
rect 16356 35544 16362 35556
rect 17604 35553 17632 35584
rect 17037 35547 17095 35553
rect 17037 35544 17049 35547
rect 16356 35516 17049 35544
rect 16356 35504 16362 35516
rect 17037 35513 17049 35516
rect 17083 35513 17095 35547
rect 17037 35507 17095 35513
rect 17589 35547 17647 35553
rect 17589 35513 17601 35547
rect 17635 35513 17647 35547
rect 17589 35507 17647 35513
rect 21836 35488 21864 35720
rect 22112 35689 22140 35720
rect 22204 35720 22508 35748
rect 22204 35689 22232 35720
rect 22097 35683 22155 35689
rect 22097 35649 22109 35683
rect 22143 35649 22155 35683
rect 22097 35643 22155 35649
rect 22189 35683 22247 35689
rect 22189 35649 22201 35683
rect 22235 35649 22247 35683
rect 22189 35643 22247 35649
rect 22278 35640 22284 35692
rect 22336 35680 22342 35692
rect 22373 35683 22431 35689
rect 22373 35680 22385 35683
rect 22336 35652 22385 35680
rect 22336 35640 22342 35652
rect 22373 35649 22385 35652
rect 22419 35680 22431 35683
rect 22462 35680 22468 35692
rect 22419 35652 22468 35680
rect 22419 35649 22431 35652
rect 22373 35643 22431 35649
rect 22462 35640 22468 35652
rect 22520 35640 22526 35692
rect 22557 35683 22615 35689
rect 22557 35649 22569 35683
rect 22603 35649 22615 35683
rect 22557 35643 22615 35649
rect 23569 35683 23627 35689
rect 23569 35649 23581 35683
rect 23615 35649 23627 35683
rect 23569 35643 23627 35649
rect 23753 35683 23811 35689
rect 23753 35649 23765 35683
rect 23799 35680 23811 35683
rect 24029 35683 24087 35689
rect 24029 35680 24041 35683
rect 23799 35652 24041 35680
rect 23799 35649 23811 35652
rect 23753 35643 23811 35649
rect 24029 35649 24041 35652
rect 24075 35649 24087 35683
rect 24029 35643 24087 35649
rect 21910 35572 21916 35624
rect 21968 35612 21974 35624
rect 22572 35612 22600 35643
rect 21968 35584 22600 35612
rect 22649 35615 22707 35621
rect 21968 35572 21974 35584
rect 22649 35581 22661 35615
rect 22695 35581 22707 35615
rect 22649 35575 22707 35581
rect 23293 35615 23351 35621
rect 23293 35581 23305 35615
rect 23339 35612 23351 35615
rect 23385 35615 23443 35621
rect 23385 35612 23397 35615
rect 23339 35584 23397 35612
rect 23339 35581 23351 35584
rect 23293 35575 23351 35581
rect 23385 35581 23397 35584
rect 23431 35581 23443 35615
rect 23385 35575 23443 35581
rect 22186 35504 22192 35556
rect 22244 35544 22250 35556
rect 22281 35547 22339 35553
rect 22281 35544 22293 35547
rect 22244 35516 22293 35544
rect 22244 35504 22250 35516
rect 22281 35513 22293 35516
rect 22327 35544 22339 35547
rect 22554 35544 22560 35556
rect 22327 35516 22560 35544
rect 22327 35513 22339 35516
rect 22281 35507 22339 35513
rect 22554 35504 22560 35516
rect 22612 35544 22618 35556
rect 22664 35544 22692 35575
rect 22612 35516 22692 35544
rect 22612 35504 22618 35516
rect 9355 35448 11284 35476
rect 11333 35479 11391 35485
rect 9355 35445 9367 35448
rect 9309 35439 9367 35445
rect 11333 35445 11345 35479
rect 11379 35476 11391 35479
rect 11698 35476 11704 35488
rect 11379 35448 11704 35476
rect 11379 35445 11391 35448
rect 11333 35439 11391 35445
rect 11698 35436 11704 35448
rect 11756 35436 11762 35488
rect 12986 35436 12992 35488
rect 13044 35476 13050 35488
rect 13357 35479 13415 35485
rect 13357 35476 13369 35479
rect 13044 35448 13369 35476
rect 13044 35436 13050 35448
rect 13357 35445 13369 35448
rect 13403 35445 13415 35479
rect 13357 35439 13415 35445
rect 14734 35436 14740 35488
rect 14792 35436 14798 35488
rect 16114 35436 16120 35488
rect 16172 35476 16178 35488
rect 16209 35479 16267 35485
rect 16209 35476 16221 35479
rect 16172 35448 16221 35476
rect 16172 35436 16178 35448
rect 16209 35445 16221 35448
rect 16255 35445 16267 35479
rect 16209 35439 16267 35445
rect 17218 35436 17224 35488
rect 17276 35436 17282 35488
rect 21266 35436 21272 35488
rect 21324 35436 21330 35488
rect 21818 35436 21824 35488
rect 21876 35436 21882 35488
rect 22646 35436 22652 35488
rect 22704 35476 22710 35488
rect 23584 35476 23612 35643
rect 24118 35640 24124 35692
rect 24176 35640 24182 35692
rect 22704 35448 23612 35476
rect 22704 35436 22710 35448
rect 1104 35386 34868 35408
rect 1104 35334 5170 35386
rect 5222 35334 5234 35386
rect 5286 35334 5298 35386
rect 5350 35334 5362 35386
rect 5414 35334 5426 35386
rect 5478 35334 13611 35386
rect 13663 35334 13675 35386
rect 13727 35334 13739 35386
rect 13791 35334 13803 35386
rect 13855 35334 13867 35386
rect 13919 35334 22052 35386
rect 22104 35334 22116 35386
rect 22168 35334 22180 35386
rect 22232 35334 22244 35386
rect 22296 35334 22308 35386
rect 22360 35334 30493 35386
rect 30545 35334 30557 35386
rect 30609 35334 30621 35386
rect 30673 35334 30685 35386
rect 30737 35334 30749 35386
rect 30801 35334 34868 35386
rect 1104 35312 34868 35334
rect 8754 35232 8760 35284
rect 8812 35272 8818 35284
rect 10873 35275 10931 35281
rect 10873 35272 10885 35275
rect 8812 35244 10885 35272
rect 8812 35232 8818 35244
rect 10873 35241 10885 35244
rect 10919 35241 10931 35275
rect 10873 35235 10931 35241
rect 12437 35275 12495 35281
rect 12437 35241 12449 35275
rect 12483 35272 12495 35275
rect 12483 35244 14320 35272
rect 12483 35241 12495 35244
rect 12437 35235 12495 35241
rect 10778 35164 10784 35216
rect 10836 35164 10842 35216
rect 14093 35207 14151 35213
rect 14093 35173 14105 35207
rect 14139 35173 14151 35207
rect 14093 35167 14151 35173
rect 9306 35096 9312 35148
rect 9364 35136 9370 35148
rect 9401 35139 9459 35145
rect 9401 35136 9413 35139
rect 9364 35108 9413 35136
rect 9364 35096 9370 35108
rect 9401 35105 9413 35108
rect 9447 35105 9459 35139
rect 9401 35099 9459 35105
rect 12069 35139 12127 35145
rect 12069 35105 12081 35139
rect 12115 35136 12127 35139
rect 12894 35136 12900 35148
rect 12115 35108 12900 35136
rect 12115 35105 12127 35108
rect 12069 35099 12127 35105
rect 12894 35096 12900 35108
rect 12952 35096 12958 35148
rect 14108 35136 14136 35167
rect 13832 35108 14136 35136
rect 9668 35071 9726 35077
rect 9668 35037 9680 35071
rect 9714 35068 9726 35071
rect 9950 35068 9956 35080
rect 9714 35040 9956 35068
rect 9714 35037 9726 35040
rect 9668 35031 9726 35037
rect 9950 35028 9956 35040
rect 10008 35028 10014 35080
rect 11057 35071 11115 35077
rect 11057 35037 11069 35071
rect 11103 35037 11115 35071
rect 11057 35031 11115 35037
rect 10042 34960 10048 35012
rect 10100 35000 10106 35012
rect 11072 35000 11100 35031
rect 11238 35028 11244 35080
rect 11296 35028 11302 35080
rect 11330 35028 11336 35080
rect 11388 35028 11394 35080
rect 11514 35068 11520 35080
rect 11440 35040 11520 35068
rect 11440 35000 11468 35040
rect 11514 35028 11520 35040
rect 11572 35028 11578 35080
rect 11606 35028 11612 35080
rect 11664 35028 11670 35080
rect 11790 35028 11796 35080
rect 11848 35068 11854 35080
rect 12253 35071 12311 35077
rect 11848 35064 12112 35068
rect 12253 35064 12265 35071
rect 11848 35040 12265 35064
rect 11848 35028 11854 35040
rect 12084 35037 12265 35040
rect 12299 35037 12311 35071
rect 12084 35036 12311 35037
rect 12253 35031 12311 35036
rect 12618 35000 12624 35012
rect 10100 34972 11468 35000
rect 11532 34972 12624 35000
rect 10100 34960 10106 34972
rect 11532 34941 11560 34972
rect 12618 34960 12624 34972
rect 12676 34960 12682 35012
rect 13664 35003 13722 35009
rect 13664 34969 13676 35003
rect 13710 35000 13722 35003
rect 13832 35000 13860 35108
rect 13909 35071 13967 35077
rect 13909 35037 13921 35071
rect 13955 35068 13967 35071
rect 13998 35068 14004 35080
rect 13955 35040 14004 35068
rect 13955 35037 13967 35040
rect 13909 35031 13967 35037
rect 13998 35028 14004 35040
rect 14056 35068 14062 35080
rect 14292 35077 14320 35244
rect 16114 35232 16120 35284
rect 16172 35232 16178 35284
rect 17218 35232 17224 35284
rect 17276 35232 17282 35284
rect 17402 35232 17408 35284
rect 17460 35272 17466 35284
rect 19061 35275 19119 35281
rect 19061 35272 19073 35275
rect 17460 35244 19073 35272
rect 17460 35232 17466 35244
rect 19061 35241 19073 35244
rect 19107 35241 19119 35275
rect 19061 35235 19119 35241
rect 19886 35232 19892 35284
rect 19944 35272 19950 35284
rect 20257 35275 20315 35281
rect 20257 35272 20269 35275
rect 19944 35244 20269 35272
rect 19944 35232 19950 35244
rect 20257 35241 20269 35244
rect 20303 35241 20315 35275
rect 20257 35235 20315 35241
rect 15933 35207 15991 35213
rect 15933 35173 15945 35207
rect 15979 35173 15991 35207
rect 15933 35167 15991 35173
rect 14550 35096 14556 35148
rect 14608 35096 14614 35148
rect 14277 35071 14335 35077
rect 14056 35040 14228 35068
rect 14056 35028 14062 35040
rect 13710 34972 13860 35000
rect 14200 35000 14228 35040
rect 14277 35037 14289 35071
rect 14323 35037 14335 35071
rect 14277 35031 14335 35037
rect 14568 35000 14596 35096
rect 15948 35068 15976 35167
rect 16025 35139 16083 35145
rect 16025 35105 16037 35139
rect 16071 35136 16083 35139
rect 16132 35136 16160 35232
rect 17037 35207 17095 35213
rect 17037 35173 17049 35207
rect 17083 35204 17095 35207
rect 17236 35204 17264 35232
rect 17083 35176 18828 35204
rect 17083 35173 17095 35176
rect 17037 35167 17095 35173
rect 17129 35139 17187 35145
rect 16071 35108 16160 35136
rect 16776 35108 16988 35136
rect 16071 35105 16083 35108
rect 16025 35099 16083 35105
rect 16209 35071 16267 35077
rect 16209 35068 16221 35071
rect 15948 35040 16221 35068
rect 16209 35037 16221 35040
rect 16255 35068 16267 35071
rect 16298 35068 16304 35080
rect 16255 35040 16304 35068
rect 16255 35037 16267 35040
rect 16209 35031 16267 35037
rect 16298 35028 16304 35040
rect 16356 35028 16362 35080
rect 16776 35077 16804 35108
rect 16393 35071 16451 35077
rect 16393 35037 16405 35071
rect 16439 35068 16451 35071
rect 16761 35071 16819 35077
rect 16761 35068 16773 35071
rect 16439 35040 16773 35068
rect 16439 35037 16451 35040
rect 16393 35031 16451 35037
rect 16761 35037 16773 35040
rect 16807 35037 16819 35071
rect 16761 35031 16819 35037
rect 16853 35071 16911 35077
rect 16853 35037 16865 35071
rect 16899 35037 16911 35071
rect 16960 35068 16988 35108
rect 17129 35105 17141 35139
rect 17175 35136 17187 35139
rect 17218 35136 17224 35148
rect 17175 35108 17224 35136
rect 17175 35105 17187 35108
rect 17129 35099 17187 35105
rect 17218 35096 17224 35108
rect 17276 35136 17282 35148
rect 18601 35139 18659 35145
rect 17276 35108 18552 35136
rect 17276 35096 17282 35108
rect 16960 35040 17264 35068
rect 16853 35031 16911 35037
rect 14200 34972 14596 35000
rect 14820 35003 14878 35009
rect 13710 34969 13722 34972
rect 13664 34963 13722 34969
rect 14820 34969 14832 35003
rect 14866 35000 14878 35003
rect 15010 35000 15016 35012
rect 14866 34972 15016 35000
rect 14866 34969 14878 34972
rect 14820 34963 14878 34969
rect 15010 34960 15016 34972
rect 15068 34960 15074 35012
rect 16868 34944 16896 35031
rect 17236 35000 17264 35040
rect 17678 35028 17684 35080
rect 17736 35068 17742 35080
rect 17773 35071 17831 35077
rect 17773 35068 17785 35071
rect 17736 35040 17785 35068
rect 17736 35028 17742 35040
rect 17773 35037 17785 35040
rect 17819 35037 17831 35071
rect 17773 35031 17831 35037
rect 18414 35028 18420 35080
rect 18472 35028 18478 35080
rect 18524 35077 18552 35108
rect 18601 35105 18613 35139
rect 18647 35105 18659 35139
rect 18601 35099 18659 35105
rect 18509 35071 18567 35077
rect 18509 35037 18521 35071
rect 18555 35037 18567 35071
rect 18509 35031 18567 35037
rect 18616 35000 18644 35099
rect 18800 35077 18828 35176
rect 18874 35164 18880 35216
rect 18932 35204 18938 35216
rect 19705 35207 19763 35213
rect 19705 35204 19717 35207
rect 18932 35176 19717 35204
rect 18932 35164 18938 35176
rect 19705 35173 19717 35176
rect 19751 35173 19763 35207
rect 19705 35167 19763 35173
rect 18785 35071 18843 35077
rect 18785 35037 18797 35071
rect 18831 35037 18843 35071
rect 18785 35031 18843 35037
rect 18877 35071 18935 35077
rect 18877 35037 18889 35071
rect 18923 35037 18935 35071
rect 18877 35031 18935 35037
rect 17236 34972 18644 35000
rect 11517 34935 11575 34941
rect 11517 34901 11529 34935
rect 11563 34901 11575 34935
rect 11517 34895 11575 34901
rect 11793 34935 11851 34941
rect 11793 34901 11805 34935
rect 11839 34932 11851 34935
rect 12250 34932 12256 34944
rect 11839 34904 12256 34932
rect 11839 34901 11851 34904
rect 11793 34895 11851 34901
rect 12250 34892 12256 34904
rect 12308 34892 12314 34944
rect 12529 34935 12587 34941
rect 12529 34901 12541 34935
rect 12575 34932 12587 34935
rect 12710 34932 12716 34944
rect 12575 34904 12716 34932
rect 12575 34901 12587 34904
rect 12529 34895 12587 34901
rect 12710 34892 12716 34904
rect 12768 34892 12774 34944
rect 15102 34892 15108 34944
rect 15160 34932 15166 34944
rect 16577 34935 16635 34941
rect 16577 34932 16589 34935
rect 15160 34904 16589 34932
rect 15160 34892 15166 34904
rect 16577 34901 16589 34904
rect 16623 34901 16635 34935
rect 16577 34895 16635 34901
rect 16850 34892 16856 34944
rect 16908 34932 16914 34944
rect 18892 34932 18920 35031
rect 19058 35028 19064 35080
rect 19116 35068 19122 35080
rect 19889 35071 19947 35077
rect 19889 35068 19901 35071
rect 19116 35040 19901 35068
rect 19116 35028 19122 35040
rect 19889 35037 19901 35040
rect 19935 35037 19947 35071
rect 19889 35031 19947 35037
rect 16908 34904 18920 34932
rect 20272 34932 20300 35235
rect 20898 35232 20904 35284
rect 20956 35272 20962 35284
rect 21729 35275 21787 35281
rect 21729 35272 21741 35275
rect 20956 35244 21741 35272
rect 20956 35232 20962 35244
rect 21729 35241 21741 35244
rect 21775 35241 21787 35275
rect 21729 35235 21787 35241
rect 21910 35232 21916 35284
rect 21968 35232 21974 35284
rect 22554 35272 22560 35284
rect 22296 35244 22560 35272
rect 21928 35136 21956 35232
rect 22296 35145 22324 35244
rect 22554 35232 22560 35244
rect 22612 35232 22618 35284
rect 23845 35275 23903 35281
rect 23845 35241 23857 35275
rect 23891 35272 23903 35275
rect 24118 35272 24124 35284
rect 23891 35244 24124 35272
rect 23891 35241 23903 35244
rect 23845 35235 23903 35241
rect 24118 35232 24124 35244
rect 24176 35232 24182 35284
rect 22005 35139 22063 35145
rect 22005 35136 22017 35139
rect 21928 35108 22017 35136
rect 22005 35105 22017 35108
rect 22051 35105 22063 35139
rect 22005 35099 22063 35105
rect 22281 35139 22339 35145
rect 22281 35105 22293 35139
rect 22327 35105 22339 35139
rect 22281 35099 22339 35105
rect 22370 35096 22376 35148
rect 22428 35096 22434 35148
rect 20806 35028 20812 35080
rect 20864 35068 20870 35080
rect 21637 35071 21695 35077
rect 21637 35068 21649 35071
rect 20864 35040 21649 35068
rect 20864 35028 20870 35040
rect 21637 35037 21649 35040
rect 21683 35037 21695 35071
rect 21637 35031 21695 35037
rect 21818 35028 21824 35080
rect 21876 35068 21882 35080
rect 21913 35071 21971 35077
rect 21913 35068 21925 35071
rect 21876 35040 21925 35068
rect 21876 35028 21882 35040
rect 21913 35037 21925 35040
rect 21959 35037 21971 35071
rect 21913 35031 21971 35037
rect 21266 34960 21272 35012
rect 21324 35000 21330 35012
rect 21370 35003 21428 35009
rect 21370 35000 21382 35003
rect 21324 34972 21382 35000
rect 21324 34960 21330 34972
rect 21370 34969 21382 34972
rect 21416 34969 21428 35003
rect 21370 34963 21428 34969
rect 21928 34932 21956 35031
rect 22462 35028 22468 35080
rect 22520 35028 22526 35080
rect 22554 35028 22560 35080
rect 22612 35028 22618 35080
rect 23566 35028 23572 35080
rect 23624 35028 23630 35080
rect 23661 35071 23719 35077
rect 23661 35037 23673 35071
rect 23707 35068 23719 35071
rect 34517 35071 34575 35077
rect 23707 35040 31754 35068
rect 23707 35037 23719 35040
rect 23661 35031 23719 35037
rect 22480 35000 22508 35028
rect 22204 34972 22508 35000
rect 22204 34941 22232 34972
rect 20272 34904 21956 34932
rect 22189 34935 22247 34941
rect 16908 34892 16914 34904
rect 22189 34901 22201 34935
rect 22235 34901 22247 34935
rect 22189 34895 22247 34901
rect 22738 34892 22744 34944
rect 22796 34892 22802 34944
rect 31726 34932 31754 35040
rect 34517 35037 34529 35071
rect 34563 35068 34575 35071
rect 34563 35040 35204 35068
rect 34563 35037 34575 35040
rect 34517 35031 34575 35037
rect 35176 34944 35204 35040
rect 34333 34935 34391 34941
rect 34333 34932 34345 34935
rect 31726 34904 34345 34932
rect 34333 34901 34345 34904
rect 34379 34901 34391 34935
rect 34333 34895 34391 34901
rect 35158 34892 35164 34944
rect 35216 34892 35222 34944
rect 1104 34842 35027 34864
rect 1104 34790 9390 34842
rect 9442 34790 9454 34842
rect 9506 34790 9518 34842
rect 9570 34790 9582 34842
rect 9634 34790 9646 34842
rect 9698 34790 17831 34842
rect 17883 34790 17895 34842
rect 17947 34790 17959 34842
rect 18011 34790 18023 34842
rect 18075 34790 18087 34842
rect 18139 34790 26272 34842
rect 26324 34790 26336 34842
rect 26388 34790 26400 34842
rect 26452 34790 26464 34842
rect 26516 34790 26528 34842
rect 26580 34790 34713 34842
rect 34765 34790 34777 34842
rect 34829 34790 34841 34842
rect 34893 34790 34905 34842
rect 34957 34790 34969 34842
rect 35021 34790 35027 34842
rect 1104 34768 35027 34790
rect 9493 34731 9551 34737
rect 9493 34697 9505 34731
rect 9539 34728 9551 34731
rect 10042 34728 10048 34740
rect 9539 34700 10048 34728
rect 9539 34697 9551 34700
rect 9493 34691 9551 34697
rect 10042 34688 10048 34700
rect 10100 34688 10106 34740
rect 10137 34731 10195 34737
rect 10137 34697 10149 34731
rect 10183 34728 10195 34731
rect 11238 34728 11244 34740
rect 10183 34700 11244 34728
rect 10183 34697 10195 34700
rect 10137 34691 10195 34697
rect 11238 34688 11244 34700
rect 11296 34688 11302 34740
rect 11330 34688 11336 34740
rect 11388 34688 11394 34740
rect 11532 34700 12388 34728
rect 9692 34632 11100 34660
rect 9125 34595 9183 34601
rect 9125 34592 9137 34595
rect 8588 34564 9137 34592
rect 8588 34536 8616 34564
rect 9125 34561 9137 34564
rect 9171 34561 9183 34595
rect 9125 34555 9183 34561
rect 8570 34484 8576 34536
rect 8628 34484 8634 34536
rect 9140 34524 9168 34555
rect 9214 34552 9220 34604
rect 9272 34552 9278 34604
rect 9692 34601 9720 34632
rect 9677 34595 9735 34601
rect 9677 34561 9689 34595
rect 9723 34561 9735 34595
rect 9677 34555 9735 34561
rect 9950 34552 9956 34604
rect 10008 34552 10014 34604
rect 10042 34552 10048 34604
rect 10100 34592 10106 34604
rect 10965 34595 11023 34601
rect 10965 34592 10977 34595
rect 10100 34564 10977 34592
rect 10100 34552 10106 34564
rect 10965 34561 10977 34564
rect 11011 34561 11023 34595
rect 10965 34555 11023 34561
rect 9769 34527 9827 34533
rect 9140 34496 9720 34524
rect 9692 34468 9720 34496
rect 9769 34493 9781 34527
rect 9815 34524 9827 34527
rect 10229 34527 10287 34533
rect 10229 34524 10241 34527
rect 9815 34496 10241 34524
rect 9815 34493 9827 34496
rect 9769 34487 9827 34493
rect 10229 34493 10241 34496
rect 10275 34493 10287 34527
rect 10229 34487 10287 34493
rect 10778 34484 10784 34536
rect 10836 34484 10842 34536
rect 11072 34524 11100 34632
rect 11149 34595 11207 34601
rect 11149 34561 11161 34595
rect 11195 34592 11207 34595
rect 11532 34592 11560 34700
rect 12360 34660 12388 34700
rect 12526 34688 12532 34740
rect 12584 34728 12590 34740
rect 12986 34728 12992 34740
rect 12584 34700 12992 34728
rect 12584 34688 12590 34700
rect 12986 34688 12992 34700
rect 13044 34688 13050 34740
rect 13354 34688 13360 34740
rect 13412 34688 13418 34740
rect 15010 34688 15016 34740
rect 15068 34688 15074 34740
rect 16022 34688 16028 34740
rect 16080 34688 16086 34740
rect 16114 34688 16120 34740
rect 16172 34688 16178 34740
rect 16206 34688 16212 34740
rect 16264 34688 16270 34740
rect 16298 34688 16304 34740
rect 16356 34688 16362 34740
rect 16393 34731 16451 34737
rect 16393 34697 16405 34731
rect 16439 34728 16451 34731
rect 16850 34728 16856 34740
rect 16439 34700 16856 34728
rect 16439 34697 16451 34700
rect 16393 34691 16451 34697
rect 16850 34688 16856 34700
rect 16908 34688 16914 34740
rect 17218 34688 17224 34740
rect 17276 34688 17282 34740
rect 17589 34731 17647 34737
rect 17589 34697 17601 34731
rect 17635 34728 17647 34731
rect 18874 34728 18880 34740
rect 17635 34700 18880 34728
rect 17635 34697 17647 34700
rect 17589 34691 17647 34697
rect 18874 34688 18880 34700
rect 18932 34728 18938 34740
rect 19058 34728 19064 34740
rect 18932 34700 19064 34728
rect 18932 34688 18938 34700
rect 19058 34688 19064 34700
rect 19116 34688 19122 34740
rect 19334 34688 19340 34740
rect 19392 34728 19398 34740
rect 20622 34728 20628 34740
rect 19392 34700 20628 34728
rect 19392 34688 19398 34700
rect 20622 34688 20628 34700
rect 20680 34688 20686 34740
rect 23385 34731 23443 34737
rect 23385 34697 23397 34731
rect 23431 34728 23443 34731
rect 24118 34728 24124 34740
rect 23431 34700 24124 34728
rect 23431 34697 23443 34700
rect 23385 34691 23443 34697
rect 24118 34688 24124 34700
rect 24176 34728 24182 34740
rect 24176 34700 25452 34728
rect 24176 34688 24182 34700
rect 13078 34660 13084 34672
rect 12360 34632 13084 34660
rect 13078 34620 13084 34632
rect 13136 34620 13142 34672
rect 13541 34663 13599 34669
rect 13541 34629 13553 34663
rect 13587 34660 13599 34663
rect 13587 34632 15700 34660
rect 13587 34629 13599 34632
rect 13541 34623 13599 34629
rect 11195 34564 11560 34592
rect 11195 34561 11207 34564
rect 11149 34555 11207 34561
rect 11606 34552 11612 34604
rect 11664 34552 11670 34604
rect 11698 34552 11704 34604
rect 11756 34592 11762 34604
rect 12244 34595 12302 34601
rect 11756 34590 12204 34592
rect 12244 34590 12256 34595
rect 11756 34564 12256 34590
rect 11756 34552 11762 34564
rect 12176 34562 12256 34564
rect 12244 34561 12256 34562
rect 12290 34561 12302 34595
rect 12244 34555 12302 34561
rect 12986 34552 12992 34604
rect 13044 34592 13050 34604
rect 13556 34592 13584 34623
rect 15672 34604 15700 34632
rect 13044 34564 13584 34592
rect 14369 34595 14427 34601
rect 13044 34552 13050 34564
rect 14369 34561 14381 34595
rect 14415 34561 14427 34595
rect 14369 34555 14427 34561
rect 11624 34524 11652 34552
rect 11977 34527 12035 34533
rect 11072 34496 11744 34524
rect 11716 34468 11744 34496
rect 11977 34493 11989 34527
rect 12023 34493 12035 34527
rect 14384 34524 14412 34555
rect 14734 34552 14740 34604
rect 14792 34592 14798 34604
rect 15197 34595 15255 34601
rect 15197 34592 15209 34595
rect 14792 34564 15209 34592
rect 14792 34552 14798 34564
rect 15197 34561 15209 34564
rect 15243 34561 15255 34595
rect 15197 34555 15255 34561
rect 15654 34552 15660 34604
rect 15712 34552 15718 34604
rect 14384 34496 15148 34524
rect 11977 34487 12035 34493
rect 9674 34416 9680 34468
rect 9732 34416 9738 34468
rect 11698 34416 11704 34468
rect 11756 34416 11762 34468
rect 8938 34348 8944 34400
rect 8996 34348 9002 34400
rect 9692 34388 9720 34416
rect 10502 34388 10508 34400
rect 9692 34360 10508 34388
rect 10502 34348 10508 34360
rect 10560 34388 10566 34400
rect 11790 34388 11796 34400
rect 10560 34360 11796 34388
rect 10560 34348 10566 34360
rect 11790 34348 11796 34360
rect 11848 34348 11854 34400
rect 11992 34388 12020 34487
rect 13817 34459 13875 34465
rect 13817 34425 13829 34459
rect 13863 34456 13875 34459
rect 14090 34456 14096 34468
rect 13863 34428 14096 34456
rect 13863 34425 13875 34428
rect 13817 34419 13875 34425
rect 14090 34416 14096 34428
rect 14148 34456 14154 34468
rect 14148 34428 14964 34456
rect 14148 34416 14154 34428
rect 14936 34400 14964 34428
rect 15120 34400 15148 34496
rect 15838 34484 15844 34536
rect 15896 34484 15902 34536
rect 16132 34524 16160 34688
rect 16224 34601 16252 34688
rect 16316 34660 16344 34688
rect 16316 34632 16528 34660
rect 16209 34595 16267 34601
rect 16209 34561 16221 34595
rect 16255 34561 16267 34595
rect 16209 34555 16267 34561
rect 16301 34595 16359 34601
rect 16301 34561 16313 34595
rect 16347 34561 16359 34595
rect 16301 34555 16359 34561
rect 16316 34524 16344 34555
rect 16390 34552 16396 34604
rect 16448 34552 16454 34604
rect 16500 34601 16528 34632
rect 18414 34620 18420 34672
rect 18472 34660 18478 34672
rect 18702 34663 18760 34669
rect 18702 34660 18714 34663
rect 18472 34632 18714 34660
rect 18472 34620 18478 34632
rect 18702 34629 18714 34632
rect 18748 34629 18760 34663
rect 18702 34623 18760 34629
rect 19150 34620 19156 34672
rect 19208 34660 19214 34672
rect 22373 34663 22431 34669
rect 19208 34632 22094 34660
rect 19208 34620 19214 34632
rect 16485 34595 16543 34601
rect 16485 34561 16497 34595
rect 16531 34561 16543 34595
rect 16485 34555 16543 34561
rect 18966 34552 18972 34604
rect 19024 34592 19030 34604
rect 19518 34601 19524 34604
rect 19245 34595 19303 34601
rect 19245 34592 19257 34595
rect 19024 34564 19257 34592
rect 19024 34552 19030 34564
rect 19245 34561 19257 34564
rect 19291 34561 19303 34595
rect 19245 34555 19303 34561
rect 19512 34555 19524 34601
rect 19518 34552 19524 34555
rect 19576 34552 19582 34604
rect 20622 34552 20628 34604
rect 20680 34592 20686 34604
rect 20717 34595 20775 34601
rect 20717 34592 20729 34595
rect 20680 34564 20729 34592
rect 20680 34552 20686 34564
rect 20717 34561 20729 34564
rect 20763 34561 20775 34595
rect 22066 34592 22094 34632
rect 22373 34629 22385 34663
rect 22419 34660 22431 34663
rect 22462 34660 22468 34672
rect 22419 34632 22468 34660
rect 22419 34629 22431 34632
rect 22373 34623 22431 34629
rect 22462 34620 22468 34632
rect 22520 34620 22526 34672
rect 22189 34595 22247 34601
rect 22189 34592 22201 34595
rect 22066 34564 22201 34592
rect 20717 34555 20775 34561
rect 22189 34561 22201 34564
rect 22235 34592 22247 34595
rect 22235 34564 22692 34592
rect 22235 34561 22247 34564
rect 22189 34555 22247 34561
rect 16132 34496 16344 34524
rect 16408 34524 16436 34552
rect 22664 34536 22692 34564
rect 24486 34552 24492 34604
rect 24544 34601 24550 34604
rect 25424 34601 25452 34700
rect 24544 34555 24556 34601
rect 25409 34595 25467 34601
rect 25409 34561 25421 34595
rect 25455 34561 25467 34595
rect 25409 34555 25467 34561
rect 24544 34552 24550 34555
rect 16761 34527 16819 34533
rect 16761 34524 16773 34527
rect 16408 34496 16773 34524
rect 16761 34493 16773 34496
rect 16807 34493 16819 34527
rect 16761 34487 16819 34493
rect 22005 34527 22063 34533
rect 22005 34493 22017 34527
rect 22051 34524 22063 34527
rect 22465 34527 22523 34533
rect 22465 34524 22477 34527
rect 22051 34496 22477 34524
rect 22051 34493 22063 34496
rect 22005 34487 22063 34493
rect 22465 34493 22477 34496
rect 22511 34493 22523 34527
rect 22465 34487 22523 34493
rect 22646 34484 22652 34536
rect 22704 34484 22710 34536
rect 23014 34484 23020 34536
rect 23072 34484 23078 34536
rect 24762 34484 24768 34536
rect 24820 34484 24826 34536
rect 17129 34459 17187 34465
rect 17129 34425 17141 34459
rect 17175 34456 17187 34459
rect 17310 34456 17316 34468
rect 17175 34428 17316 34456
rect 17175 34425 17187 34428
rect 17129 34419 17187 34425
rect 17310 34416 17316 34428
rect 17368 34416 17374 34468
rect 12158 34388 12164 34400
rect 11992 34360 12164 34388
rect 12158 34348 12164 34360
rect 12216 34348 12222 34400
rect 13354 34348 13360 34400
rect 13412 34388 13418 34400
rect 14277 34391 14335 34397
rect 14277 34388 14289 34391
rect 13412 34360 14289 34388
rect 13412 34348 13418 34360
rect 14277 34357 14289 34360
rect 14323 34357 14335 34391
rect 14277 34351 14335 34357
rect 14918 34348 14924 34400
rect 14976 34348 14982 34400
rect 15102 34348 15108 34400
rect 15160 34348 15166 34400
rect 15286 34348 15292 34400
rect 15344 34348 15350 34400
rect 15378 34348 15384 34400
rect 15436 34388 15442 34400
rect 20806 34388 20812 34400
rect 15436 34360 20812 34388
rect 15436 34348 15442 34360
rect 20806 34348 20812 34360
rect 20864 34348 20870 34400
rect 21358 34348 21364 34400
rect 21416 34348 21422 34400
rect 24854 34348 24860 34400
rect 24912 34348 24918 34400
rect 1104 34298 34868 34320
rect 1104 34246 5170 34298
rect 5222 34246 5234 34298
rect 5286 34246 5298 34298
rect 5350 34246 5362 34298
rect 5414 34246 5426 34298
rect 5478 34246 13611 34298
rect 13663 34246 13675 34298
rect 13727 34246 13739 34298
rect 13791 34246 13803 34298
rect 13855 34246 13867 34298
rect 13919 34246 22052 34298
rect 22104 34246 22116 34298
rect 22168 34246 22180 34298
rect 22232 34246 22244 34298
rect 22296 34246 22308 34298
rect 22360 34246 30493 34298
rect 30545 34246 30557 34298
rect 30609 34246 30621 34298
rect 30673 34246 30685 34298
rect 30737 34246 30749 34298
rect 30801 34246 34868 34298
rect 1104 34224 34868 34246
rect 8941 34187 8999 34193
rect 8941 34153 8953 34187
rect 8987 34184 8999 34187
rect 9214 34184 9220 34196
rect 8987 34156 9220 34184
rect 8987 34153 8999 34156
rect 8941 34147 8999 34153
rect 9214 34144 9220 34156
rect 9272 34144 9278 34196
rect 9677 34187 9735 34193
rect 9677 34153 9689 34187
rect 9723 34153 9735 34187
rect 9677 34147 9735 34153
rect 13725 34187 13783 34193
rect 13725 34153 13737 34187
rect 13771 34184 13783 34187
rect 14090 34184 14096 34196
rect 13771 34156 14096 34184
rect 13771 34153 13783 34156
rect 13725 34147 13783 34153
rect 8386 34076 8392 34128
rect 8444 34116 8450 34128
rect 9692 34116 9720 34147
rect 14090 34144 14096 34156
rect 14148 34144 14154 34196
rect 14918 34144 14924 34196
rect 14976 34184 14982 34196
rect 14976 34156 17540 34184
rect 14976 34144 14982 34156
rect 17512 34128 17540 34156
rect 17678 34144 17684 34196
rect 17736 34144 17742 34196
rect 18598 34144 18604 34196
rect 18656 34184 18662 34196
rect 18693 34187 18751 34193
rect 18693 34184 18705 34187
rect 18656 34156 18705 34184
rect 18656 34144 18662 34156
rect 18693 34153 18705 34156
rect 18739 34153 18751 34187
rect 20162 34184 20168 34196
rect 18693 34147 18751 34153
rect 18800 34156 20168 34184
rect 8444 34088 9720 34116
rect 12989 34119 13047 34125
rect 8444 34076 8450 34088
rect 12989 34085 13001 34119
rect 13035 34116 13047 34119
rect 13078 34116 13084 34128
rect 13035 34088 13084 34116
rect 13035 34085 13047 34088
rect 12989 34079 13047 34085
rect 8754 34008 8760 34060
rect 8812 34048 8818 34060
rect 9493 34051 9551 34057
rect 9493 34048 9505 34051
rect 8812 34020 9505 34048
rect 8812 34008 8818 34020
rect 9493 34017 9505 34020
rect 9539 34048 9551 34051
rect 9769 34051 9827 34057
rect 9769 34048 9781 34051
rect 9539 34020 9781 34048
rect 9539 34017 9551 34020
rect 9493 34011 9551 34017
rect 9769 34017 9781 34020
rect 9815 34017 9827 34051
rect 13004 34048 13032 34079
rect 13078 34076 13084 34088
rect 13136 34076 13142 34128
rect 13265 34119 13323 34125
rect 13265 34085 13277 34119
rect 13311 34116 13323 34119
rect 13541 34119 13599 34125
rect 13541 34116 13553 34119
rect 13311 34088 13553 34116
rect 13311 34085 13323 34088
rect 13265 34079 13323 34085
rect 13541 34085 13553 34088
rect 13587 34085 13599 34119
rect 13541 34079 13599 34085
rect 17494 34076 17500 34128
rect 17552 34116 17558 34128
rect 18800 34116 18828 34156
rect 20162 34144 20168 34156
rect 20220 34184 20226 34196
rect 23198 34184 23204 34196
rect 20220 34156 23204 34184
rect 20220 34144 20226 34156
rect 23198 34144 23204 34156
rect 23256 34144 23262 34196
rect 17552 34088 18828 34116
rect 17552 34076 17558 34088
rect 9769 34011 9827 34017
rect 12452 34020 13032 34048
rect 8478 33940 8484 33992
rect 8536 33940 8542 33992
rect 8573 33983 8631 33989
rect 8573 33949 8585 33983
rect 8619 33980 8631 33983
rect 8938 33980 8944 33992
rect 8619 33952 8944 33980
rect 8619 33949 8631 33952
rect 8573 33943 8631 33949
rect 8938 33940 8944 33952
rect 8996 33940 9002 33992
rect 9953 33983 10011 33989
rect 9953 33980 9965 33983
rect 9039 33952 9965 33980
rect 8846 33872 8852 33924
rect 8904 33912 8910 33924
rect 9039 33912 9067 33952
rect 9953 33949 9965 33952
rect 9999 33949 10011 33983
rect 9953 33943 10011 33949
rect 11974 33940 11980 33992
rect 12032 33980 12038 33992
rect 12452 33989 12480 34020
rect 13446 34008 13452 34060
rect 13504 34008 13510 34060
rect 14550 34048 14556 34060
rect 13740 34020 14556 34048
rect 12437 33983 12495 33989
rect 12437 33980 12449 33983
rect 12032 33952 12449 33980
rect 12032 33940 12038 33952
rect 12437 33949 12449 33952
rect 12483 33949 12495 33983
rect 12437 33943 12495 33949
rect 12526 33940 12532 33992
rect 12584 33940 12590 33992
rect 13173 33983 13231 33989
rect 13173 33949 13185 33983
rect 13219 33980 13231 33983
rect 13740 33980 13768 34020
rect 14550 34008 14556 34020
rect 14608 34008 14614 34060
rect 18690 34048 18696 34060
rect 17972 34020 18696 34048
rect 13219 33952 13768 33980
rect 13219 33949 13231 33952
rect 13173 33943 13231 33949
rect 13814 33940 13820 33992
rect 13872 33980 13878 33992
rect 13998 33980 14004 33992
rect 13872 33952 14004 33980
rect 13872 33940 13878 33952
rect 13998 33940 14004 33952
rect 14056 33980 14062 33992
rect 14737 33983 14795 33989
rect 14737 33980 14749 33983
rect 14056 33952 14749 33980
rect 14056 33940 14062 33952
rect 14737 33949 14749 33952
rect 14783 33949 14795 33983
rect 14737 33943 14795 33949
rect 15004 33983 15062 33989
rect 15004 33949 15016 33983
rect 15050 33980 15062 33983
rect 15286 33980 15292 33992
rect 15050 33952 15292 33980
rect 15050 33949 15062 33952
rect 15004 33943 15062 33949
rect 15286 33940 15292 33952
rect 15344 33940 15350 33992
rect 17972 33989 18000 34020
rect 18690 34008 18696 34020
rect 18748 34008 18754 34060
rect 16853 33983 16911 33989
rect 16853 33980 16865 33983
rect 16132 33952 16865 33980
rect 8904 33884 9067 33912
rect 9677 33915 9735 33921
rect 8904 33872 8910 33884
rect 9677 33881 9689 33915
rect 9723 33912 9735 33915
rect 9766 33912 9772 33924
rect 9723 33884 9772 33912
rect 9723 33881 9735 33884
rect 9677 33875 9735 33881
rect 9766 33872 9772 33884
rect 9824 33872 9830 33924
rect 10410 33872 10416 33924
rect 10468 33872 10474 33924
rect 11698 33872 11704 33924
rect 11756 33912 11762 33924
rect 12805 33915 12863 33921
rect 12805 33912 12817 33915
rect 11756 33884 12817 33912
rect 11756 33872 11762 33884
rect 12805 33881 12817 33884
rect 12851 33881 12863 33915
rect 12805 33875 12863 33881
rect 13449 33915 13507 33921
rect 13449 33881 13461 33915
rect 13495 33912 13507 33915
rect 13909 33915 13967 33921
rect 13495 33884 13860 33912
rect 13495 33881 13507 33884
rect 13449 33875 13507 33881
rect 8294 33804 8300 33856
rect 8352 33804 8358 33856
rect 8757 33847 8815 33853
rect 8757 33813 8769 33847
rect 8803 33844 8815 33847
rect 9214 33844 9220 33856
rect 8803 33816 9220 33844
rect 8803 33813 8815 33816
rect 8757 33807 8815 33813
rect 9214 33804 9220 33816
rect 9272 33804 9278 33856
rect 10137 33847 10195 33853
rect 10137 33813 10149 33847
rect 10183 33844 10195 33847
rect 10870 33844 10876 33856
rect 10183 33816 10876 33844
rect 10183 33813 10195 33816
rect 10137 33807 10195 33813
rect 10870 33804 10876 33816
rect 10928 33804 10934 33856
rect 11885 33847 11943 33853
rect 11885 33813 11897 33847
rect 11931 33844 11943 33847
rect 12158 33844 12164 33856
rect 11931 33816 12164 33844
rect 11931 33813 11943 33816
rect 11885 33807 11943 33813
rect 12158 33804 12164 33816
rect 12216 33804 12222 33856
rect 12250 33804 12256 33856
rect 12308 33804 12314 33856
rect 13722 33853 13728 33856
rect 13709 33847 13728 33853
rect 13709 33813 13721 33847
rect 13709 33807 13728 33813
rect 13722 33804 13728 33807
rect 13780 33804 13786 33856
rect 13832 33844 13860 33884
rect 13909 33881 13921 33915
rect 13955 33912 13967 33915
rect 14182 33912 14188 33924
rect 13955 33884 14188 33912
rect 13955 33881 13967 33884
rect 13909 33875 13967 33881
rect 14182 33872 14188 33884
rect 14240 33872 14246 33924
rect 14277 33915 14335 33921
rect 14277 33881 14289 33915
rect 14323 33912 14335 33915
rect 14366 33912 14372 33924
rect 14323 33884 14372 33912
rect 14323 33881 14335 33884
rect 14277 33875 14335 33881
rect 14366 33872 14372 33884
rect 14424 33872 14430 33924
rect 14461 33915 14519 33921
rect 14461 33881 14473 33915
rect 14507 33881 14519 33915
rect 14461 33875 14519 33881
rect 13998 33844 14004 33856
rect 13832 33816 14004 33844
rect 13998 33804 14004 33816
rect 14056 33804 14062 33856
rect 14476 33844 14504 33875
rect 15010 33844 15016 33856
rect 14476 33816 15016 33844
rect 15010 33804 15016 33816
rect 15068 33804 15074 33856
rect 15930 33804 15936 33856
rect 15988 33844 15994 33856
rect 16132 33853 16160 33952
rect 16853 33949 16865 33952
rect 16899 33949 16911 33983
rect 16853 33943 16911 33949
rect 17957 33983 18015 33989
rect 17957 33949 17969 33983
rect 18003 33949 18015 33983
rect 17957 33943 18015 33949
rect 18049 33983 18107 33989
rect 18049 33949 18061 33983
rect 18095 33949 18107 33983
rect 18049 33943 18107 33949
rect 18141 33983 18199 33989
rect 18141 33949 18153 33983
rect 18187 33980 18199 33983
rect 18230 33980 18236 33992
rect 18187 33952 18236 33980
rect 18187 33949 18199 33952
rect 18141 33943 18199 33949
rect 18064 33912 18092 33943
rect 18230 33940 18236 33952
rect 18288 33940 18294 33992
rect 18325 33983 18383 33989
rect 18325 33949 18337 33983
rect 18371 33980 18383 33983
rect 18800 33980 18828 34088
rect 24765 34051 24823 34057
rect 24765 34017 24777 34051
rect 24811 34048 24823 34051
rect 24854 34048 24860 34060
rect 24811 34020 24860 34048
rect 24811 34017 24823 34020
rect 24765 34011 24823 34017
rect 24854 34008 24860 34020
rect 24912 34008 24918 34060
rect 18371 33952 18828 33980
rect 18371 33949 18383 33952
rect 18325 33943 18383 33949
rect 19794 33940 19800 33992
rect 19852 33940 19858 33992
rect 20441 33983 20499 33989
rect 20441 33949 20453 33983
rect 20487 33980 20499 33983
rect 20717 33983 20775 33989
rect 20717 33980 20729 33983
rect 20487 33952 20729 33980
rect 20487 33949 20499 33952
rect 20441 33943 20499 33949
rect 20717 33949 20729 33952
rect 20763 33949 20775 33983
rect 20717 33943 20775 33949
rect 20806 33940 20812 33992
rect 20864 33980 20870 33992
rect 20901 33983 20959 33989
rect 20901 33980 20913 33983
rect 20864 33952 20913 33980
rect 20864 33940 20870 33952
rect 20901 33949 20913 33952
rect 20947 33980 20959 33983
rect 22373 33983 22431 33989
rect 20947 33952 22094 33980
rect 20947 33949 20959 33952
rect 20901 33943 20959 33949
rect 18064 33884 18552 33912
rect 18524 33856 18552 33884
rect 18782 33872 18788 33924
rect 18840 33912 18846 33924
rect 18840 33884 20760 33912
rect 18840 33872 18846 33884
rect 20732 33856 20760 33884
rect 16117 33847 16175 33853
rect 16117 33844 16129 33847
rect 15988 33816 16129 33844
rect 15988 33804 15994 33816
rect 16117 33813 16129 33816
rect 16163 33813 16175 33847
rect 16117 33807 16175 33813
rect 16669 33847 16727 33853
rect 16669 33813 16681 33847
rect 16715 33844 16727 33847
rect 16942 33844 16948 33856
rect 16715 33816 16948 33844
rect 16715 33813 16727 33816
rect 16669 33807 16727 33813
rect 16942 33804 16948 33816
rect 17000 33804 17006 33856
rect 18506 33804 18512 33856
rect 18564 33804 18570 33856
rect 19150 33804 19156 33856
rect 19208 33844 19214 33856
rect 19518 33844 19524 33856
rect 19208 33816 19524 33844
rect 19208 33804 19214 33816
rect 19518 33804 19524 33816
rect 19576 33804 19582 33856
rect 19702 33804 19708 33856
rect 19760 33844 19766 33856
rect 20533 33847 20591 33853
rect 20533 33844 20545 33847
rect 19760 33816 20545 33844
rect 19760 33804 19766 33816
rect 20533 33813 20545 33816
rect 20579 33813 20591 33847
rect 20533 33807 20591 33813
rect 20714 33804 20720 33856
rect 20772 33804 20778 33856
rect 20990 33804 20996 33856
rect 21048 33804 21054 33856
rect 22066 33844 22094 33952
rect 22373 33949 22385 33983
rect 22419 33980 22431 33983
rect 22465 33983 22523 33989
rect 22465 33980 22477 33983
rect 22419 33952 22477 33980
rect 22419 33949 22431 33952
rect 22373 33943 22431 33949
rect 22465 33949 22477 33952
rect 22511 33980 22523 33983
rect 24026 33980 24032 33992
rect 22511 33952 24032 33980
rect 22511 33949 22523 33952
rect 22465 33943 22523 33949
rect 24026 33940 24032 33952
rect 24084 33940 24090 33992
rect 24121 33983 24179 33989
rect 24121 33949 24133 33983
rect 24167 33980 24179 33983
rect 24397 33983 24455 33989
rect 24397 33980 24409 33983
rect 24167 33952 24409 33980
rect 24167 33949 24179 33952
rect 24121 33943 24179 33949
rect 24397 33949 24409 33952
rect 24443 33949 24455 33983
rect 24397 33943 24455 33949
rect 24581 33983 24639 33989
rect 24581 33949 24593 33983
rect 24627 33949 24639 33983
rect 24581 33943 24639 33949
rect 22128 33915 22186 33921
rect 22128 33881 22140 33915
rect 22174 33912 22186 33915
rect 22278 33912 22284 33924
rect 22174 33884 22284 33912
rect 22174 33881 22186 33884
rect 22128 33875 22186 33881
rect 22278 33872 22284 33884
rect 22336 33872 22342 33924
rect 22738 33921 22744 33924
rect 22732 33912 22744 33921
rect 22699 33884 22744 33912
rect 22732 33875 22744 33884
rect 22738 33872 22744 33875
rect 22796 33872 22802 33924
rect 23566 33872 23572 33924
rect 23624 33872 23630 33924
rect 24596 33912 24624 33943
rect 24320 33884 24624 33912
rect 23584 33844 23612 33872
rect 24320 33856 24348 33884
rect 22066 33816 23612 33844
rect 23842 33804 23848 33856
rect 23900 33804 23906 33856
rect 23934 33804 23940 33856
rect 23992 33804 23998 33856
rect 24302 33804 24308 33856
rect 24360 33804 24366 33856
rect 1104 33754 35027 33776
rect 1104 33702 9390 33754
rect 9442 33702 9454 33754
rect 9506 33702 9518 33754
rect 9570 33702 9582 33754
rect 9634 33702 9646 33754
rect 9698 33702 17831 33754
rect 17883 33702 17895 33754
rect 17947 33702 17959 33754
rect 18011 33702 18023 33754
rect 18075 33702 18087 33754
rect 18139 33702 26272 33754
rect 26324 33702 26336 33754
rect 26388 33702 26400 33754
rect 26452 33702 26464 33754
rect 26516 33702 26528 33754
rect 26580 33702 34713 33754
rect 34765 33702 34777 33754
rect 34829 33702 34841 33754
rect 34893 33702 34905 33754
rect 34957 33702 34969 33754
rect 35021 33702 35027 33754
rect 1104 33680 35027 33702
rect 8294 33600 8300 33652
rect 8352 33600 8358 33652
rect 8941 33643 8999 33649
rect 8941 33609 8953 33643
rect 8987 33640 8999 33643
rect 9306 33640 9312 33652
rect 8987 33612 9312 33640
rect 8987 33609 8999 33612
rect 8941 33603 8999 33609
rect 9306 33600 9312 33612
rect 9364 33640 9370 33652
rect 10042 33640 10048 33652
rect 9364 33612 10048 33640
rect 9364 33600 9370 33612
rect 10042 33600 10048 33612
rect 10100 33600 10106 33652
rect 11149 33643 11207 33649
rect 11149 33609 11161 33643
rect 11195 33609 11207 33643
rect 11149 33603 11207 33609
rect 7644 33575 7702 33581
rect 7644 33541 7656 33575
rect 7690 33572 7702 33575
rect 8312 33572 8340 33600
rect 7690 33544 8340 33572
rect 10812 33575 10870 33581
rect 7690 33541 7702 33544
rect 7644 33535 7702 33541
rect 10812 33541 10824 33575
rect 10858 33572 10870 33575
rect 11164 33572 11192 33603
rect 11238 33600 11244 33652
rect 11296 33600 11302 33652
rect 13722 33600 13728 33652
rect 13780 33640 13786 33652
rect 14274 33640 14280 33652
rect 13780 33612 14280 33640
rect 13780 33600 13786 33612
rect 14274 33600 14280 33612
rect 14332 33600 14338 33652
rect 15473 33643 15531 33649
rect 15473 33609 15485 33643
rect 15519 33640 15531 33643
rect 15838 33640 15844 33652
rect 15519 33612 15844 33640
rect 15519 33609 15531 33612
rect 15473 33603 15531 33609
rect 15838 33600 15844 33612
rect 15896 33600 15902 33652
rect 17773 33643 17831 33649
rect 15948 33612 17172 33640
rect 10858 33544 11192 33572
rect 10858 33541 10870 33544
rect 10812 33535 10870 33541
rect 11256 33504 11284 33600
rect 12158 33532 12164 33584
rect 12216 33572 12222 33584
rect 13814 33572 13820 33584
rect 12216 33544 13820 33572
rect 12216 33532 12222 33544
rect 11333 33507 11391 33513
rect 11333 33504 11345 33507
rect 11256 33476 11345 33504
rect 11333 33473 11345 33476
rect 11379 33473 11391 33507
rect 11333 33467 11391 33473
rect 12618 33464 12624 33516
rect 12676 33513 12682 33516
rect 12912 33513 12940 33544
rect 13814 33532 13820 33544
rect 13872 33532 13878 33584
rect 15948 33572 15976 33612
rect 17037 33575 17095 33581
rect 17037 33572 17049 33575
rect 14568 33544 15976 33572
rect 16040 33544 17049 33572
rect 12676 33504 12688 33513
rect 12897 33507 12955 33513
rect 12676 33476 12721 33504
rect 12676 33467 12688 33476
rect 12897 33473 12909 33507
rect 12943 33473 12955 33507
rect 12897 33467 12955 33473
rect 12676 33464 12682 33467
rect 13538 33464 13544 33516
rect 13596 33504 13602 33516
rect 14568 33513 14596 33544
rect 14553 33507 14611 33513
rect 14553 33504 14565 33507
rect 13596 33476 14565 33504
rect 13596 33464 13602 33476
rect 14553 33473 14565 33476
rect 14599 33473 14611 33507
rect 14553 33467 14611 33473
rect 14734 33464 14740 33516
rect 14792 33464 14798 33516
rect 14829 33507 14887 33513
rect 14829 33473 14841 33507
rect 14875 33504 14887 33507
rect 14918 33504 14924 33516
rect 14875 33476 14924 33504
rect 14875 33473 14887 33476
rect 14829 33467 14887 33473
rect 14918 33464 14924 33476
rect 14976 33464 14982 33516
rect 15120 33513 15148 33544
rect 15013 33507 15071 33513
rect 15013 33473 15025 33507
rect 15059 33473 15071 33507
rect 15013 33467 15071 33473
rect 15105 33507 15163 33513
rect 15105 33473 15117 33507
rect 15151 33473 15163 33507
rect 15105 33467 15163 33473
rect 15197 33507 15255 33513
rect 15197 33473 15209 33507
rect 15243 33504 15255 33507
rect 15470 33504 15476 33516
rect 15243 33476 15476 33504
rect 15243 33473 15255 33476
rect 15197 33467 15255 33473
rect 7374 33396 7380 33448
rect 7432 33396 7438 33448
rect 9585 33439 9643 33445
rect 9585 33405 9597 33439
rect 9631 33405 9643 33439
rect 9585 33399 9643 33405
rect 11057 33439 11115 33445
rect 11057 33405 11069 33439
rect 11103 33436 11115 33439
rect 11103 33408 11948 33436
rect 11103 33405 11115 33408
rect 11057 33399 11115 33405
rect 9600 33368 9628 33399
rect 9677 33371 9735 33377
rect 9677 33368 9689 33371
rect 9600 33340 9689 33368
rect 9677 33337 9689 33340
rect 9723 33337 9735 33371
rect 9677 33331 9735 33337
rect 8754 33260 8760 33312
rect 8812 33260 8818 33312
rect 11514 33260 11520 33312
rect 11572 33260 11578 33312
rect 11920 33300 11948 33408
rect 13354 33396 13360 33448
rect 13412 33436 13418 33448
rect 13633 33439 13691 33445
rect 13633 33436 13645 33439
rect 13412 33408 13645 33436
rect 13412 33396 13418 33408
rect 13633 33405 13645 33408
rect 13679 33405 13691 33439
rect 13633 33399 13691 33405
rect 14458 33396 14464 33448
rect 14516 33396 14522 33448
rect 14645 33439 14703 33445
rect 14645 33405 14657 33439
rect 14691 33436 14703 33439
rect 15028 33436 15056 33467
rect 15470 33464 15476 33476
rect 15528 33464 15534 33516
rect 15565 33507 15623 33513
rect 15565 33473 15577 33507
rect 15611 33504 15623 33507
rect 15933 33507 15991 33513
rect 15611 33476 15792 33504
rect 15611 33473 15623 33476
rect 15565 33467 15623 33473
rect 15764 33448 15792 33476
rect 15933 33473 15945 33507
rect 15979 33504 15991 33507
rect 16040 33504 16068 33544
rect 17037 33541 17049 33544
rect 17083 33541 17095 33575
rect 17144 33572 17172 33612
rect 17773 33609 17785 33643
rect 17819 33640 17831 33643
rect 18230 33640 18236 33652
rect 17819 33612 18236 33640
rect 17819 33609 17831 33612
rect 17773 33603 17831 33609
rect 18230 33600 18236 33612
rect 18288 33600 18294 33652
rect 19702 33640 19708 33652
rect 18984 33612 19708 33640
rect 17144 33544 17816 33572
rect 17037 33535 17095 33541
rect 15979 33476 16068 33504
rect 15979 33473 15991 33476
rect 15933 33467 15991 33473
rect 14691 33408 15056 33436
rect 14691 33405 14703 33408
rect 14645 33399 14703 33405
rect 15746 33396 15752 33448
rect 15804 33396 15810 33448
rect 15841 33439 15899 33445
rect 15841 33405 15853 33439
rect 15887 33436 15899 33439
rect 15948 33436 15976 33467
rect 16114 33464 16120 33516
rect 16172 33464 16178 33516
rect 16574 33464 16580 33516
rect 16632 33504 16638 33516
rect 16669 33507 16727 33513
rect 16669 33504 16681 33507
rect 16632 33476 16681 33504
rect 16632 33464 16638 33476
rect 16669 33473 16681 33476
rect 16715 33473 16727 33507
rect 16669 33467 16727 33473
rect 16850 33464 16856 33516
rect 16908 33464 16914 33516
rect 16942 33464 16948 33516
rect 17000 33464 17006 33516
rect 17126 33464 17132 33516
rect 17184 33464 17190 33516
rect 15887 33408 15976 33436
rect 15887 33405 15899 33408
rect 15841 33399 15899 33405
rect 16206 33396 16212 33448
rect 16264 33436 16270 33448
rect 16960 33436 16988 33464
rect 17788 33445 17816 33544
rect 18046 33464 18052 33516
rect 18104 33464 18110 33516
rect 18984 33513 19012 33612
rect 19702 33600 19708 33612
rect 19760 33600 19766 33652
rect 19794 33600 19800 33652
rect 19852 33600 19858 33652
rect 22649 33643 22707 33649
rect 22649 33609 22661 33643
rect 22695 33640 22707 33643
rect 23014 33640 23020 33652
rect 22695 33612 23020 33640
rect 22695 33609 22707 33612
rect 22649 33603 22707 33609
rect 23014 33600 23020 33612
rect 23072 33600 23078 33652
rect 23934 33600 23940 33652
rect 23992 33600 23998 33652
rect 24486 33600 24492 33652
rect 24544 33640 24550 33652
rect 24581 33643 24639 33649
rect 24581 33640 24593 33643
rect 24544 33612 24593 33640
rect 24544 33600 24550 33612
rect 24581 33609 24593 33612
rect 24627 33609 24639 33643
rect 24581 33603 24639 33609
rect 24762 33600 24768 33652
rect 24820 33600 24826 33652
rect 19150 33532 19156 33584
rect 19208 33532 19214 33584
rect 19543 33575 19601 33581
rect 19543 33541 19555 33575
rect 19589 33572 19601 33575
rect 19812 33572 19840 33600
rect 20349 33575 20407 33581
rect 20349 33572 20361 33575
rect 19589 33544 19840 33572
rect 19904 33544 20361 33572
rect 19589 33541 19601 33544
rect 19543 33535 19601 33541
rect 18969 33507 19027 33513
rect 18969 33473 18981 33507
rect 19015 33473 19027 33507
rect 18969 33467 19027 33473
rect 17773 33439 17831 33445
rect 16264 33408 17356 33436
rect 16264 33396 16270 33408
rect 17328 33380 17356 33408
rect 17773 33405 17785 33439
rect 17819 33436 17831 33439
rect 17819 33408 18552 33436
rect 17819 33405 17831 33408
rect 17773 33399 17831 33405
rect 18524 33380 18552 33408
rect 15654 33328 15660 33380
rect 15712 33368 15718 33380
rect 16025 33371 16083 33377
rect 16025 33368 16037 33371
rect 15712 33340 16037 33368
rect 15712 33328 15718 33340
rect 16025 33337 16037 33340
rect 16071 33337 16083 33371
rect 16025 33331 16083 33337
rect 17310 33328 17316 33380
rect 17368 33328 17374 33380
rect 18506 33328 18512 33380
rect 18564 33328 18570 33380
rect 19168 33377 19196 33532
rect 19245 33507 19303 33513
rect 19245 33473 19257 33507
rect 19291 33473 19303 33507
rect 19904 33504 19932 33544
rect 20349 33541 20361 33544
rect 20395 33541 20407 33575
rect 21358 33572 21364 33584
rect 20349 33535 20407 33541
rect 20916 33544 21364 33572
rect 19245 33467 19303 33473
rect 19444 33476 19932 33504
rect 19153 33371 19211 33377
rect 19153 33337 19165 33371
rect 19199 33337 19211 33371
rect 19153 33331 19211 33337
rect 12710 33300 12716 33312
rect 11920 33272 12716 33300
rect 12710 33260 12716 33272
rect 12768 33260 12774 33312
rect 13078 33260 13084 33312
rect 13136 33260 13142 33312
rect 13817 33303 13875 33309
rect 13817 33269 13829 33303
rect 13863 33300 13875 33303
rect 14366 33300 14372 33312
rect 13863 33272 14372 33300
rect 13863 33269 13875 33272
rect 13817 33263 13875 33269
rect 14366 33260 14372 33272
rect 14424 33300 14430 33312
rect 14918 33300 14924 33312
rect 14424 33272 14924 33300
rect 14424 33260 14430 33272
rect 14918 33260 14924 33272
rect 14976 33260 14982 33312
rect 15562 33260 15568 33312
rect 15620 33300 15626 33312
rect 15749 33303 15807 33309
rect 15749 33300 15761 33303
rect 15620 33272 15761 33300
rect 15620 33260 15626 33272
rect 15749 33269 15761 33272
rect 15795 33300 15807 33303
rect 16298 33300 16304 33312
rect 15795 33272 16304 33300
rect 15795 33269 15807 33272
rect 15749 33263 15807 33269
rect 16298 33260 16304 33272
rect 16356 33260 16362 33312
rect 16853 33303 16911 33309
rect 16853 33269 16865 33303
rect 16899 33300 16911 33303
rect 17957 33303 18015 33309
rect 17957 33300 17969 33303
rect 16899 33272 17969 33300
rect 16899 33269 16911 33272
rect 16853 33263 16911 33269
rect 17957 33269 17969 33272
rect 18003 33300 18015 33303
rect 18690 33300 18696 33312
rect 18003 33272 18696 33300
rect 18003 33269 18015 33272
rect 17957 33263 18015 33269
rect 18690 33260 18696 33272
rect 18748 33260 18754 33312
rect 19260 33300 19288 33467
rect 19444 33445 19472 33476
rect 20162 33464 20168 33516
rect 20220 33504 20226 33516
rect 20916 33513 20944 33544
rect 21358 33532 21364 33544
rect 21416 33532 21422 33584
rect 23784 33575 23842 33581
rect 23784 33541 23796 33575
rect 23830 33572 23842 33575
rect 23952 33572 23980 33600
rect 24780 33572 24808 33600
rect 23830 33544 23980 33572
rect 24044 33544 24808 33572
rect 23830 33541 23842 33544
rect 23784 33535 23842 33541
rect 24044 33516 24072 33544
rect 20441 33507 20499 33513
rect 20441 33504 20453 33507
rect 20220 33476 20453 33504
rect 20220 33464 20226 33476
rect 20441 33473 20453 33476
rect 20487 33473 20499 33507
rect 20441 33467 20499 33473
rect 20625 33507 20683 33513
rect 20625 33473 20637 33507
rect 20671 33473 20683 33507
rect 20625 33467 20683 33473
rect 20901 33507 20959 33513
rect 20901 33473 20913 33507
rect 20947 33473 20959 33507
rect 20901 33467 20959 33473
rect 19429 33439 19487 33445
rect 19429 33405 19441 33439
rect 19475 33405 19487 33439
rect 19705 33439 19763 33445
rect 19705 33436 19717 33439
rect 19429 33399 19487 33405
rect 19536 33408 19717 33436
rect 19536 33380 19564 33408
rect 19705 33405 19717 33408
rect 19751 33405 19763 33439
rect 19705 33399 19763 33405
rect 20073 33439 20131 33445
rect 20073 33405 20085 33439
rect 20119 33436 20131 33439
rect 20640 33436 20668 33467
rect 20990 33464 20996 33516
rect 21048 33504 21054 33516
rect 21821 33507 21879 33513
rect 21821 33504 21833 33507
rect 21048 33476 21833 33504
rect 21048 33464 21054 33476
rect 21821 33473 21833 33476
rect 21867 33473 21879 33507
rect 21821 33467 21879 33473
rect 24026 33464 24032 33516
rect 24084 33464 24090 33516
rect 24210 33464 24216 33516
rect 24268 33464 24274 33516
rect 24302 33464 24308 33516
rect 24360 33464 24366 33516
rect 24489 33507 24547 33513
rect 24489 33473 24501 33507
rect 24535 33504 24547 33507
rect 24765 33507 24823 33513
rect 24765 33504 24777 33507
rect 24535 33476 24777 33504
rect 24535 33473 24547 33476
rect 24489 33467 24547 33473
rect 24765 33473 24777 33476
rect 24811 33473 24823 33507
rect 24765 33467 24823 33473
rect 20119 33408 21128 33436
rect 20119 33405 20131 33408
rect 20073 33399 20131 33405
rect 19337 33371 19395 33377
rect 19337 33337 19349 33371
rect 19383 33368 19395 33371
rect 19518 33368 19524 33380
rect 19383 33340 19524 33368
rect 19383 33337 19395 33340
rect 19337 33331 19395 33337
rect 19518 33328 19524 33340
rect 19576 33328 19582 33380
rect 19610 33328 19616 33380
rect 19668 33328 19674 33380
rect 20809 33371 20867 33377
rect 20809 33368 20821 33371
rect 19720 33340 20821 33368
rect 19720 33300 19748 33340
rect 20809 33337 20821 33340
rect 20855 33337 20867 33371
rect 20809 33331 20867 33337
rect 21100 33312 21128 33408
rect 22465 33371 22523 33377
rect 22465 33337 22477 33371
rect 22511 33368 22523 33371
rect 22511 33340 22876 33368
rect 22511 33337 22523 33340
rect 22465 33331 22523 33337
rect 22848 33312 22876 33340
rect 19260 33272 19748 33300
rect 19794 33260 19800 33312
rect 19852 33300 19858 33312
rect 20162 33300 20168 33312
rect 19852 33272 20168 33300
rect 19852 33260 19858 33272
rect 20162 33260 20168 33272
rect 20220 33260 20226 33312
rect 20438 33260 20444 33312
rect 20496 33260 20502 33312
rect 21082 33260 21088 33312
rect 21140 33260 21146 33312
rect 22830 33260 22836 33312
rect 22888 33260 22894 33312
rect 23290 33260 23296 33312
rect 23348 33300 23354 33312
rect 24320 33300 24348 33464
rect 23348 33272 24348 33300
rect 23348 33260 23354 33272
rect 1104 33210 34868 33232
rect 1104 33158 5170 33210
rect 5222 33158 5234 33210
rect 5286 33158 5298 33210
rect 5350 33158 5362 33210
rect 5414 33158 5426 33210
rect 5478 33158 13611 33210
rect 13663 33158 13675 33210
rect 13727 33158 13739 33210
rect 13791 33158 13803 33210
rect 13855 33158 13867 33210
rect 13919 33158 22052 33210
rect 22104 33158 22116 33210
rect 22168 33158 22180 33210
rect 22232 33158 22244 33210
rect 22296 33158 22308 33210
rect 22360 33158 30493 33210
rect 30545 33158 30557 33210
rect 30609 33158 30621 33210
rect 30673 33158 30685 33210
rect 30737 33158 30749 33210
rect 30801 33158 34868 33210
rect 1104 33136 34868 33158
rect 8021 33099 8079 33105
rect 8021 33065 8033 33099
rect 8067 33096 8079 33099
rect 8478 33096 8484 33108
rect 8067 33068 8484 33096
rect 8067 33065 8079 33068
rect 8021 33059 8079 33065
rect 8478 33056 8484 33068
rect 8536 33056 8542 33108
rect 10042 33056 10048 33108
rect 10100 33096 10106 33108
rect 10321 33099 10379 33105
rect 10321 33096 10333 33099
rect 10100 33068 10333 33096
rect 10100 33056 10106 33068
rect 10321 33065 10333 33068
rect 10367 33096 10379 33099
rect 10778 33096 10784 33108
rect 10367 33068 10784 33096
rect 10367 33065 10379 33068
rect 10321 33059 10379 33065
rect 10778 33056 10784 33068
rect 10836 33056 10842 33108
rect 12253 33099 12311 33105
rect 12253 33065 12265 33099
rect 12299 33096 12311 33099
rect 12526 33096 12532 33108
rect 12299 33068 12532 33096
rect 12299 33065 12311 33068
rect 12253 33059 12311 33065
rect 12526 33056 12532 33068
rect 12584 33056 12590 33108
rect 14090 33056 14096 33108
rect 14148 33056 14154 33108
rect 14734 33056 14740 33108
rect 14792 33096 14798 33108
rect 15013 33099 15071 33105
rect 15013 33096 15025 33099
rect 14792 33068 15025 33096
rect 14792 33056 14798 33068
rect 15013 33065 15025 33068
rect 15059 33065 15071 33099
rect 15013 33059 15071 33065
rect 16114 33056 16120 33108
rect 16172 33056 16178 33108
rect 16850 33056 16856 33108
rect 16908 33096 16914 33108
rect 17037 33099 17095 33105
rect 17037 33096 17049 33099
rect 16908 33068 17049 33096
rect 16908 33056 16914 33068
rect 17037 33065 17049 33068
rect 17083 33096 17095 33099
rect 17083 33068 17908 33096
rect 17083 33065 17095 33068
rect 17037 33059 17095 33065
rect 7926 32988 7932 33040
rect 7984 33028 7990 33040
rect 8754 33028 8760 33040
rect 7984 33000 8760 33028
rect 7984 32988 7990 33000
rect 8754 32988 8760 33000
rect 8812 32988 8818 33040
rect 13909 33031 13967 33037
rect 13909 32997 13921 33031
rect 13955 32997 13967 33031
rect 14108 33028 14136 33056
rect 14108 33000 14780 33028
rect 13909 32991 13967 32997
rect 7653 32963 7711 32969
rect 7653 32929 7665 32963
rect 7699 32960 7711 32963
rect 8113 32963 8171 32969
rect 8113 32960 8125 32963
rect 7699 32932 8125 32960
rect 7699 32929 7711 32932
rect 7653 32923 7711 32929
rect 8113 32929 8125 32932
rect 8159 32929 8171 32963
rect 12250 32960 12256 32972
rect 8113 32923 8171 32929
rect 11348 32932 12256 32960
rect 7837 32895 7895 32901
rect 7837 32861 7849 32895
rect 7883 32892 7895 32895
rect 8570 32892 8576 32904
rect 7883 32864 8576 32892
rect 7883 32861 7895 32864
rect 7837 32855 7895 32861
rect 8312 32836 8340 32864
rect 8570 32852 8576 32864
rect 8628 32852 8634 32904
rect 8757 32895 8815 32901
rect 8757 32861 8769 32895
rect 8803 32861 8815 32895
rect 8757 32855 8815 32861
rect 8941 32895 8999 32901
rect 8941 32861 8953 32895
rect 8987 32892 8999 32895
rect 9030 32892 9036 32904
rect 8987 32864 9036 32892
rect 8987 32861 8999 32864
rect 8941 32855 8999 32861
rect 8294 32784 8300 32836
rect 8352 32784 8358 32836
rect 7834 32716 7840 32768
rect 7892 32756 7898 32768
rect 8772 32756 8800 32855
rect 9030 32852 9036 32864
rect 9088 32852 9094 32904
rect 9214 32901 9220 32904
rect 9208 32892 9220 32901
rect 9175 32864 9220 32892
rect 9208 32855 9220 32864
rect 9214 32852 9220 32855
rect 9272 32852 9278 32904
rect 11348 32901 11376 32932
rect 12250 32920 12256 32932
rect 12308 32920 12314 32972
rect 13924 32960 13952 32991
rect 14752 32972 14780 33000
rect 15470 32988 15476 33040
rect 15528 33028 15534 33040
rect 17402 33028 17408 33040
rect 15528 33000 15976 33028
rect 15528 32988 15534 33000
rect 14458 32960 14464 32972
rect 13924 32932 14464 32960
rect 14458 32920 14464 32932
rect 14516 32920 14522 32972
rect 14734 32920 14740 32972
rect 14792 32920 14798 32972
rect 15381 32963 15439 32969
rect 15381 32929 15393 32963
rect 15427 32960 15439 32963
rect 15654 32960 15660 32972
rect 15427 32932 15660 32960
rect 15427 32929 15439 32932
rect 15381 32923 15439 32929
rect 15654 32920 15660 32932
rect 15712 32920 15718 32972
rect 15746 32920 15752 32972
rect 15804 32920 15810 32972
rect 10505 32895 10563 32901
rect 10505 32861 10517 32895
rect 10551 32861 10563 32895
rect 10505 32855 10563 32861
rect 11333 32895 11391 32901
rect 11333 32861 11345 32895
rect 11379 32861 11391 32895
rect 11333 32855 11391 32861
rect 9122 32784 9128 32836
rect 9180 32824 9186 32836
rect 10520 32824 10548 32855
rect 11514 32852 11520 32904
rect 11572 32892 11578 32904
rect 11609 32895 11667 32901
rect 11609 32892 11621 32895
rect 11572 32864 11621 32892
rect 11572 32852 11578 32864
rect 11609 32861 11621 32864
rect 11655 32861 11667 32895
rect 11609 32855 11667 32861
rect 12529 32895 12587 32901
rect 12529 32861 12541 32895
rect 12575 32892 12587 32895
rect 12796 32895 12854 32901
rect 12575 32864 12756 32892
rect 12575 32861 12587 32864
rect 12529 32855 12587 32861
rect 9180 32796 10548 32824
rect 9180 32784 9186 32796
rect 12728 32768 12756 32864
rect 12796 32861 12808 32895
rect 12842 32892 12854 32895
rect 13078 32892 13084 32904
rect 12842 32864 13084 32892
rect 12842 32861 12854 32864
rect 12796 32855 12854 32861
rect 13078 32852 13084 32864
rect 13136 32852 13142 32904
rect 14093 32895 14151 32901
rect 14093 32861 14105 32895
rect 14139 32892 14151 32895
rect 14274 32892 14280 32904
rect 14139 32864 14280 32892
rect 14139 32861 14151 32864
rect 14093 32855 14151 32861
rect 14274 32852 14280 32864
rect 14332 32852 14338 32904
rect 14642 32852 14648 32904
rect 14700 32852 14706 32904
rect 15289 32895 15347 32901
rect 15289 32861 15301 32895
rect 15335 32892 15347 32895
rect 15764 32892 15792 32920
rect 15948 32901 15976 33000
rect 16408 33000 17408 33028
rect 15335 32864 15792 32892
rect 15933 32895 15991 32901
rect 15335 32861 15347 32864
rect 15289 32855 15347 32861
rect 15933 32861 15945 32895
rect 15979 32892 15991 32895
rect 16206 32892 16212 32904
rect 15979 32864 16212 32892
rect 15979 32861 15991 32864
rect 15933 32855 15991 32861
rect 14292 32824 14320 32852
rect 14826 32824 14832 32836
rect 14292 32796 14832 32824
rect 14826 32784 14832 32796
rect 14884 32784 14890 32836
rect 9766 32756 9772 32768
rect 7892 32728 9772 32756
rect 7892 32716 7898 32728
rect 9766 32716 9772 32728
rect 9824 32756 9830 32768
rect 10318 32756 10324 32768
rect 9824 32728 10324 32756
rect 9824 32716 9830 32728
rect 10318 32716 10324 32728
rect 10376 32716 10382 32768
rect 11149 32759 11207 32765
rect 11149 32725 11161 32759
rect 11195 32756 11207 32759
rect 11330 32756 11336 32768
rect 11195 32728 11336 32756
rect 11195 32725 11207 32728
rect 11149 32719 11207 32725
rect 11330 32716 11336 32728
rect 11388 32716 11394 32768
rect 11514 32716 11520 32768
rect 11572 32716 11578 32768
rect 12710 32716 12716 32768
rect 12768 32716 12774 32768
rect 14645 32759 14703 32765
rect 14645 32725 14657 32759
rect 14691 32756 14703 32759
rect 15304 32756 15332 32855
rect 16206 32852 16212 32864
rect 16264 32852 16270 32904
rect 16301 32895 16359 32901
rect 16301 32861 16313 32895
rect 16347 32892 16359 32895
rect 16408 32892 16436 33000
rect 17402 32988 17408 33000
rect 17460 32988 17466 33040
rect 17221 32963 17279 32969
rect 17221 32929 17233 32963
rect 17267 32929 17279 32963
rect 17221 32923 17279 32929
rect 16347 32864 16436 32892
rect 16347 32861 16359 32864
rect 16301 32855 16359 32861
rect 15470 32784 15476 32836
rect 15528 32824 15534 32836
rect 15749 32827 15807 32833
rect 15749 32824 15761 32827
rect 15528 32796 15761 32824
rect 15528 32784 15534 32796
rect 15749 32793 15761 32796
rect 15795 32824 15807 32827
rect 16316 32824 16344 32855
rect 17126 32824 17132 32836
rect 15795 32796 16344 32824
rect 16408 32796 17132 32824
rect 15795 32793 15807 32796
rect 15749 32787 15807 32793
rect 14691 32728 15332 32756
rect 14691 32725 14703 32728
rect 14645 32719 14703 32725
rect 16206 32716 16212 32768
rect 16264 32756 16270 32768
rect 16408 32765 16436 32796
rect 17126 32784 17132 32796
rect 17184 32824 17190 32836
rect 17236 32824 17264 32923
rect 17313 32895 17371 32901
rect 17313 32861 17325 32895
rect 17359 32861 17371 32895
rect 17313 32855 17371 32861
rect 17681 32895 17739 32901
rect 17681 32861 17693 32895
rect 17727 32861 17739 32895
rect 17681 32855 17739 32861
rect 17184 32796 17264 32824
rect 17184 32784 17190 32796
rect 16393 32759 16451 32765
rect 16393 32756 16405 32759
rect 16264 32728 16405 32756
rect 16264 32716 16270 32728
rect 16393 32725 16405 32728
rect 16439 32725 16451 32759
rect 17328 32756 17356 32855
rect 17586 32784 17592 32836
rect 17644 32824 17650 32836
rect 17696 32824 17724 32855
rect 17770 32852 17776 32904
rect 17828 32852 17834 32904
rect 17880 32901 17908 33068
rect 18046 33056 18052 33108
rect 18104 33096 18110 33108
rect 19245 33099 19303 33105
rect 19245 33096 19257 33099
rect 18104 33068 19257 33096
rect 18104 33056 18110 33068
rect 19245 33065 19257 33068
rect 19291 33065 19303 33099
rect 19245 33059 19303 33065
rect 19610 33056 19616 33108
rect 19668 33096 19674 33108
rect 20438 33096 20444 33108
rect 19668 33068 20444 33096
rect 19668 33056 19674 33068
rect 20438 33056 20444 33068
rect 20496 33096 20502 33108
rect 20533 33099 20591 33105
rect 20533 33096 20545 33099
rect 20496 33068 20545 33096
rect 20496 33056 20502 33068
rect 20533 33065 20545 33068
rect 20579 33065 20591 33099
rect 20533 33059 20591 33065
rect 21082 33056 21088 33108
rect 21140 33056 21146 33108
rect 22281 33099 22339 33105
rect 22281 33065 22293 33099
rect 22327 33096 22339 33099
rect 22370 33096 22376 33108
rect 22327 33068 22376 33096
rect 22327 33065 22339 33068
rect 22281 33059 22339 33065
rect 22370 33056 22376 33068
rect 22428 33056 22434 33108
rect 22554 33056 22560 33108
rect 22612 33056 22618 33108
rect 24210 33056 24216 33108
rect 24268 33096 24274 33108
rect 24673 33099 24731 33105
rect 24673 33096 24685 33099
rect 24268 33068 24685 33096
rect 24268 33056 24274 33068
rect 24673 33065 24685 33068
rect 24719 33065 24731 33099
rect 24673 33059 24731 33065
rect 18141 33031 18199 33037
rect 18141 32997 18153 33031
rect 18187 33028 18199 33031
rect 19794 33028 19800 33040
rect 18187 33000 19800 33028
rect 18187 32997 18199 33000
rect 18141 32991 18199 32997
rect 19794 32988 19800 33000
rect 19852 32988 19858 33040
rect 20070 32988 20076 33040
rect 20128 33028 20134 33040
rect 22189 33031 22247 33037
rect 20128 33000 20852 33028
rect 20128 32988 20134 33000
rect 18877 32963 18935 32969
rect 18877 32929 18889 32963
rect 18923 32960 18935 32963
rect 20714 32960 20720 32972
rect 18923 32932 20720 32960
rect 18923 32929 18935 32932
rect 18877 32923 18935 32929
rect 20714 32920 20720 32932
rect 20772 32920 20778 32972
rect 17865 32895 17923 32901
rect 17865 32861 17877 32895
rect 17911 32861 17923 32895
rect 17865 32855 17923 32861
rect 17957 32895 18015 32901
rect 17957 32861 17969 32895
rect 18003 32892 18015 32895
rect 18138 32892 18144 32904
rect 18003 32864 18144 32892
rect 18003 32861 18015 32864
rect 17957 32855 18015 32861
rect 17644 32796 17724 32824
rect 17880 32824 17908 32855
rect 18138 32852 18144 32864
rect 18196 32852 18202 32904
rect 18325 32895 18383 32901
rect 18325 32861 18337 32895
rect 18371 32892 18383 32895
rect 18598 32892 18604 32904
rect 18371 32864 18604 32892
rect 18371 32861 18383 32864
rect 18325 32855 18383 32861
rect 18598 32852 18604 32864
rect 18656 32852 18662 32904
rect 19429 32895 19487 32901
rect 19429 32861 19441 32895
rect 19475 32861 19487 32895
rect 19429 32855 19487 32861
rect 19435 32824 19463 32855
rect 19518 32852 19524 32904
rect 19576 32852 19582 32904
rect 19705 32895 19763 32901
rect 19705 32861 19717 32895
rect 19751 32861 19763 32895
rect 19705 32855 19763 32861
rect 19889 32895 19947 32901
rect 19889 32861 19901 32895
rect 19935 32892 19947 32895
rect 20070 32892 20076 32904
rect 19935 32864 20076 32892
rect 19935 32861 19947 32864
rect 19889 32855 19947 32861
rect 19720 32824 19748 32855
rect 20070 32852 20076 32864
rect 20128 32852 20134 32904
rect 20346 32852 20352 32904
rect 20404 32852 20410 32904
rect 20625 32895 20683 32901
rect 20625 32861 20637 32895
rect 20671 32861 20683 32895
rect 20824 32892 20852 33000
rect 22189 32997 22201 33031
rect 22235 33028 22247 33031
rect 22572 33028 22600 33056
rect 22235 33000 22600 33028
rect 22235 32997 22247 33000
rect 22189 32991 22247 32997
rect 21821 32963 21879 32969
rect 21821 32929 21833 32963
rect 21867 32960 21879 32963
rect 22830 32960 22836 32972
rect 21867 32932 22836 32960
rect 21867 32929 21879 32932
rect 21821 32923 21879 32929
rect 22830 32920 22836 32932
rect 22888 32920 22894 32972
rect 23290 32960 23296 32972
rect 23032 32932 23296 32960
rect 21177 32895 21235 32901
rect 21177 32892 21189 32895
rect 20824 32864 21189 32892
rect 20625 32855 20683 32861
rect 21177 32861 21189 32864
rect 21223 32861 21235 32895
rect 21177 32855 21235 32861
rect 20640 32824 20668 32855
rect 21358 32852 21364 32904
rect 21416 32852 21422 32904
rect 22005 32895 22063 32901
rect 22005 32861 22017 32895
rect 22051 32861 22063 32895
rect 22005 32855 22063 32861
rect 20717 32827 20775 32833
rect 20717 32824 20729 32827
rect 17880 32796 19463 32824
rect 19628 32796 19748 32824
rect 20088 32796 20729 32824
rect 17644 32784 17650 32796
rect 18782 32756 18788 32768
rect 17328 32728 18788 32756
rect 16393 32719 16451 32725
rect 18782 32716 18788 32728
rect 18840 32716 18846 32768
rect 19334 32716 19340 32768
rect 19392 32756 19398 32768
rect 19628 32756 19656 32796
rect 19392 32728 19656 32756
rect 19392 32716 19398 32728
rect 19794 32716 19800 32768
rect 19852 32756 19858 32768
rect 20088 32765 20116 32796
rect 20717 32793 20729 32796
rect 20763 32793 20775 32827
rect 20717 32787 20775 32793
rect 20901 32827 20959 32833
rect 20901 32793 20913 32827
rect 20947 32824 20959 32827
rect 21269 32827 21327 32833
rect 21269 32824 21281 32827
rect 20947 32796 21281 32824
rect 20947 32793 20959 32796
rect 20901 32787 20959 32793
rect 21269 32793 21281 32796
rect 21315 32793 21327 32827
rect 22020 32824 22048 32855
rect 22462 32852 22468 32904
rect 22520 32852 22526 32904
rect 23032 32892 23060 32932
rect 23216 32901 23244 32932
rect 23290 32920 23296 32932
rect 23348 32920 23354 32972
rect 23385 32963 23443 32969
rect 23385 32929 23397 32963
rect 23431 32960 23443 32963
rect 23431 32932 24624 32960
rect 23431 32929 23443 32932
rect 23385 32923 23443 32929
rect 22756 32864 23060 32892
rect 23109 32895 23167 32901
rect 22756 32836 22784 32864
rect 23109 32861 23121 32895
rect 23155 32861 23167 32895
rect 23109 32855 23167 32861
rect 23201 32895 23259 32901
rect 23201 32861 23213 32895
rect 23247 32861 23259 32895
rect 23201 32855 23259 32861
rect 22738 32824 22744 32836
rect 22020 32796 22744 32824
rect 21269 32787 21327 32793
rect 22738 32784 22744 32796
rect 22796 32784 22802 32836
rect 23124 32824 23152 32855
rect 23842 32852 23848 32904
rect 23900 32892 23906 32904
rect 24596 32901 24624 32932
rect 24029 32895 24087 32901
rect 24029 32892 24041 32895
rect 23900 32864 24041 32892
rect 23900 32852 23906 32864
rect 24029 32861 24041 32864
rect 24075 32861 24087 32895
rect 24029 32855 24087 32861
rect 24581 32895 24639 32901
rect 24581 32861 24593 32895
rect 24627 32861 24639 32895
rect 24581 32855 24639 32861
rect 25314 32852 25320 32904
rect 25372 32852 25378 32904
rect 25498 32824 25504 32836
rect 23124 32796 25504 32824
rect 25498 32784 25504 32796
rect 25556 32784 25562 32836
rect 20073 32759 20131 32765
rect 20073 32756 20085 32759
rect 19852 32728 20085 32756
rect 19852 32716 19858 32728
rect 20073 32725 20085 32728
rect 20119 32725 20131 32759
rect 20073 32719 20131 32725
rect 20165 32759 20223 32765
rect 20165 32725 20177 32759
rect 20211 32756 20223 32759
rect 20254 32756 20260 32768
rect 20211 32728 20260 32756
rect 20211 32725 20223 32728
rect 20165 32719 20223 32725
rect 20254 32716 20260 32728
rect 20312 32716 20318 32768
rect 23474 32716 23480 32768
rect 23532 32716 23538 32768
rect 24394 32716 24400 32768
rect 24452 32716 24458 32768
rect 1104 32666 35027 32688
rect 1104 32614 9390 32666
rect 9442 32614 9454 32666
rect 9506 32614 9518 32666
rect 9570 32614 9582 32666
rect 9634 32614 9646 32666
rect 9698 32614 17831 32666
rect 17883 32614 17895 32666
rect 17947 32614 17959 32666
rect 18011 32614 18023 32666
rect 18075 32614 18087 32666
rect 18139 32614 26272 32666
rect 26324 32614 26336 32666
rect 26388 32614 26400 32666
rect 26452 32614 26464 32666
rect 26516 32614 26528 32666
rect 26580 32614 34713 32666
rect 34765 32614 34777 32666
rect 34829 32614 34841 32666
rect 34893 32614 34905 32666
rect 34957 32614 34969 32666
rect 35021 32614 35027 32666
rect 1104 32592 35027 32614
rect 7653 32555 7711 32561
rect 7653 32521 7665 32555
rect 7699 32552 7711 32555
rect 7699 32524 8984 32552
rect 7699 32521 7711 32524
rect 7653 32515 7711 32521
rect 8478 32484 8484 32496
rect 7392 32456 8484 32484
rect 7392 32425 7420 32456
rect 8478 32444 8484 32456
rect 8536 32444 8542 32496
rect 7377 32419 7435 32425
rect 7377 32385 7389 32419
rect 7423 32385 7435 32419
rect 7377 32379 7435 32385
rect 7834 32376 7840 32428
rect 7892 32376 7898 32428
rect 7926 32376 7932 32428
rect 7984 32376 7990 32428
rect 8021 32419 8079 32425
rect 8021 32385 8033 32419
rect 8067 32416 8079 32419
rect 8110 32416 8116 32428
rect 8067 32388 8116 32416
rect 8067 32385 8079 32388
rect 8021 32379 8079 32385
rect 8110 32376 8116 32388
rect 8168 32416 8174 32428
rect 8168 32388 8248 32416
rect 8168 32376 8174 32388
rect 8220 32348 8248 32388
rect 8386 32348 8392 32360
rect 8220 32320 8392 32348
rect 8386 32308 8392 32320
rect 8444 32308 8450 32360
rect 8846 32348 8852 32360
rect 8772 32320 8852 32348
rect 7561 32283 7619 32289
rect 7561 32249 7573 32283
rect 7607 32280 7619 32283
rect 8205 32283 8263 32289
rect 7607 32252 8156 32280
rect 7607 32249 7619 32252
rect 7561 32243 7619 32249
rect 8128 32212 8156 32252
rect 8205 32249 8217 32283
rect 8251 32280 8263 32283
rect 8772 32280 8800 32320
rect 8846 32308 8852 32320
rect 8904 32308 8910 32360
rect 8956 32348 8984 32524
rect 10226 32512 10232 32564
rect 10284 32512 10290 32564
rect 10778 32512 10784 32564
rect 10836 32552 10842 32564
rect 10836 32524 11284 32552
rect 10836 32512 10842 32524
rect 9033 32487 9091 32493
rect 9033 32453 9045 32487
rect 9079 32484 9091 32487
rect 9122 32484 9128 32496
rect 9079 32456 9128 32484
rect 9079 32453 9091 32456
rect 9033 32447 9091 32453
rect 9122 32444 9128 32456
rect 9180 32444 9186 32496
rect 9769 32487 9827 32493
rect 9769 32484 9781 32487
rect 9508 32456 9781 32484
rect 9306 32376 9312 32428
rect 9364 32376 9370 32428
rect 9508 32425 9536 32456
rect 9769 32453 9781 32456
rect 9815 32453 9827 32487
rect 9769 32447 9827 32453
rect 9858 32444 9864 32496
rect 9916 32484 9922 32496
rect 10321 32487 10379 32493
rect 9916 32456 10180 32484
rect 9916 32444 9922 32456
rect 9401 32419 9459 32425
rect 9401 32385 9413 32419
rect 9447 32385 9459 32419
rect 9401 32379 9459 32385
rect 9493 32419 9551 32425
rect 9493 32385 9505 32419
rect 9539 32385 9551 32419
rect 9493 32379 9551 32385
rect 9416 32348 9444 32379
rect 9674 32376 9680 32428
rect 9732 32376 9738 32428
rect 9950 32376 9956 32428
rect 10008 32376 10014 32428
rect 10042 32376 10048 32428
rect 10100 32376 10106 32428
rect 10152 32416 10180 32456
rect 10321 32453 10333 32487
rect 10367 32484 10379 32487
rect 10594 32484 10600 32496
rect 10367 32456 10600 32484
rect 10367 32453 10379 32456
rect 10321 32447 10379 32453
rect 10594 32444 10600 32456
rect 10652 32444 10658 32496
rect 10686 32444 10692 32496
rect 10744 32484 10750 32496
rect 11146 32484 11152 32496
rect 10744 32456 11152 32484
rect 10744 32444 10750 32456
rect 10413 32419 10471 32425
rect 10336 32416 10425 32419
rect 10152 32391 10425 32416
rect 10152 32388 10364 32391
rect 10413 32385 10425 32391
rect 10459 32385 10471 32419
rect 10413 32379 10471 32385
rect 10502 32376 10508 32428
rect 10560 32416 10566 32428
rect 10796 32425 10824 32456
rect 11146 32444 11152 32456
rect 11204 32444 11210 32496
rect 10781 32419 10839 32425
rect 10560 32388 10732 32416
rect 10560 32376 10566 32388
rect 10704 32348 10732 32388
rect 10781 32385 10793 32419
rect 10827 32385 10839 32419
rect 10781 32379 10839 32385
rect 10870 32376 10876 32428
rect 10928 32376 10934 32428
rect 11256 32425 11284 32524
rect 11514 32512 11520 32564
rect 11572 32552 11578 32564
rect 11572 32524 12434 32552
rect 11572 32512 11578 32524
rect 11241 32419 11299 32425
rect 11241 32385 11253 32419
rect 11287 32385 11299 32419
rect 12406 32416 12434 32524
rect 13354 32512 13360 32564
rect 13412 32512 13418 32564
rect 13998 32512 14004 32564
rect 14056 32512 14062 32564
rect 14185 32555 14243 32561
rect 14185 32521 14197 32555
rect 14231 32552 14243 32555
rect 14642 32552 14648 32564
rect 14231 32524 14648 32552
rect 14231 32521 14243 32524
rect 14185 32515 14243 32521
rect 14642 32512 14648 32524
rect 14700 32512 14706 32564
rect 14734 32512 14740 32564
rect 14792 32512 14798 32564
rect 14826 32512 14832 32564
rect 14884 32552 14890 32564
rect 14884 32524 14964 32552
rect 14884 32512 14890 32524
rect 13446 32444 13452 32496
rect 13504 32484 13510 32496
rect 14016 32484 14044 32512
rect 14461 32487 14519 32493
rect 14461 32484 14473 32487
rect 13504 32456 13768 32484
rect 13504 32444 13510 32456
rect 13740 32425 13768 32456
rect 13832 32456 14044 32484
rect 14200 32456 14473 32484
rect 13832 32425 13860 32456
rect 14200 32428 14228 32456
rect 14461 32453 14473 32456
rect 14507 32453 14519 32487
rect 14752 32484 14780 32512
rect 14461 32447 14519 32453
rect 14660 32456 14780 32484
rect 12630 32419 12688 32425
rect 12630 32416 12642 32419
rect 12406 32388 12642 32416
rect 11241 32379 11299 32385
rect 12630 32385 12642 32388
rect 12676 32385 12688 32419
rect 12630 32379 12688 32385
rect 13633 32419 13691 32425
rect 13633 32385 13645 32419
rect 13679 32385 13691 32419
rect 13633 32379 13691 32385
rect 13725 32419 13783 32425
rect 13725 32385 13737 32419
rect 13771 32385 13783 32419
rect 13725 32379 13783 32385
rect 13817 32419 13875 32425
rect 13817 32385 13829 32419
rect 13863 32385 13875 32419
rect 13817 32379 13875 32385
rect 14001 32419 14059 32425
rect 14001 32385 14013 32419
rect 14047 32385 14059 32419
rect 14001 32379 14059 32385
rect 11057 32351 11115 32357
rect 11057 32348 11069 32351
rect 8956 32320 9352 32348
rect 9416 32340 10088 32348
rect 9416 32320 10226 32340
rect 10704 32320 11069 32348
rect 9214 32280 9220 32292
rect 8251 32252 8800 32280
rect 8864 32252 9220 32280
rect 8251 32249 8263 32252
rect 8205 32243 8263 32249
rect 8864 32212 8892 32252
rect 9214 32240 9220 32252
rect 9272 32240 9278 32292
rect 8128 32184 8892 32212
rect 8938 32172 8944 32224
rect 8996 32172 9002 32224
rect 9324 32212 9352 32320
rect 10060 32312 10226 32320
rect 10198 32280 10226 32312
rect 11057 32317 11069 32320
rect 11103 32317 11115 32351
rect 11057 32311 11115 32317
rect 12897 32351 12955 32357
rect 12897 32317 12909 32351
rect 12943 32317 12955 32351
rect 13648 32348 13676 32379
rect 14016 32348 14044 32379
rect 14090 32376 14096 32428
rect 14148 32376 14154 32428
rect 14182 32376 14188 32428
rect 14240 32376 14246 32428
rect 14660 32425 14688 32456
rect 14369 32419 14427 32425
rect 14369 32385 14381 32419
rect 14415 32385 14427 32419
rect 14369 32379 14427 32385
rect 14645 32419 14703 32425
rect 14645 32385 14657 32419
rect 14691 32385 14703 32419
rect 14645 32379 14703 32385
rect 14737 32419 14795 32425
rect 14737 32385 14749 32419
rect 14783 32385 14795 32419
rect 14737 32379 14795 32385
rect 14274 32348 14280 32360
rect 13648 32320 13768 32348
rect 14016 32320 14280 32348
rect 12897 32311 12955 32317
rect 11072 32280 11100 32311
rect 11517 32283 11575 32289
rect 11517 32280 11529 32283
rect 10198 32252 10548 32280
rect 11072 32252 11529 32280
rect 9858 32212 9864 32224
rect 9324 32184 9864 32212
rect 9858 32172 9864 32184
rect 9916 32172 9922 32224
rect 10520 32221 10548 32252
rect 11517 32249 11529 32252
rect 11563 32249 11575 32283
rect 11517 32243 11575 32249
rect 10505 32215 10563 32221
rect 10505 32181 10517 32215
rect 10551 32181 10563 32215
rect 10505 32175 10563 32181
rect 10594 32172 10600 32224
rect 10652 32212 10658 32224
rect 10965 32215 11023 32221
rect 10965 32212 10977 32215
rect 10652 32184 10977 32212
rect 10652 32172 10658 32184
rect 10965 32181 10977 32184
rect 11011 32212 11023 32215
rect 11422 32212 11428 32224
rect 11011 32184 11428 32212
rect 11011 32181 11023 32184
rect 10965 32175 11023 32181
rect 11422 32172 11428 32184
rect 11480 32172 11486 32224
rect 12710 32172 12716 32224
rect 12768 32212 12774 32224
rect 12912 32212 12940 32311
rect 13740 32280 13768 32320
rect 14274 32308 14280 32320
rect 14332 32308 14338 32360
rect 14090 32280 14096 32292
rect 13740 32252 14096 32280
rect 14090 32240 14096 32252
rect 14148 32240 14154 32292
rect 14384 32280 14412 32379
rect 14752 32348 14780 32379
rect 14826 32376 14832 32428
rect 14884 32376 14890 32428
rect 14936 32348 14964 32524
rect 15470 32512 15476 32564
rect 15528 32512 15534 32564
rect 15654 32512 15660 32564
rect 15712 32512 15718 32564
rect 15749 32555 15807 32561
rect 15749 32521 15761 32555
rect 15795 32552 15807 32555
rect 16574 32552 16580 32564
rect 15795 32524 16580 32552
rect 15795 32521 15807 32524
rect 15749 32515 15807 32521
rect 16574 32512 16580 32524
rect 16632 32512 16638 32564
rect 18325 32555 18383 32561
rect 18325 32552 18337 32555
rect 17880 32524 18337 32552
rect 15010 32376 15016 32428
rect 15068 32416 15074 32428
rect 15488 32416 15516 32512
rect 15672 32484 15700 32512
rect 17497 32487 17555 32493
rect 17497 32484 17509 32487
rect 15672 32456 16068 32484
rect 15068 32388 15516 32416
rect 15068 32376 15074 32388
rect 15562 32376 15568 32428
rect 15620 32376 15626 32428
rect 15657 32419 15715 32425
rect 15657 32385 15669 32419
rect 15703 32385 15715 32419
rect 15657 32379 15715 32385
rect 14752 32320 14964 32348
rect 15102 32308 15108 32360
rect 15160 32348 15166 32360
rect 15286 32348 15292 32360
rect 15160 32320 15292 32348
rect 15160 32308 15166 32320
rect 15286 32308 15292 32320
rect 15344 32348 15350 32360
rect 15381 32351 15439 32357
rect 15381 32348 15393 32351
rect 15344 32320 15393 32348
rect 15344 32308 15350 32320
rect 15381 32317 15393 32320
rect 15427 32317 15439 32351
rect 15672 32348 15700 32379
rect 15746 32376 15752 32428
rect 15804 32416 15810 32428
rect 16040 32425 16068 32456
rect 16224 32456 17509 32484
rect 16224 32425 16252 32456
rect 17497 32453 17509 32456
rect 17543 32453 17555 32487
rect 17497 32447 17555 32453
rect 15933 32419 15991 32425
rect 15933 32416 15945 32419
rect 15804 32388 15945 32416
rect 15804 32376 15810 32388
rect 15933 32385 15945 32388
rect 15979 32385 15991 32419
rect 15933 32379 15991 32385
rect 16025 32419 16083 32425
rect 16025 32385 16037 32419
rect 16071 32385 16083 32419
rect 16025 32379 16083 32385
rect 16209 32419 16267 32425
rect 16209 32385 16221 32419
rect 16255 32385 16267 32419
rect 16209 32379 16267 32385
rect 16298 32376 16304 32428
rect 16356 32416 16362 32428
rect 16669 32419 16727 32425
rect 16669 32416 16681 32419
rect 16356 32388 16681 32416
rect 16356 32376 16362 32388
rect 16669 32385 16681 32388
rect 16715 32385 16727 32419
rect 16669 32379 16727 32385
rect 16761 32419 16819 32425
rect 16761 32385 16773 32419
rect 16807 32385 16819 32419
rect 16945 32419 17003 32425
rect 16945 32416 16957 32419
rect 16761 32379 16819 32385
rect 16868 32388 16957 32416
rect 15838 32348 15844 32360
rect 15672 32320 15844 32348
rect 15381 32311 15439 32317
rect 15838 32308 15844 32320
rect 15896 32348 15902 32360
rect 16117 32351 16175 32357
rect 16117 32348 16129 32351
rect 15896 32320 16129 32348
rect 15896 32308 15902 32320
rect 16117 32317 16129 32320
rect 16163 32348 16175 32351
rect 16776 32348 16804 32379
rect 16163 32320 16804 32348
rect 16163 32317 16175 32320
rect 16117 32311 16175 32317
rect 15473 32283 15531 32289
rect 14384 32252 15424 32280
rect 12768 32184 12940 32212
rect 12768 32172 12774 32184
rect 14366 32172 14372 32224
rect 14424 32172 14430 32224
rect 14461 32215 14519 32221
rect 14461 32181 14473 32215
rect 14507 32212 14519 32215
rect 14550 32212 14556 32224
rect 14507 32184 14556 32212
rect 14507 32181 14519 32184
rect 14461 32175 14519 32181
rect 14550 32172 14556 32184
rect 14608 32172 14614 32224
rect 15396 32212 15424 32252
rect 15473 32249 15485 32283
rect 15519 32280 15531 32283
rect 16868 32280 16896 32388
rect 16945 32385 16957 32388
rect 16991 32385 17003 32419
rect 16945 32379 17003 32385
rect 17126 32376 17132 32428
rect 17184 32376 17190 32428
rect 17218 32376 17224 32428
rect 17276 32376 17282 32428
rect 17310 32376 17316 32428
rect 17368 32376 17374 32428
rect 17880 32425 17908 32524
rect 18325 32521 18337 32524
rect 18371 32521 18383 32555
rect 18325 32515 18383 32521
rect 18782 32512 18788 32564
rect 18840 32512 18846 32564
rect 19889 32555 19947 32561
rect 19889 32521 19901 32555
rect 19935 32552 19947 32555
rect 20346 32552 20352 32564
rect 19935 32524 20352 32552
rect 19935 32521 19947 32524
rect 19889 32515 19947 32521
rect 18800 32484 18828 32512
rect 19904 32484 19932 32515
rect 20346 32512 20352 32524
rect 20404 32512 20410 32564
rect 23658 32512 23664 32564
rect 23716 32512 23722 32564
rect 23842 32512 23848 32564
rect 23900 32512 23906 32564
rect 24026 32512 24032 32564
rect 24084 32512 24090 32564
rect 24394 32512 24400 32564
rect 24452 32512 24458 32564
rect 24486 32512 24492 32564
rect 24544 32552 24550 32564
rect 25314 32552 25320 32564
rect 24544 32524 25320 32552
rect 24544 32512 24550 32524
rect 25314 32512 25320 32524
rect 25372 32552 25378 32564
rect 25409 32555 25467 32561
rect 25409 32552 25421 32555
rect 25372 32524 25421 32552
rect 25372 32512 25378 32524
rect 25409 32521 25421 32524
rect 25455 32521 25467 32555
rect 25409 32515 25467 32521
rect 25498 32512 25504 32564
rect 25556 32512 25562 32564
rect 23293 32487 23351 32493
rect 23293 32484 23305 32487
rect 18800 32456 19104 32484
rect 17865 32419 17923 32425
rect 17865 32416 17877 32419
rect 17696 32388 17877 32416
rect 17144 32348 17172 32376
rect 17696 32360 17724 32388
rect 17865 32385 17877 32388
rect 17911 32385 17923 32419
rect 17865 32379 17923 32385
rect 18693 32419 18751 32425
rect 18693 32385 18705 32419
rect 18739 32416 18751 32419
rect 18782 32416 18788 32428
rect 18739 32388 18788 32416
rect 18739 32385 18751 32388
rect 18693 32379 18751 32385
rect 18782 32376 18788 32388
rect 18840 32416 18846 32428
rect 19076 32425 19104 32456
rect 19536 32456 19932 32484
rect 23032 32456 23305 32484
rect 18969 32419 19027 32425
rect 18969 32416 18981 32419
rect 18840 32388 18981 32416
rect 18840 32376 18846 32388
rect 18969 32385 18981 32388
rect 19015 32385 19027 32419
rect 18969 32379 19027 32385
rect 19061 32419 19119 32425
rect 19061 32385 19073 32419
rect 19107 32385 19119 32419
rect 19061 32379 19119 32385
rect 19337 32419 19395 32425
rect 19337 32385 19349 32419
rect 19383 32416 19395 32419
rect 19426 32416 19432 32428
rect 19383 32388 19432 32416
rect 19383 32385 19395 32388
rect 19337 32379 19395 32385
rect 19426 32376 19432 32388
rect 19484 32376 19490 32428
rect 19536 32425 19564 32456
rect 19521 32419 19579 32425
rect 19521 32385 19533 32419
rect 19567 32385 19579 32419
rect 19521 32379 19579 32385
rect 19610 32376 19616 32428
rect 19668 32425 19674 32428
rect 19668 32419 19717 32425
rect 19668 32385 19671 32419
rect 19705 32385 19717 32419
rect 19668 32379 19717 32385
rect 19668 32376 19674 32379
rect 19794 32376 19800 32428
rect 19852 32376 19858 32428
rect 20070 32376 20076 32428
rect 20128 32416 20134 32428
rect 20257 32419 20315 32425
rect 20128 32388 20208 32416
rect 20128 32376 20134 32388
rect 17497 32351 17555 32357
rect 17497 32348 17509 32351
rect 17144 32320 17509 32348
rect 17497 32317 17509 32320
rect 17543 32317 17555 32351
rect 17497 32311 17555 32317
rect 15519 32252 15976 32280
rect 15519 32249 15531 32252
rect 15473 32243 15531 32249
rect 15654 32212 15660 32224
rect 15396 32184 15660 32212
rect 15654 32172 15660 32184
rect 15712 32172 15718 32224
rect 15948 32212 15976 32252
rect 16776 32252 16896 32280
rect 17512 32280 17540 32311
rect 17678 32308 17684 32360
rect 17736 32308 17742 32360
rect 17770 32308 17776 32360
rect 17828 32308 17834 32360
rect 18230 32308 18236 32360
rect 18288 32308 18294 32360
rect 20180 32357 20208 32388
rect 20257 32385 20269 32419
rect 20303 32416 20315 32419
rect 20533 32419 20591 32425
rect 20533 32416 20545 32419
rect 20303 32388 20545 32416
rect 20303 32385 20315 32388
rect 20257 32379 20315 32385
rect 20533 32385 20545 32388
rect 20579 32385 20591 32419
rect 20533 32379 20591 32385
rect 18601 32351 18659 32357
rect 18601 32317 18613 32351
rect 18647 32348 18659 32351
rect 19245 32351 19303 32357
rect 19245 32348 19257 32351
rect 18647 32320 19257 32348
rect 18647 32317 18659 32320
rect 18601 32311 18659 32317
rect 18616 32280 18644 32311
rect 18984 32292 19012 32320
rect 19245 32317 19257 32320
rect 19291 32317 19303 32351
rect 20165 32351 20223 32357
rect 20165 32348 20177 32351
rect 19245 32311 19303 32317
rect 19418 32320 20177 32348
rect 17512 32252 18644 32280
rect 16776 32212 16804 32252
rect 18966 32240 18972 32292
rect 19024 32240 19030 32292
rect 19150 32240 19156 32292
rect 19208 32240 19214 32292
rect 19260 32280 19288 32311
rect 19418 32280 19446 32320
rect 20165 32317 20177 32320
rect 20211 32317 20223 32351
rect 20165 32311 20223 32317
rect 19260 32252 19446 32280
rect 20070 32240 20076 32292
rect 20128 32280 20134 32292
rect 20272 32280 20300 32379
rect 22830 32376 22836 32428
rect 22888 32376 22894 32428
rect 22922 32376 22928 32428
rect 22980 32376 22986 32428
rect 23032 32425 23060 32456
rect 23293 32453 23305 32456
rect 23339 32453 23351 32487
rect 23293 32447 23351 32453
rect 23382 32444 23388 32496
rect 23440 32484 23446 32496
rect 23860 32484 23888 32512
rect 23440 32456 23888 32484
rect 23440 32444 23446 32456
rect 23017 32419 23075 32425
rect 23017 32385 23029 32419
rect 23063 32385 23075 32419
rect 23017 32379 23075 32385
rect 23198 32376 23204 32428
rect 23256 32376 23262 32428
rect 24044 32425 24072 32512
rect 24296 32487 24354 32493
rect 24296 32453 24308 32487
rect 24342 32484 24354 32487
rect 24412 32484 24440 32512
rect 24342 32456 24440 32484
rect 24342 32453 24354 32456
rect 24296 32447 24354 32453
rect 23569 32419 23627 32425
rect 23569 32385 23581 32419
rect 23615 32385 23627 32419
rect 23569 32379 23627 32385
rect 24029 32419 24087 32425
rect 24029 32385 24041 32419
rect 24075 32385 24087 32419
rect 24029 32379 24087 32385
rect 21082 32308 21088 32360
rect 21140 32308 21146 32360
rect 21913 32351 21971 32357
rect 21913 32317 21925 32351
rect 21959 32348 21971 32351
rect 22557 32351 22615 32357
rect 22557 32348 22569 32351
rect 21959 32320 22569 32348
rect 21959 32317 21971 32320
rect 21913 32311 21971 32317
rect 22557 32317 22569 32320
rect 22603 32317 22615 32351
rect 22557 32311 22615 32317
rect 23477 32351 23535 32357
rect 23477 32317 23489 32351
rect 23523 32317 23535 32351
rect 23477 32311 23535 32317
rect 20128 32252 20300 32280
rect 20128 32240 20134 32252
rect 21450 32240 21456 32292
rect 21508 32280 21514 32292
rect 23198 32280 23204 32292
rect 21508 32252 23204 32280
rect 21508 32240 21514 32252
rect 23198 32240 23204 32252
rect 23256 32280 23262 32292
rect 23492 32280 23520 32311
rect 23256 32252 23520 32280
rect 23256 32240 23262 32252
rect 15948 32184 16804 32212
rect 16850 32172 16856 32224
rect 16908 32212 16914 32224
rect 17129 32215 17187 32221
rect 17129 32212 17141 32215
rect 16908 32184 17141 32212
rect 16908 32172 16914 32184
rect 17129 32181 17141 32184
rect 17175 32181 17187 32215
rect 17129 32175 17187 32181
rect 17586 32172 17592 32224
rect 17644 32172 17650 32224
rect 19426 32172 19432 32224
rect 19484 32172 19490 32224
rect 22462 32172 22468 32224
rect 22520 32172 22526 32224
rect 23014 32172 23020 32224
rect 23072 32212 23078 32224
rect 23290 32212 23296 32224
rect 23072 32184 23296 32212
rect 23072 32172 23078 32184
rect 23290 32172 23296 32184
rect 23348 32212 23354 32224
rect 23584 32212 23612 32379
rect 23934 32308 23940 32360
rect 23992 32308 23998 32360
rect 26053 32351 26111 32357
rect 26053 32317 26065 32351
rect 26099 32317 26111 32351
rect 26053 32311 26111 32317
rect 23348 32184 23612 32212
rect 23348 32172 23354 32184
rect 25774 32172 25780 32224
rect 25832 32212 25838 32224
rect 26068 32212 26096 32311
rect 25832 32184 26096 32212
rect 25832 32172 25838 32184
rect 1104 32122 34868 32144
rect 1104 32070 5170 32122
rect 5222 32070 5234 32122
rect 5286 32070 5298 32122
rect 5350 32070 5362 32122
rect 5414 32070 5426 32122
rect 5478 32070 13611 32122
rect 13663 32070 13675 32122
rect 13727 32070 13739 32122
rect 13791 32070 13803 32122
rect 13855 32070 13867 32122
rect 13919 32070 22052 32122
rect 22104 32070 22116 32122
rect 22168 32070 22180 32122
rect 22232 32070 22244 32122
rect 22296 32070 22308 32122
rect 22360 32070 30493 32122
rect 30545 32070 30557 32122
rect 30609 32070 30621 32122
rect 30673 32070 30685 32122
rect 30737 32070 30749 32122
rect 30801 32070 34868 32122
rect 1104 32048 34868 32070
rect 8757 32011 8815 32017
rect 8757 31977 8769 32011
rect 8803 32008 8815 32011
rect 8846 32008 8852 32020
rect 8803 31980 8852 32008
rect 8803 31977 8815 31980
rect 8757 31971 8815 31977
rect 8846 31968 8852 31980
rect 8904 31968 8910 32020
rect 9674 31968 9680 32020
rect 9732 32008 9738 32020
rect 11054 32008 11060 32020
rect 9732 31980 11060 32008
rect 9732 31968 9738 31980
rect 11054 31968 11060 31980
rect 11112 31968 11118 32020
rect 11146 31968 11152 32020
rect 11204 32008 11210 32020
rect 12253 32011 12311 32017
rect 12253 32008 12265 32011
rect 11204 31980 12265 32008
rect 11204 31968 11210 31980
rect 12253 31977 12265 31980
rect 12299 31977 12311 32011
rect 12253 31971 12311 31977
rect 10318 31900 10324 31952
rect 10376 31900 10382 31952
rect 12268 31884 12296 31971
rect 14090 31968 14096 32020
rect 14148 32008 14154 32020
rect 14826 32008 14832 32020
rect 14148 31980 14832 32008
rect 14148 31968 14154 31980
rect 14826 31968 14832 31980
rect 14884 31968 14890 32020
rect 15838 31968 15844 32020
rect 15896 31968 15902 32020
rect 18414 32008 18420 32020
rect 16868 31980 18420 32008
rect 14553 31943 14611 31949
rect 14553 31909 14565 31943
rect 14599 31940 14611 31943
rect 14642 31940 14648 31952
rect 14599 31912 14648 31940
rect 14599 31909 14611 31912
rect 14553 31903 14611 31909
rect 14642 31900 14648 31912
rect 14700 31900 14706 31952
rect 7374 31832 7380 31884
rect 7432 31832 7438 31884
rect 12250 31832 12256 31884
rect 12308 31872 12314 31884
rect 12897 31875 12955 31881
rect 12897 31872 12909 31875
rect 12308 31844 12909 31872
rect 12308 31832 12314 31844
rect 12897 31841 12909 31844
rect 12943 31841 12955 31875
rect 12897 31835 12955 31841
rect 13814 31832 13820 31884
rect 13872 31832 13878 31884
rect 16206 31832 16212 31884
rect 16264 31832 16270 31884
rect 7392 31804 7420 31832
rect 8941 31807 8999 31813
rect 8941 31804 8953 31807
rect 7392 31776 8953 31804
rect 8941 31773 8953 31776
rect 8987 31804 8999 31807
rect 9030 31804 9036 31816
rect 8987 31776 9036 31804
rect 8987 31773 8999 31776
rect 8941 31767 8999 31773
rect 9030 31764 9036 31776
rect 9088 31764 9094 31816
rect 9214 31813 9220 31816
rect 9208 31804 9220 31813
rect 9175 31776 9220 31804
rect 9208 31767 9220 31776
rect 9214 31764 9220 31767
rect 9272 31764 9278 31816
rect 10873 31807 10931 31813
rect 10873 31773 10885 31807
rect 10919 31804 10931 31807
rect 12710 31804 12716 31816
rect 10919 31776 12716 31804
rect 10919 31773 10931 31776
rect 10873 31767 10931 31773
rect 12710 31764 12716 31776
rect 12768 31764 12774 31816
rect 13446 31764 13452 31816
rect 13504 31804 13510 31816
rect 14090 31804 14096 31816
rect 13504 31776 14096 31804
rect 13504 31764 13510 31776
rect 14090 31764 14096 31776
rect 14148 31764 14154 31816
rect 14182 31764 14188 31816
rect 14240 31804 14246 31816
rect 14369 31807 14427 31813
rect 14369 31804 14381 31807
rect 14240 31776 14381 31804
rect 14240 31764 14246 31776
rect 14369 31773 14381 31776
rect 14415 31773 14427 31807
rect 14369 31767 14427 31773
rect 15930 31764 15936 31816
rect 15988 31804 15994 31816
rect 16117 31807 16175 31813
rect 16117 31804 16129 31807
rect 15988 31776 16129 31804
rect 15988 31764 15994 31776
rect 16117 31773 16129 31776
rect 16163 31804 16175 31807
rect 16163 31776 16574 31804
rect 16163 31773 16175 31776
rect 16117 31767 16175 31773
rect 7644 31739 7702 31745
rect 7644 31705 7656 31739
rect 7690 31736 7702 31739
rect 8018 31736 8024 31748
rect 7690 31708 8024 31736
rect 7690 31705 7702 31708
rect 7644 31699 7702 31705
rect 8018 31696 8024 31708
rect 8076 31696 8082 31748
rect 11140 31739 11198 31745
rect 11140 31705 11152 31739
rect 11186 31736 11198 31739
rect 11330 31736 11336 31748
rect 11186 31708 11336 31736
rect 11186 31705 11198 31708
rect 11140 31699 11198 31705
rect 11330 31696 11336 31708
rect 11388 31696 11394 31748
rect 12342 31628 12348 31680
rect 12400 31628 12406 31680
rect 13262 31628 13268 31680
rect 13320 31628 13326 31680
rect 14274 31628 14280 31680
rect 14332 31668 14338 31680
rect 14734 31668 14740 31680
rect 14332 31640 14740 31668
rect 14332 31628 14338 31640
rect 14734 31628 14740 31640
rect 14792 31668 14798 31680
rect 15470 31668 15476 31680
rect 14792 31640 15476 31668
rect 14792 31628 14798 31640
rect 15470 31628 15476 31640
rect 15528 31628 15534 31680
rect 16546 31668 16574 31776
rect 16666 31764 16672 31816
rect 16724 31764 16730 31816
rect 16868 31813 16896 31980
rect 18414 31968 18420 31980
rect 18472 31968 18478 32020
rect 18782 32008 18788 32020
rect 18524 31980 18788 32008
rect 17126 31900 17132 31952
rect 17184 31940 17190 31952
rect 17221 31943 17279 31949
rect 17221 31940 17233 31943
rect 17184 31912 17233 31940
rect 17184 31900 17190 31912
rect 17221 31909 17233 31912
rect 17267 31909 17279 31943
rect 17678 31940 17684 31952
rect 17221 31903 17279 31909
rect 17512 31912 17684 31940
rect 16853 31807 16911 31813
rect 16853 31773 16865 31807
rect 16899 31773 16911 31807
rect 16853 31767 16911 31773
rect 17034 31764 17040 31816
rect 17092 31764 17098 31816
rect 17512 31813 17540 31912
rect 17678 31900 17684 31912
rect 17736 31900 17742 31952
rect 17770 31900 17776 31952
rect 17828 31900 17834 31952
rect 17957 31943 18015 31949
rect 17957 31909 17969 31943
rect 18003 31940 18015 31943
rect 18230 31940 18236 31952
rect 18003 31912 18236 31940
rect 18003 31909 18015 31912
rect 17957 31903 18015 31909
rect 18230 31900 18236 31912
rect 18288 31940 18294 31952
rect 18524 31940 18552 31980
rect 18782 31968 18788 31980
rect 18840 31968 18846 32020
rect 19702 31968 19708 32020
rect 19760 32008 19766 32020
rect 20254 32008 20260 32020
rect 19760 31980 20260 32008
rect 19760 31968 19766 31980
rect 20254 31968 20260 31980
rect 20312 31968 20318 32020
rect 21174 31968 21180 32020
rect 21232 31968 21238 32020
rect 21361 32011 21419 32017
rect 21361 31977 21373 32011
rect 21407 32008 21419 32011
rect 22094 32008 22100 32020
rect 21407 31980 22100 32008
rect 21407 31977 21419 31980
rect 21361 31971 21419 31977
rect 22094 31968 22100 31980
rect 22152 31968 22158 32020
rect 22922 31968 22928 32020
rect 22980 31968 22986 32020
rect 23382 31968 23388 32020
rect 23440 31968 23446 32020
rect 23477 32011 23535 32017
rect 23477 31977 23489 32011
rect 23523 32008 23535 32011
rect 23658 32008 23664 32020
rect 23523 31980 23664 32008
rect 23523 31977 23535 31980
rect 23477 31971 23535 31977
rect 23658 31968 23664 31980
rect 23716 31968 23722 32020
rect 24026 31968 24032 32020
rect 24084 31968 24090 32020
rect 24213 32011 24271 32017
rect 24213 31977 24225 32011
rect 24259 32008 24271 32011
rect 24302 32008 24308 32020
rect 24259 31980 24308 32008
rect 24259 31977 24271 31980
rect 24213 31971 24271 31977
rect 24302 31968 24308 31980
rect 24360 31968 24366 32020
rect 24762 31968 24768 32020
rect 24820 32008 24826 32020
rect 25774 32008 25780 32020
rect 24820 31980 25780 32008
rect 24820 31968 24826 31980
rect 25774 31968 25780 31980
rect 25832 31968 25838 32020
rect 18288 31912 18552 31940
rect 18288 31900 18294 31912
rect 18598 31900 18604 31952
rect 18656 31940 18662 31952
rect 21192 31940 21220 31968
rect 18656 31912 21220 31940
rect 18656 31900 18662 31912
rect 21450 31900 21456 31952
rect 21508 31900 21514 31952
rect 23293 31943 23351 31949
rect 23293 31909 23305 31943
rect 23339 31940 23351 31943
rect 23753 31943 23811 31949
rect 23753 31940 23765 31943
rect 23339 31912 23765 31940
rect 23339 31909 23351 31912
rect 23293 31903 23351 31909
rect 23753 31909 23765 31912
rect 23799 31909 23811 31943
rect 23753 31903 23811 31909
rect 17788 31872 17816 31900
rect 18509 31875 18567 31881
rect 18509 31872 18521 31875
rect 17696 31844 18521 31872
rect 17696 31813 17724 31844
rect 18509 31841 18521 31844
rect 18555 31841 18567 31875
rect 18509 31835 18567 31841
rect 19426 31832 19432 31884
rect 19484 31872 19490 31884
rect 19797 31875 19855 31881
rect 19797 31872 19809 31875
rect 19484 31844 19809 31872
rect 19484 31832 19490 31844
rect 19797 31841 19809 31844
rect 19843 31841 19855 31875
rect 19797 31835 19855 31841
rect 22833 31875 22891 31881
rect 22833 31841 22845 31875
rect 22879 31872 22891 31875
rect 24044 31872 24072 31968
rect 24397 31875 24455 31881
rect 24397 31872 24409 31875
rect 22879 31844 24409 31872
rect 22879 31841 22891 31844
rect 22833 31835 22891 31841
rect 24397 31841 24409 31844
rect 24443 31841 24455 31875
rect 24397 31835 24455 31841
rect 17497 31807 17555 31813
rect 17497 31773 17509 31807
rect 17543 31773 17555 31807
rect 17497 31767 17555 31773
rect 17681 31807 17739 31813
rect 17681 31773 17693 31807
rect 17727 31773 17739 31807
rect 17681 31767 17739 31773
rect 17773 31807 17831 31813
rect 17773 31773 17785 31807
rect 17819 31773 17831 31807
rect 17773 31767 17831 31773
rect 16942 31696 16948 31748
rect 17000 31696 17006 31748
rect 17218 31696 17224 31748
rect 17276 31696 17282 31748
rect 17788 31736 17816 31767
rect 18690 31764 18696 31816
rect 18748 31764 18754 31816
rect 18874 31804 18880 31816
rect 18800 31776 18880 31804
rect 18800 31748 18828 31776
rect 18874 31764 18880 31776
rect 18932 31764 18938 31816
rect 18966 31764 18972 31816
rect 19024 31764 19030 31816
rect 19518 31764 19524 31816
rect 19576 31764 19582 31816
rect 19702 31764 19708 31816
rect 19760 31764 19766 31816
rect 19889 31807 19947 31813
rect 19889 31804 19901 31807
rect 19812 31776 19901 31804
rect 17512 31708 17816 31736
rect 17236 31668 17264 31696
rect 17512 31680 17540 31708
rect 18506 31696 18512 31748
rect 18564 31696 18570 31748
rect 18782 31696 18788 31748
rect 18840 31696 18846 31748
rect 19812 31736 19840 31776
rect 19889 31773 19901 31776
rect 19935 31773 19947 31807
rect 19889 31767 19947 31773
rect 20070 31764 20076 31816
rect 20128 31764 20134 31816
rect 20257 31807 20315 31813
rect 20257 31773 20269 31807
rect 20303 31804 20315 31807
rect 20349 31807 20407 31813
rect 20349 31804 20361 31807
rect 20303 31776 20361 31804
rect 20303 31773 20315 31776
rect 20257 31767 20315 31773
rect 20349 31773 20361 31776
rect 20395 31773 20407 31807
rect 20349 31767 20407 31773
rect 21177 31807 21235 31813
rect 21177 31773 21189 31807
rect 21223 31804 21235 31807
rect 22848 31804 22876 31835
rect 21223 31776 21772 31804
rect 21223 31773 21235 31776
rect 21177 31767 21235 31773
rect 19260 31708 19840 31736
rect 16546 31640 17264 31668
rect 17494 31628 17500 31680
rect 17552 31628 17558 31680
rect 17586 31628 17592 31680
rect 17644 31628 17650 31680
rect 18524 31668 18552 31696
rect 19260 31668 19288 31708
rect 18524 31640 19288 31668
rect 20990 31628 20996 31680
rect 21048 31628 21054 31680
rect 21744 31668 21772 31776
rect 22112 31776 22876 31804
rect 21818 31696 21824 31748
rect 21876 31736 21882 31748
rect 22112 31736 22140 31776
rect 23198 31764 23204 31816
rect 23256 31764 23262 31816
rect 23290 31764 23296 31816
rect 23348 31764 23354 31816
rect 23661 31807 23719 31813
rect 23661 31773 23673 31807
rect 23707 31804 23719 31807
rect 23937 31807 23995 31813
rect 23707 31776 23741 31804
rect 23707 31773 23719 31776
rect 23661 31767 23719 31773
rect 23937 31773 23949 31807
rect 23983 31773 23995 31807
rect 23937 31767 23995 31773
rect 24029 31807 24087 31813
rect 24029 31773 24041 31807
rect 24075 31804 24087 31807
rect 24118 31804 24124 31816
rect 24075 31776 24124 31804
rect 24075 31773 24087 31776
rect 24029 31767 24087 31773
rect 21876 31708 22140 31736
rect 21876 31696 21882 31708
rect 22554 31696 22560 31748
rect 22612 31745 22618 31748
rect 22612 31699 22624 31745
rect 23308 31736 23336 31764
rect 23676 31736 23704 31767
rect 23952 31736 23980 31767
rect 24118 31764 24124 31776
rect 24176 31764 24182 31816
rect 24213 31807 24271 31813
rect 24213 31773 24225 31807
rect 24259 31804 24271 31807
rect 24486 31804 24492 31816
rect 24259 31776 24492 31804
rect 24259 31773 24271 31776
rect 24213 31767 24271 31773
rect 24486 31764 24492 31776
rect 24544 31764 24550 31816
rect 24642 31739 24700 31745
rect 24642 31736 24654 31739
rect 23308 31708 23704 31736
rect 23768 31708 23980 31736
rect 24044 31708 24654 31736
rect 22612 31696 22618 31699
rect 23768 31680 23796 31708
rect 22646 31668 22652 31680
rect 21744 31640 22652 31668
rect 22646 31628 22652 31640
rect 22704 31628 22710 31680
rect 23750 31628 23756 31680
rect 23808 31628 23814 31680
rect 23842 31628 23848 31680
rect 23900 31668 23906 31680
rect 24044 31668 24072 31708
rect 24642 31705 24654 31708
rect 24688 31705 24700 31739
rect 24642 31699 24700 31705
rect 23900 31640 24072 31668
rect 23900 31628 23906 31640
rect 1104 31578 35027 31600
rect 1104 31526 9390 31578
rect 9442 31526 9454 31578
rect 9506 31526 9518 31578
rect 9570 31526 9582 31578
rect 9634 31526 9646 31578
rect 9698 31526 17831 31578
rect 17883 31526 17895 31578
rect 17947 31526 17959 31578
rect 18011 31526 18023 31578
rect 18075 31526 18087 31578
rect 18139 31526 26272 31578
rect 26324 31526 26336 31578
rect 26388 31526 26400 31578
rect 26452 31526 26464 31578
rect 26516 31526 26528 31578
rect 26580 31526 34713 31578
rect 34765 31526 34777 31578
rect 34829 31526 34841 31578
rect 34893 31526 34905 31578
rect 34957 31526 34969 31578
rect 35021 31526 35027 31578
rect 1104 31504 35027 31526
rect 8018 31424 8024 31476
rect 8076 31424 8082 31476
rect 8478 31424 8484 31476
rect 8536 31464 8542 31476
rect 9493 31467 9551 31473
rect 9493 31464 9505 31467
rect 8536 31436 9505 31464
rect 8536 31424 8542 31436
rect 9493 31433 9505 31436
rect 9539 31433 9551 31467
rect 9493 31427 9551 31433
rect 11532 31436 13400 31464
rect 8938 31396 8944 31408
rect 8680 31368 8944 31396
rect 8205 31331 8263 31337
rect 8205 31297 8217 31331
rect 8251 31328 8263 31331
rect 8297 31331 8355 31337
rect 8297 31328 8309 31331
rect 8251 31300 8309 31328
rect 8251 31297 8263 31300
rect 8205 31291 8263 31297
rect 8297 31297 8309 31300
rect 8343 31297 8355 31331
rect 8297 31291 8355 31297
rect 8478 31288 8484 31340
rect 8536 31288 8542 31340
rect 8680 31337 8708 31368
rect 8938 31356 8944 31368
rect 8996 31356 9002 31408
rect 8665 31331 8723 31337
rect 8665 31297 8677 31331
rect 8711 31297 8723 31331
rect 8665 31291 8723 31297
rect 8754 31288 8760 31340
rect 8812 31288 8818 31340
rect 9677 31331 9735 31337
rect 9677 31328 9689 31331
rect 8864 31300 9689 31328
rect 8496 31260 8524 31288
rect 8864 31260 8892 31300
rect 9677 31297 9689 31300
rect 9723 31297 9735 31331
rect 9677 31291 9735 31297
rect 10226 31288 10232 31340
rect 10284 31288 10290 31340
rect 11054 31288 11060 31340
rect 11112 31328 11118 31340
rect 11532 31337 11560 31436
rect 12980 31399 13038 31405
rect 12980 31365 12992 31399
rect 13026 31396 13038 31399
rect 13262 31396 13268 31408
rect 13026 31368 13268 31396
rect 13026 31365 13038 31368
rect 12980 31359 13038 31365
rect 13262 31356 13268 31368
rect 13320 31356 13326 31408
rect 13372 31396 13400 31436
rect 13814 31424 13820 31476
rect 13872 31464 13878 31476
rect 14185 31467 14243 31473
rect 14185 31464 14197 31467
rect 13872 31436 14197 31464
rect 13872 31424 13878 31436
rect 14185 31433 14197 31436
rect 14231 31433 14243 31467
rect 14185 31427 14243 31433
rect 14550 31424 14556 31476
rect 14608 31464 14614 31476
rect 17129 31467 17187 31473
rect 14608 31436 15792 31464
rect 14608 31424 14614 31436
rect 14274 31396 14280 31408
rect 13372 31368 14280 31396
rect 14274 31356 14280 31368
rect 14332 31356 14338 31408
rect 15473 31399 15531 31405
rect 15473 31396 15485 31399
rect 14476 31368 15485 31396
rect 14476 31340 14504 31368
rect 15473 31365 15485 31368
rect 15519 31365 15531 31399
rect 15473 31359 15531 31365
rect 11517 31331 11575 31337
rect 11517 31328 11529 31331
rect 11112 31300 11529 31328
rect 11112 31288 11118 31300
rect 11517 31297 11529 31300
rect 11563 31297 11575 31331
rect 11517 31291 11575 31297
rect 11606 31288 11612 31340
rect 11664 31328 11670 31340
rect 11701 31331 11759 31337
rect 11701 31328 11713 31331
rect 11664 31300 11713 31328
rect 11664 31288 11670 31300
rect 11701 31297 11713 31300
rect 11747 31297 11759 31331
rect 11701 31291 11759 31297
rect 11790 31288 11796 31340
rect 11848 31288 11854 31340
rect 11885 31331 11943 31337
rect 11885 31297 11897 31331
rect 11931 31297 11943 31331
rect 11885 31291 11943 31297
rect 8496 31232 8892 31260
rect 9401 31263 9459 31269
rect 9401 31229 9413 31263
rect 9447 31260 9459 31263
rect 9861 31263 9919 31269
rect 9861 31260 9873 31263
rect 9447 31232 9873 31260
rect 9447 31229 9459 31232
rect 9401 31223 9459 31229
rect 9861 31229 9873 31232
rect 9907 31229 9919 31263
rect 9861 31223 9919 31229
rect 10502 31220 10508 31272
rect 10560 31220 10566 31272
rect 11900 31260 11928 31291
rect 12342 31288 12348 31340
rect 12400 31288 12406 31340
rect 12434 31288 12440 31340
rect 12492 31328 12498 31340
rect 13354 31328 13360 31340
rect 12492 31300 13360 31328
rect 12492 31288 12498 31300
rect 13354 31288 13360 31300
rect 13412 31328 13418 31340
rect 13412 31300 13768 31328
rect 13412 31288 13418 31300
rect 11164 31232 11928 31260
rect 11164 31136 11192 31232
rect 12710 31220 12716 31272
rect 12768 31220 12774 31272
rect 13740 31192 13768 31300
rect 13998 31288 14004 31340
rect 14056 31288 14062 31340
rect 14366 31288 14372 31340
rect 14424 31288 14430 31340
rect 14458 31288 14464 31340
rect 14516 31288 14522 31340
rect 14642 31288 14648 31340
rect 14700 31288 14706 31340
rect 14829 31331 14887 31337
rect 14829 31297 14841 31331
rect 14875 31297 14887 31331
rect 14829 31291 14887 31297
rect 14016 31260 14044 31288
rect 14553 31263 14611 31269
rect 14553 31260 14565 31263
rect 14016 31232 14565 31260
rect 14553 31229 14565 31232
rect 14599 31229 14611 31263
rect 14553 31223 14611 31229
rect 14568 31192 14596 31223
rect 14642 31192 14648 31204
rect 13740 31164 14320 31192
rect 14568 31164 14648 31192
rect 10042 31084 10048 31136
rect 10100 31084 10106 31136
rect 11146 31084 11152 31136
rect 11204 31084 11210 31136
rect 12161 31127 12219 31133
rect 12161 31093 12173 31127
rect 12207 31124 12219 31127
rect 12526 31124 12532 31136
rect 12207 31096 12532 31124
rect 12207 31093 12219 31096
rect 12161 31087 12219 31093
rect 12526 31084 12532 31096
rect 12584 31084 12590 31136
rect 12621 31127 12679 31133
rect 12621 31093 12633 31127
rect 12667 31124 12679 31127
rect 13446 31124 13452 31136
rect 12667 31096 13452 31124
rect 12667 31093 12679 31096
rect 12621 31087 12679 31093
rect 13446 31084 13452 31096
rect 13504 31084 13510 31136
rect 14093 31127 14151 31133
rect 14093 31093 14105 31127
rect 14139 31124 14151 31127
rect 14182 31124 14188 31136
rect 14139 31096 14188 31124
rect 14139 31093 14151 31096
rect 14093 31087 14151 31093
rect 14182 31084 14188 31096
rect 14240 31084 14246 31136
rect 14292 31124 14320 31164
rect 14642 31152 14648 31164
rect 14700 31152 14706 31204
rect 14844 31124 14872 31291
rect 15010 31288 15016 31340
rect 15068 31328 15074 31340
rect 15764 31337 15792 31436
rect 17129 31433 17141 31467
rect 17175 31464 17187 31467
rect 17218 31464 17224 31476
rect 17175 31436 17224 31464
rect 17175 31433 17187 31436
rect 17129 31427 17187 31433
rect 17218 31424 17224 31436
rect 17276 31424 17282 31476
rect 17586 31424 17592 31476
rect 17644 31424 17650 31476
rect 19610 31424 19616 31476
rect 19668 31464 19674 31476
rect 19889 31467 19947 31473
rect 19889 31464 19901 31467
rect 19668 31436 19901 31464
rect 19668 31424 19674 31436
rect 19889 31433 19901 31436
rect 19935 31464 19947 31467
rect 21082 31464 21088 31476
rect 19935 31436 21088 31464
rect 19935 31433 19947 31436
rect 19889 31427 19947 31433
rect 21082 31424 21088 31436
rect 21140 31424 21146 31476
rect 23201 31467 23259 31473
rect 23201 31433 23213 31467
rect 23247 31464 23259 31467
rect 23658 31464 23664 31476
rect 23247 31436 23664 31464
rect 23247 31433 23259 31436
rect 23201 31427 23259 31433
rect 23658 31424 23664 31436
rect 23716 31424 23722 31476
rect 23842 31424 23848 31476
rect 23900 31424 23906 31476
rect 23934 31424 23940 31476
rect 23992 31424 23998 31476
rect 24118 31424 24124 31476
rect 24176 31464 24182 31476
rect 24213 31467 24271 31473
rect 24213 31464 24225 31467
rect 24176 31436 24225 31464
rect 24176 31424 24182 31436
rect 24213 31433 24225 31436
rect 24259 31433 24271 31467
rect 24213 31427 24271 31433
rect 24302 31424 24308 31476
rect 24360 31424 24366 31476
rect 24486 31424 24492 31476
rect 24544 31424 24550 31476
rect 16942 31356 16948 31408
rect 17000 31396 17006 31408
rect 17604 31396 17632 31424
rect 18506 31396 18512 31408
rect 17000 31368 17356 31396
rect 17604 31368 17816 31396
rect 17000 31356 17006 31368
rect 17328 31337 17356 31368
rect 17788 31337 17816 31368
rect 17972 31368 18512 31396
rect 15289 31331 15347 31337
rect 15289 31328 15301 31331
rect 15068 31300 15301 31328
rect 15068 31288 15074 31300
rect 15289 31297 15301 31300
rect 15335 31297 15347 31331
rect 15289 31291 15347 31297
rect 15749 31331 15807 31337
rect 15749 31297 15761 31331
rect 15795 31297 15807 31331
rect 15749 31291 15807 31297
rect 15841 31331 15899 31337
rect 15841 31297 15853 31331
rect 15887 31297 15899 31331
rect 15841 31291 15899 31297
rect 16025 31331 16083 31337
rect 16025 31297 16037 31331
rect 16071 31297 16083 31331
rect 16025 31291 16083 31297
rect 17313 31331 17371 31337
rect 17313 31297 17325 31331
rect 17359 31297 17371 31331
rect 17313 31291 17371 31297
rect 17589 31331 17647 31337
rect 17589 31297 17601 31331
rect 17635 31297 17647 31331
rect 17589 31291 17647 31297
rect 17773 31331 17831 31337
rect 17773 31297 17785 31331
rect 17819 31297 17831 31331
rect 17773 31291 17831 31297
rect 15304 31260 15332 31291
rect 15856 31260 15884 31291
rect 15304 31232 15884 31260
rect 15562 31152 15568 31204
rect 15620 31192 15626 31204
rect 16040 31192 16068 31291
rect 16758 31220 16764 31272
rect 16816 31260 16822 31272
rect 17604 31260 17632 31291
rect 17862 31288 17868 31340
rect 17920 31288 17926 31340
rect 17972 31337 18000 31368
rect 18506 31356 18512 31368
rect 18564 31356 18570 31408
rect 20990 31356 20996 31408
rect 21048 31405 21054 31408
rect 22094 31405 22100 31408
rect 21048 31396 21060 31405
rect 21048 31368 21093 31396
rect 21048 31359 21060 31368
rect 22088 31359 22100 31405
rect 22152 31396 22158 31408
rect 24504 31396 24532 31424
rect 22152 31368 22188 31396
rect 24136 31368 24532 31396
rect 21048 31356 21054 31359
rect 22094 31356 22100 31359
rect 22152 31356 22158 31368
rect 17957 31331 18015 31337
rect 17957 31297 17969 31331
rect 18003 31297 18015 31331
rect 17957 31291 18015 31297
rect 18141 31331 18199 31337
rect 18141 31297 18153 31331
rect 18187 31328 18199 31331
rect 18230 31328 18236 31340
rect 18187 31300 18236 31328
rect 18187 31297 18199 31300
rect 18141 31291 18199 31297
rect 18230 31288 18236 31300
rect 18288 31288 18294 31340
rect 21269 31331 21327 31337
rect 21269 31328 21281 31331
rect 19812 31300 21281 31328
rect 19812 31272 19840 31300
rect 21269 31297 21281 31300
rect 21315 31328 21327 31331
rect 21818 31328 21824 31340
rect 21315 31300 21824 31328
rect 21315 31297 21327 31300
rect 21269 31291 21327 31297
rect 21818 31288 21824 31300
rect 21876 31288 21882 31340
rect 23658 31288 23664 31340
rect 23716 31288 23722 31340
rect 24136 31337 24164 31368
rect 24121 31331 24179 31337
rect 24121 31297 24133 31331
rect 24167 31297 24179 31331
rect 24121 31291 24179 31297
rect 24302 31288 24308 31340
rect 24360 31328 24366 31340
rect 24670 31328 24676 31340
rect 24360 31300 24676 31328
rect 24360 31288 24366 31300
rect 24670 31288 24676 31300
rect 24728 31328 24734 31340
rect 24857 31331 24915 31337
rect 24857 31328 24869 31331
rect 24728 31300 24869 31328
rect 24728 31288 24734 31300
rect 24857 31297 24869 31300
rect 24903 31297 24915 31331
rect 24857 31291 24915 31297
rect 16816 31232 17632 31260
rect 18325 31263 18383 31269
rect 16816 31220 16822 31232
rect 18325 31229 18337 31263
rect 18371 31260 18383 31263
rect 18417 31263 18475 31269
rect 18417 31260 18429 31263
rect 18371 31232 18429 31260
rect 18371 31229 18383 31232
rect 18325 31223 18383 31229
rect 18417 31229 18429 31232
rect 18463 31229 18475 31263
rect 18417 31223 18475 31229
rect 19794 31220 19800 31272
rect 19852 31220 19858 31272
rect 23750 31220 23756 31272
rect 23808 31260 23814 31272
rect 24489 31263 24547 31269
rect 24489 31260 24501 31263
rect 23808 31232 24501 31260
rect 23808 31220 23814 31232
rect 24489 31229 24501 31232
rect 24535 31260 24547 31263
rect 24762 31260 24768 31272
rect 24535 31232 24768 31260
rect 24535 31229 24547 31232
rect 24489 31223 24547 31229
rect 24762 31220 24768 31232
rect 24820 31220 24826 31272
rect 15620 31164 20392 31192
rect 15620 31152 15626 31164
rect 20364 31136 20392 31164
rect 14292 31096 14872 31124
rect 15010 31084 15016 31136
rect 15068 31124 15074 31136
rect 15105 31127 15163 31133
rect 15105 31124 15117 31127
rect 15068 31096 15117 31124
rect 15068 31084 15074 31096
rect 15105 31093 15117 31096
rect 15151 31093 15163 31127
rect 15105 31087 15163 31093
rect 15654 31084 15660 31136
rect 15712 31084 15718 31136
rect 16022 31084 16028 31136
rect 16080 31084 16086 31136
rect 18966 31084 18972 31136
rect 19024 31124 19030 31136
rect 19061 31127 19119 31133
rect 19061 31124 19073 31127
rect 19024 31096 19073 31124
rect 19024 31084 19030 31096
rect 19061 31093 19073 31096
rect 19107 31093 19119 31127
rect 19061 31087 19119 31093
rect 20346 31084 20352 31136
rect 20404 31084 20410 31136
rect 25498 31084 25504 31136
rect 25556 31084 25562 31136
rect 1104 31034 34868 31056
rect 1104 30982 5170 31034
rect 5222 30982 5234 31034
rect 5286 30982 5298 31034
rect 5350 30982 5362 31034
rect 5414 30982 5426 31034
rect 5478 30982 13611 31034
rect 13663 30982 13675 31034
rect 13727 30982 13739 31034
rect 13791 30982 13803 31034
rect 13855 30982 13867 31034
rect 13919 30982 22052 31034
rect 22104 30982 22116 31034
rect 22168 30982 22180 31034
rect 22232 30982 22244 31034
rect 22296 30982 22308 31034
rect 22360 30982 30493 31034
rect 30545 30982 30557 31034
rect 30609 30982 30621 31034
rect 30673 30982 30685 31034
rect 30737 30982 30749 31034
rect 30801 30982 34868 31034
rect 1104 30960 34868 30982
rect 8110 30880 8116 30932
rect 8168 30920 8174 30932
rect 8205 30923 8263 30929
rect 8205 30920 8217 30923
rect 8168 30892 8217 30920
rect 8168 30880 8174 30892
rect 8205 30889 8217 30892
rect 8251 30889 8263 30923
rect 8205 30883 8263 30889
rect 10321 30923 10379 30929
rect 10321 30889 10333 30923
rect 10367 30920 10379 30923
rect 10502 30920 10508 30932
rect 10367 30892 10508 30920
rect 10367 30889 10379 30892
rect 10321 30883 10379 30889
rect 10502 30880 10508 30892
rect 10560 30880 10566 30932
rect 13817 30923 13875 30929
rect 13817 30889 13829 30923
rect 13863 30920 13875 30923
rect 15746 30920 15752 30932
rect 13863 30892 15752 30920
rect 13863 30889 13875 30892
rect 13817 30883 13875 30889
rect 15746 30880 15752 30892
rect 15804 30880 15810 30932
rect 16758 30920 16764 30932
rect 15856 30892 16764 30920
rect 15010 30812 15016 30864
rect 15068 30852 15074 30864
rect 15856 30852 15884 30892
rect 16758 30880 16764 30892
rect 16816 30880 16822 30932
rect 16942 30880 16948 30932
rect 17000 30920 17006 30932
rect 17221 30923 17279 30929
rect 17221 30920 17233 30923
rect 17000 30892 17233 30920
rect 17000 30880 17006 30892
rect 17221 30889 17233 30892
rect 17267 30889 17279 30923
rect 17221 30883 17279 30889
rect 17494 30880 17500 30932
rect 17552 30920 17558 30932
rect 17678 30920 17684 30932
rect 17552 30892 17684 30920
rect 17552 30880 17558 30892
rect 17678 30880 17684 30892
rect 17736 30880 17742 30932
rect 20717 30923 20775 30929
rect 18156 30892 20024 30920
rect 15068 30824 15884 30852
rect 16776 30852 16804 30880
rect 18156 30852 18184 30892
rect 16776 30824 18184 30852
rect 19996 30852 20024 30892
rect 20717 30889 20729 30923
rect 20763 30920 20775 30923
rect 20763 30892 22600 30920
rect 20763 30889 20775 30892
rect 20717 30883 20775 30889
rect 21542 30852 21548 30864
rect 19996 30824 21548 30852
rect 15068 30812 15074 30824
rect 12161 30787 12219 30793
rect 12161 30753 12173 30787
rect 12207 30784 12219 30787
rect 12710 30784 12716 30796
rect 12207 30756 12716 30784
rect 12207 30753 12219 30756
rect 12161 30747 12219 30753
rect 6825 30719 6883 30725
rect 6825 30685 6837 30719
rect 6871 30716 6883 30719
rect 8938 30716 8944 30728
rect 6871 30688 8944 30716
rect 6871 30685 6883 30688
rect 6825 30679 6883 30685
rect 8938 30676 8944 30688
rect 8996 30716 9002 30728
rect 12176 30716 12204 30747
rect 12710 30744 12716 30756
rect 12768 30744 12774 30796
rect 19061 30787 19119 30793
rect 19061 30753 19073 30787
rect 19107 30784 19119 30787
rect 19794 30784 19800 30796
rect 19107 30756 19800 30784
rect 19107 30753 19119 30756
rect 19061 30747 19119 30753
rect 19794 30744 19800 30756
rect 19852 30744 19858 30796
rect 8996 30688 12204 30716
rect 8996 30676 9002 30688
rect 12526 30676 12532 30728
rect 12584 30716 12590 30728
rect 12805 30719 12863 30725
rect 12805 30716 12817 30719
rect 12584 30688 12817 30716
rect 12584 30676 12590 30688
rect 12805 30685 12817 30688
rect 12851 30685 12863 30719
rect 12805 30679 12863 30685
rect 13354 30676 13360 30728
rect 13412 30676 13418 30728
rect 13446 30676 13452 30728
rect 13504 30716 13510 30728
rect 14277 30719 14335 30725
rect 14277 30716 14289 30719
rect 13504 30688 14289 30716
rect 13504 30676 13510 30688
rect 14277 30685 14289 30688
rect 14323 30685 14335 30719
rect 14277 30679 14335 30685
rect 14369 30719 14427 30725
rect 14369 30685 14381 30719
rect 14415 30685 14427 30719
rect 14369 30679 14427 30685
rect 6914 30608 6920 30660
rect 6972 30648 6978 30660
rect 7070 30651 7128 30657
rect 7070 30648 7082 30651
rect 6972 30620 7082 30648
rect 6972 30608 6978 30620
rect 7070 30617 7082 30620
rect 7116 30617 7128 30651
rect 7070 30611 7128 30617
rect 9208 30651 9266 30657
rect 9208 30617 9220 30651
rect 9254 30648 9266 30651
rect 9858 30648 9864 30660
rect 9254 30620 9864 30648
rect 9254 30617 9266 30620
rect 9208 30611 9266 30617
rect 9858 30608 9864 30620
rect 9916 30608 9922 30660
rect 10410 30608 10416 30660
rect 10468 30608 10474 30660
rect 13372 30648 13400 30676
rect 13541 30651 13599 30657
rect 13541 30648 13553 30651
rect 13372 30620 13553 30648
rect 13541 30617 13553 30620
rect 13587 30617 13599 30651
rect 13541 30611 13599 30617
rect 14182 30608 14188 30660
rect 14240 30648 14246 30660
rect 14384 30648 14412 30679
rect 14458 30676 14464 30728
rect 14516 30716 14522 30728
rect 14645 30719 14703 30725
rect 14645 30716 14657 30719
rect 14516 30688 14657 30716
rect 14516 30676 14522 30688
rect 14645 30685 14657 30688
rect 14691 30685 14703 30719
rect 14645 30679 14703 30685
rect 14734 30676 14740 30728
rect 14792 30676 14798 30728
rect 15102 30676 15108 30728
rect 15160 30676 15166 30728
rect 15378 30676 15384 30728
rect 15436 30716 15442 30728
rect 15841 30719 15899 30725
rect 15841 30716 15853 30719
rect 15436 30688 15853 30716
rect 15436 30676 15442 30688
rect 15841 30685 15853 30688
rect 15887 30685 15899 30719
rect 15841 30679 15899 30685
rect 17589 30719 17647 30725
rect 17589 30685 17601 30719
rect 17635 30716 17647 30719
rect 18230 30716 18236 30728
rect 17635 30688 18236 30716
rect 17635 30685 17647 30688
rect 17589 30679 17647 30685
rect 18230 30676 18236 30688
rect 18288 30676 18294 30728
rect 18805 30719 18863 30725
rect 18805 30685 18817 30719
rect 18851 30716 18863 30719
rect 18966 30716 18972 30728
rect 18851 30688 18972 30716
rect 18851 30685 18863 30688
rect 18805 30679 18863 30685
rect 18966 30676 18972 30688
rect 19024 30676 19030 30728
rect 19334 30676 19340 30728
rect 19392 30676 19398 30728
rect 19610 30676 19616 30728
rect 19668 30676 19674 30728
rect 19705 30719 19763 30725
rect 19705 30685 19717 30719
rect 19751 30716 19763 30719
rect 19886 30716 19892 30728
rect 19751 30688 19892 30716
rect 19751 30685 19763 30688
rect 19705 30679 19763 30685
rect 19886 30676 19892 30688
rect 19944 30676 19950 30728
rect 19996 30725 20024 30824
rect 21542 30812 21548 30824
rect 21600 30812 21606 30864
rect 21818 30812 21824 30864
rect 21876 30852 21882 30864
rect 22002 30852 22008 30864
rect 21876 30824 22008 30852
rect 21876 30812 21882 30824
rect 22002 30812 22008 30824
rect 22060 30852 22066 30864
rect 22097 30855 22155 30861
rect 22097 30852 22109 30855
rect 22060 30824 22109 30852
rect 22060 30812 22066 30824
rect 22097 30821 22109 30824
rect 22143 30821 22155 30855
rect 22572 30852 22600 30892
rect 22646 30880 22652 30932
rect 22704 30880 22710 30932
rect 23106 30880 23112 30932
rect 23164 30880 23170 30932
rect 23658 30880 23664 30932
rect 23716 30920 23722 30932
rect 24581 30923 24639 30929
rect 24581 30920 24593 30923
rect 23716 30892 24593 30920
rect 23716 30880 23722 30892
rect 24581 30889 24593 30892
rect 24627 30889 24639 30923
rect 24581 30883 24639 30889
rect 25498 30880 25504 30932
rect 25556 30880 25562 30932
rect 23124 30852 23152 30880
rect 22572 30824 23152 30852
rect 22097 30815 22155 30821
rect 23017 30787 23075 30793
rect 23017 30753 23029 30787
rect 23063 30784 23075 30787
rect 23474 30784 23480 30796
rect 23063 30756 23480 30784
rect 23063 30753 23075 30756
rect 23017 30747 23075 30753
rect 23474 30744 23480 30756
rect 23532 30744 23538 30796
rect 24949 30787 25007 30793
rect 24949 30753 24961 30787
rect 24995 30784 25007 30787
rect 25516 30784 25544 30880
rect 24995 30756 25544 30784
rect 24995 30753 25007 30756
rect 24949 30747 25007 30753
rect 19981 30719 20039 30725
rect 19981 30685 19993 30719
rect 20027 30685 20039 30719
rect 19981 30679 20039 30685
rect 20165 30719 20223 30725
rect 20165 30685 20177 30719
rect 20211 30685 20223 30719
rect 20165 30679 20223 30685
rect 14240 30620 14412 30648
rect 14240 30608 14246 30620
rect 14550 30608 14556 30660
rect 14608 30608 14614 30660
rect 14752 30648 14780 30676
rect 16086 30651 16144 30657
rect 16086 30648 16098 30651
rect 14660 30620 14780 30648
rect 15948 30620 16098 30648
rect 12066 30540 12072 30592
rect 12124 30580 12130 30592
rect 12253 30583 12311 30589
rect 12253 30580 12265 30583
rect 12124 30552 12265 30580
rect 12124 30540 12130 30552
rect 12253 30549 12265 30552
rect 12299 30549 12311 30583
rect 12253 30543 12311 30549
rect 14090 30540 14096 30592
rect 14148 30540 14154 30592
rect 14274 30540 14280 30592
rect 14332 30580 14338 30592
rect 14660 30580 14688 30620
rect 14332 30552 14688 30580
rect 14921 30583 14979 30589
rect 14332 30540 14338 30552
rect 14921 30549 14933 30583
rect 14967 30580 14979 30583
rect 15286 30580 15292 30592
rect 14967 30552 15292 30580
rect 14967 30549 14979 30552
rect 14921 30543 14979 30549
rect 15286 30540 15292 30552
rect 15344 30540 15350 30592
rect 15749 30583 15807 30589
rect 15749 30549 15761 30583
rect 15795 30580 15807 30583
rect 15948 30580 15976 30620
rect 16086 30617 16098 30620
rect 16132 30617 16144 30651
rect 16086 30611 16144 30617
rect 19518 30608 19524 30660
rect 19576 30608 19582 30660
rect 15795 30552 15976 30580
rect 15795 30549 15807 30552
rect 15749 30543 15807 30549
rect 17494 30540 17500 30592
rect 17552 30540 17558 30592
rect 19889 30583 19947 30589
rect 19889 30549 19901 30583
rect 19935 30580 19947 30583
rect 20180 30580 20208 30679
rect 20254 30676 20260 30728
rect 20312 30676 20318 30728
rect 20349 30719 20407 30725
rect 20349 30685 20361 30719
rect 20395 30716 20407 30719
rect 20438 30716 20444 30728
rect 20395 30688 20444 30716
rect 20395 30685 20407 30688
rect 20349 30679 20407 30685
rect 20438 30676 20444 30688
rect 20496 30676 20502 30728
rect 20533 30719 20591 30725
rect 20533 30685 20545 30719
rect 20579 30716 20591 30719
rect 21082 30716 21088 30728
rect 20579 30688 21088 30716
rect 20579 30685 20591 30688
rect 20533 30679 20591 30685
rect 21082 30676 21088 30688
rect 21140 30676 21146 30728
rect 22830 30676 22836 30728
rect 22888 30676 22894 30728
rect 23198 30676 23204 30728
rect 23256 30716 23262 30728
rect 23293 30719 23351 30725
rect 23293 30716 23305 30719
rect 23256 30688 23305 30716
rect 23256 30676 23262 30688
rect 23293 30685 23305 30688
rect 23339 30685 23351 30719
rect 23293 30679 23351 30685
rect 24765 30719 24823 30725
rect 24765 30685 24777 30719
rect 24811 30685 24823 30719
rect 24765 30679 24823 30685
rect 20809 30651 20867 30657
rect 20809 30617 20821 30651
rect 20855 30617 20867 30651
rect 22848 30648 22876 30676
rect 24780 30648 24808 30679
rect 22848 30620 24808 30648
rect 20809 30611 20867 30617
rect 19935 30552 20208 30580
rect 19935 30549 19947 30552
rect 19889 30543 19947 30549
rect 20530 30540 20536 30592
rect 20588 30580 20594 30592
rect 20824 30580 20852 30611
rect 20588 30552 20852 30580
rect 20588 30540 20594 30552
rect 23934 30540 23940 30592
rect 23992 30540 23998 30592
rect 1104 30490 35027 30512
rect 1104 30438 9390 30490
rect 9442 30438 9454 30490
rect 9506 30438 9518 30490
rect 9570 30438 9582 30490
rect 9634 30438 9646 30490
rect 9698 30438 17831 30490
rect 17883 30438 17895 30490
rect 17947 30438 17959 30490
rect 18011 30438 18023 30490
rect 18075 30438 18087 30490
rect 18139 30438 26272 30490
rect 26324 30438 26336 30490
rect 26388 30438 26400 30490
rect 26452 30438 26464 30490
rect 26516 30438 26528 30490
rect 26580 30438 34713 30490
rect 34765 30438 34777 30490
rect 34829 30438 34841 30490
rect 34893 30438 34905 30490
rect 34957 30438 34969 30490
rect 35021 30438 35027 30490
rect 1104 30416 35027 30438
rect 10226 30376 10232 30388
rect 9784 30348 10232 30376
rect 9493 30311 9551 30317
rect 9493 30277 9505 30311
rect 9539 30308 9551 30311
rect 9784 30308 9812 30348
rect 10226 30336 10232 30348
rect 10284 30336 10290 30388
rect 14642 30336 14648 30388
rect 14700 30336 14706 30388
rect 14829 30379 14887 30385
rect 14829 30345 14841 30379
rect 14875 30376 14887 30379
rect 15102 30376 15108 30388
rect 14875 30348 15108 30376
rect 14875 30345 14887 30348
rect 14829 30339 14887 30345
rect 15102 30336 15108 30348
rect 15160 30336 15166 30388
rect 16942 30336 16948 30388
rect 17000 30336 17006 30388
rect 17678 30336 17684 30388
rect 17736 30376 17742 30388
rect 19705 30379 19763 30385
rect 17736 30348 19288 30376
rect 17736 30336 17742 30348
rect 9539 30280 9812 30308
rect 9852 30311 9910 30317
rect 9539 30277 9551 30280
rect 9493 30271 9551 30277
rect 9852 30277 9864 30311
rect 9898 30308 9910 30311
rect 10042 30308 10048 30320
rect 9898 30280 10048 30308
rect 9898 30277 9910 30280
rect 9852 30271 9910 30277
rect 10042 30268 10048 30280
rect 10100 30268 10106 30320
rect 12152 30311 12210 30317
rect 12152 30277 12164 30311
rect 12198 30308 12210 30311
rect 14090 30308 14096 30320
rect 12198 30280 14096 30308
rect 12198 30277 12210 30280
rect 12152 30271 12210 30277
rect 14090 30268 14096 30280
rect 14148 30268 14154 30320
rect 14660 30308 14688 30336
rect 15930 30308 15936 30320
rect 14660 30280 14964 30308
rect 6546 30200 6552 30252
rect 6604 30200 6610 30252
rect 8110 30200 8116 30252
rect 8168 30200 8174 30252
rect 8938 30200 8944 30252
rect 8996 30240 9002 30252
rect 9309 30243 9367 30249
rect 8996 30212 9260 30240
rect 8996 30200 9002 30212
rect 6914 30172 6920 30184
rect 6748 30144 6920 30172
rect 6748 30113 6776 30144
rect 6914 30132 6920 30144
rect 6972 30132 6978 30184
rect 9125 30175 9183 30181
rect 9125 30141 9137 30175
rect 9171 30141 9183 30175
rect 9232 30172 9260 30212
rect 9309 30209 9321 30243
rect 9355 30240 9367 30243
rect 9398 30240 9404 30252
rect 9355 30212 9404 30240
rect 9355 30209 9367 30212
rect 9309 30203 9367 30209
rect 9398 30200 9404 30212
rect 9456 30200 9462 30252
rect 11514 30200 11520 30252
rect 11572 30200 11578 30252
rect 11885 30243 11943 30249
rect 11885 30209 11897 30243
rect 11931 30240 11943 30243
rect 12710 30240 12716 30252
rect 11931 30212 12716 30240
rect 11931 30209 11943 30212
rect 11885 30203 11943 30209
rect 12710 30200 12716 30212
rect 12768 30200 12774 30252
rect 13725 30243 13783 30249
rect 13725 30209 13737 30243
rect 13771 30240 13783 30243
rect 13771 30212 14872 30240
rect 13771 30209 13783 30212
rect 13725 30203 13783 30209
rect 9585 30175 9643 30181
rect 9585 30172 9597 30175
rect 9232 30144 9597 30172
rect 9125 30135 9183 30141
rect 9585 30141 9597 30144
rect 9631 30141 9643 30175
rect 9585 30135 9643 30141
rect 6733 30107 6791 30113
rect 6733 30073 6745 30107
rect 6779 30073 6791 30107
rect 6733 30067 6791 30073
rect 7926 29996 7932 30048
rect 7984 29996 7990 30048
rect 9140 30036 9168 30135
rect 13998 30132 14004 30184
rect 14056 30132 14062 30184
rect 14093 30175 14151 30181
rect 14093 30141 14105 30175
rect 14139 30141 14151 30175
rect 14093 30135 14151 30141
rect 11146 30104 11152 30116
rect 10888 30076 11152 30104
rect 10888 30036 10916 30076
rect 11146 30064 11152 30076
rect 11204 30064 11210 30116
rect 13541 30107 13599 30113
rect 13541 30073 13553 30107
rect 13587 30104 13599 30107
rect 14108 30104 14136 30135
rect 14550 30132 14556 30184
rect 14608 30132 14614 30184
rect 13587 30076 14136 30104
rect 13587 30073 13599 30076
rect 13541 30067 13599 30073
rect 9140 30008 10916 30036
rect 10962 29996 10968 30048
rect 11020 29996 11026 30048
rect 11698 29996 11704 30048
rect 11756 29996 11762 30048
rect 13262 29996 13268 30048
rect 13320 29996 13326 30048
rect 13909 30039 13967 30045
rect 13909 30005 13921 30039
rect 13955 30036 13967 30039
rect 13998 30036 14004 30048
rect 13955 30008 14004 30036
rect 13955 30005 13967 30008
rect 13909 29999 13967 30005
rect 13998 29996 14004 30008
rect 14056 30036 14062 30048
rect 14568 30036 14596 30132
rect 14844 30104 14872 30212
rect 14936 30172 14964 30280
rect 15120 30280 15936 30308
rect 15120 30249 15148 30280
rect 15930 30268 15936 30280
rect 15988 30268 15994 30320
rect 16960 30308 16988 30336
rect 18340 30317 18368 30348
rect 18233 30311 18291 30317
rect 18233 30308 18245 30311
rect 16960 30280 17356 30308
rect 15105 30243 15163 30249
rect 15105 30209 15117 30243
rect 15151 30209 15163 30243
rect 15105 30203 15163 30209
rect 15197 30243 15255 30249
rect 15197 30209 15209 30243
rect 15243 30209 15255 30243
rect 15197 30203 15255 30209
rect 15289 30243 15347 30249
rect 15289 30209 15301 30243
rect 15335 30209 15347 30243
rect 15289 30203 15347 30209
rect 15212 30172 15240 30203
rect 14936 30144 15240 30172
rect 15304 30172 15332 30203
rect 15470 30200 15476 30252
rect 15528 30200 15534 30252
rect 15562 30200 15568 30252
rect 15620 30200 15626 30252
rect 16758 30200 16764 30252
rect 16816 30200 16822 30252
rect 16942 30200 16948 30252
rect 17000 30200 17006 30252
rect 17034 30200 17040 30252
rect 17092 30200 17098 30252
rect 17218 30200 17224 30252
rect 17276 30200 17282 30252
rect 17328 30249 17356 30280
rect 17512 30280 18245 30308
rect 17512 30252 17540 30280
rect 18233 30277 18245 30280
rect 18279 30277 18291 30311
rect 18233 30271 18291 30277
rect 18325 30311 18383 30317
rect 18325 30277 18337 30311
rect 18371 30277 18383 30311
rect 18325 30271 18383 30277
rect 18616 30280 19196 30308
rect 17313 30243 17371 30249
rect 17313 30209 17325 30243
rect 17359 30209 17371 30243
rect 17313 30203 17371 30209
rect 17405 30243 17463 30249
rect 17405 30209 17417 30243
rect 17451 30240 17463 30243
rect 17494 30240 17500 30252
rect 17451 30212 17500 30240
rect 17451 30209 17463 30212
rect 17405 30203 17463 30209
rect 17494 30200 17500 30212
rect 17552 30200 17558 30252
rect 17589 30243 17647 30249
rect 17589 30209 17601 30243
rect 17635 30209 17647 30243
rect 17589 30203 17647 30209
rect 17773 30243 17831 30249
rect 17773 30209 17785 30243
rect 17819 30240 17831 30243
rect 17957 30243 18015 30249
rect 17957 30240 17969 30243
rect 17819 30212 17969 30240
rect 17819 30209 17831 30212
rect 17773 30203 17831 30209
rect 17957 30209 17969 30212
rect 18003 30209 18015 30243
rect 17957 30203 18015 30209
rect 18105 30243 18163 30249
rect 18105 30209 18117 30243
rect 18151 30240 18163 30243
rect 18463 30243 18521 30249
rect 18151 30209 18184 30240
rect 18105 30203 18184 30209
rect 18463 30209 18475 30243
rect 18509 30240 18521 30243
rect 18616 30240 18644 30280
rect 19168 30252 19196 30280
rect 18509 30212 18644 30240
rect 18509 30209 18521 30212
rect 18463 30203 18521 30209
rect 16850 30172 16856 30184
rect 15304 30144 16856 30172
rect 16850 30132 16856 30144
rect 16908 30132 16914 30184
rect 16022 30104 16028 30116
rect 14844 30076 16028 30104
rect 16022 30064 16028 30076
rect 16080 30064 16086 30116
rect 16574 30064 16580 30116
rect 16632 30104 16638 30116
rect 17236 30104 17264 30200
rect 17604 30172 17632 30203
rect 18156 30172 18184 30203
rect 18690 30200 18696 30252
rect 18748 30200 18754 30252
rect 18874 30200 18880 30252
rect 18932 30200 18938 30252
rect 18969 30243 19027 30249
rect 18969 30209 18981 30243
rect 19015 30209 19027 30243
rect 18969 30203 19027 30209
rect 18984 30172 19012 30203
rect 19150 30200 19156 30252
rect 19208 30200 19214 30252
rect 19260 30249 19288 30348
rect 19705 30345 19717 30379
rect 19751 30376 19763 30379
rect 20254 30376 20260 30388
rect 19751 30348 20260 30376
rect 19751 30345 19763 30348
rect 19705 30339 19763 30345
rect 20254 30336 20260 30348
rect 20312 30336 20318 30388
rect 20438 30336 20444 30388
rect 20496 30376 20502 30388
rect 20533 30379 20591 30385
rect 20533 30376 20545 30379
rect 20496 30348 20545 30376
rect 20496 30336 20502 30348
rect 20533 30345 20545 30348
rect 20579 30345 20591 30379
rect 20533 30339 20591 30345
rect 24670 30336 24676 30388
rect 24728 30336 24734 30388
rect 19886 30268 19892 30320
rect 19944 30308 19950 30320
rect 20456 30308 20484 30336
rect 19944 30280 20484 30308
rect 19944 30268 19950 30280
rect 21726 30268 21732 30320
rect 21784 30308 21790 30320
rect 22097 30311 22155 30317
rect 22097 30308 22109 30311
rect 21784 30280 22109 30308
rect 21784 30268 21790 30280
rect 22097 30277 22109 30280
rect 22143 30308 22155 30311
rect 23198 30308 23204 30320
rect 22143 30280 23204 30308
rect 22143 30277 22155 30280
rect 22097 30271 22155 30277
rect 23198 30268 23204 30280
rect 23256 30268 23262 30320
rect 19245 30243 19303 30249
rect 19245 30209 19257 30243
rect 19291 30209 19303 30243
rect 19245 30203 19303 30209
rect 19426 30200 19432 30252
rect 19484 30240 19490 30252
rect 19521 30243 19579 30249
rect 19521 30240 19533 30243
rect 19484 30212 19533 30240
rect 19484 30200 19490 30212
rect 19521 30209 19533 30212
rect 19567 30209 19579 30243
rect 19521 30203 19579 30209
rect 19981 30243 20039 30249
rect 19981 30209 19993 30243
rect 20027 30209 20039 30243
rect 19981 30203 20039 30209
rect 20073 30243 20131 30249
rect 20073 30209 20085 30243
rect 20119 30240 20131 30243
rect 20162 30240 20168 30252
rect 20119 30212 20168 30240
rect 20119 30209 20131 30212
rect 20073 30203 20131 30209
rect 17604 30144 18184 30172
rect 16632 30076 17264 30104
rect 16632 30064 16638 30076
rect 14056 30008 14596 30036
rect 14056 29996 14062 30008
rect 14734 29996 14740 30048
rect 14792 29996 14798 30048
rect 15746 29996 15752 30048
rect 15804 29996 15810 30048
rect 16945 30039 17003 30045
rect 16945 30005 16957 30039
rect 16991 30036 17003 30039
rect 17126 30036 17132 30048
rect 16991 30008 17132 30036
rect 16991 30005 17003 30008
rect 16945 29999 17003 30005
rect 17126 29996 17132 30008
rect 17184 29996 17190 30048
rect 18156 30036 18184 30144
rect 18616 30144 19012 30172
rect 19337 30175 19395 30181
rect 18616 30113 18644 30144
rect 19337 30141 19349 30175
rect 19383 30172 19395 30175
rect 19886 30172 19892 30184
rect 19383 30144 19892 30172
rect 19383 30141 19395 30144
rect 19337 30135 19395 30141
rect 19536 30116 19564 30144
rect 19886 30132 19892 30144
rect 19944 30132 19950 30184
rect 19996 30172 20024 30203
rect 20162 30200 20168 30212
rect 20220 30200 20226 30252
rect 20257 30243 20315 30249
rect 20257 30209 20269 30243
rect 20303 30240 20315 30243
rect 20346 30240 20352 30252
rect 20303 30212 20352 30240
rect 20303 30209 20315 30212
rect 20257 30203 20315 30209
rect 20346 30200 20352 30212
rect 20404 30200 20410 30252
rect 20625 30243 20683 30249
rect 20625 30209 20637 30243
rect 20671 30240 20683 30243
rect 20990 30240 20996 30252
rect 20671 30212 20996 30240
rect 20671 30209 20683 30212
rect 20625 30203 20683 30209
rect 20990 30200 20996 30212
rect 21048 30200 21054 30252
rect 21634 30200 21640 30252
rect 21692 30240 21698 30252
rect 21821 30243 21879 30249
rect 21821 30240 21833 30243
rect 21692 30212 21833 30240
rect 21692 30200 21698 30212
rect 21821 30209 21833 30212
rect 21867 30209 21879 30243
rect 21821 30203 21879 30209
rect 22002 30200 22008 30252
rect 22060 30240 22066 30252
rect 23293 30243 23351 30249
rect 23293 30240 23305 30243
rect 22060 30212 23305 30240
rect 22060 30200 22066 30212
rect 23293 30209 23305 30212
rect 23339 30209 23351 30243
rect 23293 30203 23351 30209
rect 23560 30243 23618 30249
rect 23560 30209 23572 30243
rect 23606 30240 23618 30243
rect 23842 30240 23848 30252
rect 23606 30212 23848 30240
rect 23606 30209 23618 30212
rect 23560 30203 23618 30209
rect 23842 30200 23848 30212
rect 23900 30200 23906 30252
rect 19996 30144 20576 30172
rect 18601 30107 18659 30113
rect 18601 30073 18613 30107
rect 18647 30073 18659 30107
rect 18601 30067 18659 30073
rect 18782 30064 18788 30116
rect 18840 30064 18846 30116
rect 18966 30064 18972 30116
rect 19024 30104 19030 30116
rect 19024 30076 19380 30104
rect 19024 30064 19030 30076
rect 18800 30036 18828 30064
rect 19352 30048 19380 30076
rect 19518 30064 19524 30116
rect 19576 30064 19582 30116
rect 18156 30008 18828 30036
rect 18874 29996 18880 30048
rect 18932 29996 18938 30048
rect 19334 29996 19340 30048
rect 19392 30036 19398 30048
rect 19996 30036 20024 30144
rect 20548 30048 20576 30144
rect 20714 30132 20720 30184
rect 20772 30172 20778 30184
rect 20772 30144 22876 30172
rect 20772 30132 20778 30144
rect 21266 30064 21272 30116
rect 21324 30104 21330 30116
rect 22373 30107 22431 30113
rect 22373 30104 22385 30107
rect 21324 30076 22385 30104
rect 21324 30064 21330 30076
rect 22373 30073 22385 30076
rect 22419 30073 22431 30107
rect 22373 30067 22431 30073
rect 19392 30008 20024 30036
rect 19392 29996 19398 30008
rect 20254 29996 20260 30048
rect 20312 29996 20318 30048
rect 20530 29996 20536 30048
rect 20588 29996 20594 30048
rect 21818 29996 21824 30048
rect 21876 30036 21882 30048
rect 22005 30039 22063 30045
rect 22005 30036 22017 30039
rect 21876 30008 22017 30036
rect 21876 29996 21882 30008
rect 22005 30005 22017 30008
rect 22051 30005 22063 30039
rect 22005 29999 22063 30005
rect 22557 30039 22615 30045
rect 22557 30005 22569 30039
rect 22603 30036 22615 30039
rect 22646 30036 22652 30048
rect 22603 30008 22652 30036
rect 22603 30005 22615 30008
rect 22557 29999 22615 30005
rect 22646 29996 22652 30008
rect 22704 29996 22710 30048
rect 22848 30036 22876 30144
rect 23566 30036 23572 30048
rect 22848 30008 23572 30036
rect 23566 29996 23572 30008
rect 23624 29996 23630 30048
rect 1104 29946 34868 29968
rect 1104 29894 5170 29946
rect 5222 29894 5234 29946
rect 5286 29894 5298 29946
rect 5350 29894 5362 29946
rect 5414 29894 5426 29946
rect 5478 29894 13611 29946
rect 13663 29894 13675 29946
rect 13727 29894 13739 29946
rect 13791 29894 13803 29946
rect 13855 29894 13867 29946
rect 13919 29894 22052 29946
rect 22104 29894 22116 29946
rect 22168 29894 22180 29946
rect 22232 29894 22244 29946
rect 22296 29894 22308 29946
rect 22360 29894 30493 29946
rect 30545 29894 30557 29946
rect 30609 29894 30621 29946
rect 30673 29894 30685 29946
rect 30737 29894 30749 29946
rect 30801 29894 34868 29946
rect 1104 29872 34868 29894
rect 6273 29835 6331 29841
rect 6273 29801 6285 29835
rect 6319 29832 6331 29835
rect 6546 29832 6552 29844
rect 6319 29804 6552 29832
rect 6319 29801 6331 29804
rect 6273 29795 6331 29801
rect 6546 29792 6552 29804
rect 6604 29792 6610 29844
rect 9858 29792 9864 29844
rect 9916 29832 9922 29844
rect 10505 29835 10563 29841
rect 10505 29832 10517 29835
rect 9916 29804 10517 29832
rect 9916 29792 9922 29804
rect 10505 29801 10517 29804
rect 10551 29801 10563 29835
rect 11974 29832 11980 29844
rect 10505 29795 10563 29801
rect 11072 29804 11980 29832
rect 10226 29724 10232 29776
rect 10284 29764 10290 29776
rect 10962 29764 10968 29776
rect 10284 29736 10968 29764
rect 10284 29724 10290 29736
rect 10962 29724 10968 29736
rect 11020 29724 11026 29776
rect 5905 29699 5963 29705
rect 5905 29665 5917 29699
rect 5951 29696 5963 29699
rect 5994 29696 6000 29708
rect 5951 29668 6000 29696
rect 5951 29665 5963 29668
rect 5905 29659 5963 29665
rect 5994 29656 6000 29668
rect 6052 29656 6058 29708
rect 8846 29656 8852 29708
rect 8904 29696 8910 29708
rect 9398 29696 9404 29708
rect 8904 29668 9404 29696
rect 8904 29656 8910 29668
rect 9398 29656 9404 29668
rect 9456 29696 9462 29708
rect 11072 29696 11100 29804
rect 11974 29792 11980 29804
rect 12032 29792 12038 29844
rect 12710 29792 12716 29844
rect 12768 29832 12774 29844
rect 15378 29832 15384 29844
rect 12768 29804 15384 29832
rect 12768 29792 12774 29804
rect 14108 29705 14136 29804
rect 15378 29792 15384 29804
rect 15436 29792 15442 29844
rect 15473 29835 15531 29841
rect 15473 29801 15485 29835
rect 15519 29832 15531 29835
rect 15562 29832 15568 29844
rect 15519 29804 15568 29832
rect 15519 29801 15531 29804
rect 15473 29795 15531 29801
rect 15562 29792 15568 29804
rect 15620 29792 15626 29844
rect 16117 29835 16175 29841
rect 16117 29801 16129 29835
rect 16163 29832 16175 29835
rect 16666 29832 16672 29844
rect 16163 29804 16672 29832
rect 16163 29801 16175 29804
rect 16117 29795 16175 29801
rect 16666 29792 16672 29804
rect 16724 29792 16730 29844
rect 16776 29804 18368 29832
rect 9456 29668 11100 29696
rect 14093 29699 14151 29705
rect 9456 29656 9462 29668
rect 6086 29588 6092 29640
rect 6144 29588 6150 29640
rect 7374 29588 7380 29640
rect 7432 29588 7438 29640
rect 7644 29631 7702 29637
rect 7644 29597 7656 29631
rect 7690 29628 7702 29631
rect 7926 29628 7932 29640
rect 7690 29600 7932 29628
rect 7690 29597 7702 29600
rect 7644 29591 7702 29597
rect 7926 29588 7932 29600
rect 7984 29588 7990 29640
rect 9306 29588 9312 29640
rect 9364 29628 9370 29640
rect 10244 29637 10272 29668
rect 14093 29665 14105 29699
rect 14139 29665 14151 29699
rect 15470 29696 15476 29708
rect 14093 29659 14151 29665
rect 15212 29668 15476 29696
rect 9493 29631 9551 29637
rect 9493 29628 9505 29631
rect 9364 29600 9505 29628
rect 9364 29588 9370 29600
rect 9493 29597 9505 29600
rect 9539 29597 9551 29631
rect 9493 29591 9551 29597
rect 10137 29631 10195 29637
rect 10137 29597 10149 29631
rect 10183 29597 10195 29631
rect 10137 29591 10195 29597
rect 10229 29631 10287 29637
rect 10229 29597 10241 29631
rect 10275 29597 10287 29631
rect 10229 29591 10287 29597
rect 10413 29631 10471 29637
rect 10413 29597 10425 29631
rect 10459 29628 10471 29631
rect 10689 29631 10747 29637
rect 10689 29628 10701 29631
rect 10459 29600 10701 29628
rect 10459 29597 10471 29600
rect 10413 29591 10471 29597
rect 10689 29597 10701 29600
rect 10735 29597 10747 29631
rect 10689 29591 10747 29597
rect 11905 29631 11963 29637
rect 11905 29597 11917 29631
rect 11951 29628 11963 29631
rect 12066 29628 12072 29640
rect 11951 29600 12072 29628
rect 11951 29597 11963 29600
rect 11905 29591 11963 29597
rect 8478 29452 8484 29504
rect 8536 29492 8542 29504
rect 8757 29495 8815 29501
rect 8757 29492 8769 29495
rect 8536 29464 8769 29492
rect 8536 29452 8542 29464
rect 8757 29461 8769 29464
rect 8803 29461 8815 29495
rect 8757 29455 8815 29461
rect 8938 29452 8944 29504
rect 8996 29452 9002 29504
rect 10152 29492 10180 29591
rect 12066 29588 12072 29600
rect 12124 29588 12130 29640
rect 12158 29588 12164 29640
rect 12216 29588 12222 29640
rect 12253 29631 12311 29637
rect 12253 29597 12265 29631
rect 12299 29597 12311 29631
rect 12253 29591 12311 29597
rect 13081 29631 13139 29637
rect 13081 29597 13093 29631
rect 13127 29628 13139 29631
rect 13354 29628 13360 29640
rect 13127 29600 13360 29628
rect 13127 29597 13139 29600
rect 13081 29591 13139 29597
rect 10686 29492 10692 29504
rect 10152 29464 10692 29492
rect 10686 29452 10692 29464
rect 10744 29452 10750 29504
rect 10778 29452 10784 29504
rect 10836 29492 10842 29504
rect 12268 29492 12296 29591
rect 13354 29588 13360 29600
rect 13412 29588 13418 29640
rect 14360 29631 14418 29637
rect 14360 29597 14372 29631
rect 14406 29628 14418 29631
rect 14734 29628 14740 29640
rect 14406 29600 14740 29628
rect 14406 29597 14418 29600
rect 14360 29591 14418 29597
rect 14734 29588 14740 29600
rect 14792 29588 14798 29640
rect 12434 29520 12440 29572
rect 12492 29560 12498 29572
rect 13449 29563 13507 29569
rect 13449 29560 13461 29563
rect 12492 29532 13461 29560
rect 12492 29520 12498 29532
rect 13449 29529 13461 29532
rect 13495 29560 13507 29563
rect 15212 29560 15240 29668
rect 15470 29656 15476 29668
rect 15528 29696 15534 29708
rect 16776 29696 16804 29804
rect 18340 29764 18368 29804
rect 18414 29792 18420 29844
rect 18472 29792 18478 29844
rect 18969 29835 19027 29841
rect 18969 29801 18981 29835
rect 19015 29832 19027 29835
rect 19150 29832 19156 29844
rect 19015 29804 19156 29832
rect 19015 29801 19027 29804
rect 18969 29795 19027 29801
rect 19150 29792 19156 29804
rect 19208 29792 19214 29844
rect 19245 29835 19303 29841
rect 19245 29801 19257 29835
rect 19291 29832 19303 29835
rect 19334 29832 19340 29844
rect 19291 29804 19340 29832
rect 19291 29801 19303 29804
rect 19245 29795 19303 29801
rect 19334 29792 19340 29804
rect 19392 29792 19398 29844
rect 19429 29835 19487 29841
rect 19429 29801 19441 29835
rect 19475 29801 19487 29835
rect 19429 29795 19487 29801
rect 18506 29764 18512 29776
rect 18340 29736 18512 29764
rect 18506 29724 18512 29736
rect 18564 29724 18570 29776
rect 19058 29724 19064 29776
rect 19116 29764 19122 29776
rect 19444 29764 19472 29795
rect 19886 29792 19892 29844
rect 19944 29832 19950 29844
rect 20717 29835 20775 29841
rect 20717 29832 20729 29835
rect 19944 29804 20729 29832
rect 19944 29792 19950 29804
rect 20717 29801 20729 29804
rect 20763 29801 20775 29835
rect 20717 29795 20775 29801
rect 21634 29792 21640 29844
rect 21692 29832 21698 29844
rect 23385 29835 23443 29841
rect 23385 29832 23397 29835
rect 21692 29804 23397 29832
rect 21692 29792 21698 29804
rect 23385 29801 23397 29804
rect 23431 29801 23443 29835
rect 23385 29795 23443 29801
rect 23842 29792 23848 29844
rect 23900 29792 23906 29844
rect 19116 29736 19472 29764
rect 19116 29724 19122 29736
rect 19978 29724 19984 29776
rect 20036 29764 20042 29776
rect 20346 29764 20352 29776
rect 20036 29736 20352 29764
rect 20036 29724 20042 29736
rect 20346 29724 20352 29736
rect 20404 29724 20410 29776
rect 21726 29724 21732 29776
rect 21784 29724 21790 29776
rect 15528 29668 16804 29696
rect 18064 29668 22048 29696
rect 15528 29656 15534 29668
rect 15286 29588 15292 29640
rect 15344 29628 15350 29640
rect 15565 29631 15623 29637
rect 15565 29628 15577 29631
rect 15344 29600 15577 29628
rect 15344 29588 15350 29600
rect 15565 29597 15577 29600
rect 15611 29597 15623 29631
rect 15565 29591 15623 29597
rect 15654 29588 15660 29640
rect 15712 29628 15718 29640
rect 15749 29631 15807 29637
rect 15749 29628 15761 29631
rect 15712 29600 15761 29628
rect 15712 29588 15718 29600
rect 15749 29597 15761 29600
rect 15795 29597 15807 29631
rect 15749 29591 15807 29597
rect 15838 29588 15844 29640
rect 15896 29588 15902 29640
rect 15933 29631 15991 29637
rect 15933 29597 15945 29631
rect 15979 29597 15991 29631
rect 18064 29628 18092 29668
rect 15933 29591 15991 29597
rect 17972 29600 18092 29628
rect 13495 29532 15240 29560
rect 15948 29560 15976 29591
rect 17862 29560 17868 29572
rect 15948 29532 17868 29560
rect 13495 29529 13507 29532
rect 13449 29523 13507 29529
rect 10836 29464 12296 29492
rect 10836 29452 10842 29464
rect 12342 29452 12348 29504
rect 12400 29492 12406 29504
rect 12897 29495 12955 29501
rect 12897 29492 12909 29495
rect 12400 29464 12909 29492
rect 12400 29452 12406 29464
rect 12897 29461 12909 29464
rect 12943 29461 12955 29495
rect 12897 29455 12955 29461
rect 14458 29452 14464 29504
rect 14516 29492 14522 29504
rect 15948 29492 15976 29532
rect 17862 29520 17868 29532
rect 17920 29520 17926 29572
rect 17972 29569 18000 29600
rect 18414 29588 18420 29640
rect 18472 29628 18478 29640
rect 18509 29631 18567 29637
rect 18509 29628 18521 29631
rect 18472 29600 18521 29628
rect 18472 29588 18478 29600
rect 18509 29597 18521 29600
rect 18555 29628 18567 29631
rect 18598 29628 18604 29640
rect 18555 29600 18604 29628
rect 18555 29597 18567 29600
rect 18509 29591 18567 29597
rect 18598 29588 18604 29600
rect 18656 29588 18662 29640
rect 18693 29631 18751 29637
rect 18693 29597 18705 29631
rect 18739 29628 18751 29631
rect 18966 29628 18972 29640
rect 18739 29600 18972 29628
rect 18739 29597 18751 29600
rect 18693 29591 18751 29597
rect 18966 29588 18972 29600
rect 19024 29588 19030 29640
rect 19058 29588 19064 29640
rect 19116 29588 19122 29640
rect 19334 29588 19340 29640
rect 19392 29588 19398 29640
rect 20438 29588 20444 29640
rect 20496 29588 20502 29640
rect 20622 29588 20628 29640
rect 20680 29588 20686 29640
rect 20714 29588 20720 29640
rect 20772 29588 20778 29640
rect 20806 29588 20812 29640
rect 20864 29628 20870 29640
rect 20901 29631 20959 29637
rect 20901 29628 20913 29631
rect 20864 29600 20913 29628
rect 20864 29588 20870 29600
rect 20901 29597 20913 29600
rect 20947 29597 20959 29631
rect 20901 29591 20959 29597
rect 21085 29631 21143 29637
rect 21085 29597 21097 29631
rect 21131 29597 21143 29631
rect 21085 29591 21143 29597
rect 17957 29563 18015 29569
rect 17957 29529 17969 29563
rect 18003 29529 18015 29563
rect 17957 29523 18015 29529
rect 18046 29520 18052 29572
rect 18104 29520 18110 29572
rect 18138 29520 18144 29572
rect 18196 29560 18202 29572
rect 18233 29563 18291 29569
rect 18233 29560 18245 29563
rect 18196 29532 18245 29560
rect 18196 29520 18202 29532
rect 18233 29529 18245 29532
rect 18279 29529 18291 29563
rect 19352 29560 19380 29588
rect 19613 29563 19671 29569
rect 19352 29532 19463 29560
rect 18233 29523 18291 29529
rect 14516 29464 15976 29492
rect 16669 29495 16727 29501
rect 14516 29452 14522 29464
rect 16669 29461 16681 29495
rect 16715 29492 16727 29495
rect 18322 29492 18328 29504
rect 16715 29464 18328 29492
rect 16715 29461 16727 29464
rect 16669 29455 16727 29461
rect 18322 29452 18328 29464
rect 18380 29452 18386 29504
rect 18598 29452 18604 29504
rect 18656 29452 18662 29504
rect 18690 29452 18696 29504
rect 18748 29492 18754 29504
rect 19150 29492 19156 29504
rect 18748 29464 19156 29492
rect 18748 29452 18754 29464
rect 19150 29452 19156 29464
rect 19208 29452 19214 29504
rect 19435 29501 19463 29532
rect 19613 29529 19625 29563
rect 19659 29560 19671 29563
rect 19702 29560 19708 29572
rect 19659 29532 19708 29560
rect 19659 29529 19671 29532
rect 19613 29523 19671 29529
rect 19702 29520 19708 29532
rect 19760 29520 19766 29572
rect 20732 29560 20760 29588
rect 21100 29560 21128 29591
rect 21266 29588 21272 29640
rect 21324 29628 21330 29640
rect 21361 29631 21419 29637
rect 21361 29628 21373 29631
rect 21324 29600 21373 29628
rect 21324 29588 21330 29600
rect 21361 29597 21373 29600
rect 21407 29597 21419 29631
rect 21361 29591 21419 29597
rect 21818 29588 21824 29640
rect 21876 29588 21882 29640
rect 21910 29588 21916 29640
rect 21968 29588 21974 29640
rect 22020 29628 22048 29668
rect 23492 29668 29040 29696
rect 23492 29628 23520 29668
rect 29012 29640 29040 29668
rect 22020 29600 23520 29628
rect 23566 29588 23572 29640
rect 23624 29588 23630 29640
rect 23753 29631 23811 29637
rect 23753 29597 23765 29631
rect 23799 29628 23811 29631
rect 23934 29628 23940 29640
rect 23799 29600 23940 29628
rect 23799 29597 23811 29600
rect 23753 29591 23811 29597
rect 23934 29588 23940 29600
rect 23992 29588 23998 29640
rect 24026 29588 24032 29640
rect 24084 29588 24090 29640
rect 28994 29588 29000 29640
rect 29052 29588 29058 29640
rect 20732 29532 21128 29560
rect 21836 29560 21864 29588
rect 22158 29563 22216 29569
rect 22158 29560 22170 29563
rect 21836 29532 22170 29560
rect 22158 29529 22170 29532
rect 22204 29529 22216 29563
rect 22158 29523 22216 29529
rect 19403 29495 19463 29501
rect 19403 29461 19415 29495
rect 19449 29464 19463 29495
rect 19449 29461 19461 29464
rect 19403 29455 19461 29461
rect 19886 29452 19892 29504
rect 19944 29452 19950 29504
rect 21174 29452 21180 29504
rect 21232 29492 21238 29504
rect 21269 29495 21327 29501
rect 21269 29492 21281 29495
rect 21232 29464 21281 29492
rect 21232 29452 21238 29464
rect 21269 29461 21281 29464
rect 21315 29461 21327 29495
rect 21269 29455 21327 29461
rect 21821 29495 21879 29501
rect 21821 29461 21833 29495
rect 21867 29492 21879 29495
rect 22738 29492 22744 29504
rect 21867 29464 22744 29492
rect 21867 29461 21879 29464
rect 21821 29455 21879 29461
rect 22738 29452 22744 29464
rect 22796 29452 22802 29504
rect 23290 29452 23296 29504
rect 23348 29452 23354 29504
rect 1104 29402 35027 29424
rect 1104 29350 9390 29402
rect 9442 29350 9454 29402
rect 9506 29350 9518 29402
rect 9570 29350 9582 29402
rect 9634 29350 9646 29402
rect 9698 29350 17831 29402
rect 17883 29350 17895 29402
rect 17947 29350 17959 29402
rect 18011 29350 18023 29402
rect 18075 29350 18087 29402
rect 18139 29350 26272 29402
rect 26324 29350 26336 29402
rect 26388 29350 26400 29402
rect 26452 29350 26464 29402
rect 26516 29350 26528 29402
rect 26580 29350 34713 29402
rect 34765 29350 34777 29402
rect 34829 29350 34841 29402
rect 34893 29350 34905 29402
rect 34957 29350 34969 29402
rect 35021 29350 35027 29402
rect 1104 29328 35027 29350
rect 1581 29291 1639 29297
rect 1581 29257 1593 29291
rect 1627 29288 1639 29291
rect 6086 29288 6092 29300
rect 1627 29260 6092 29288
rect 1627 29257 1639 29260
rect 1581 29251 1639 29257
rect 6086 29248 6092 29260
rect 6144 29248 6150 29300
rect 8021 29291 8079 29297
rect 8021 29257 8033 29291
rect 8067 29288 8079 29291
rect 8110 29288 8116 29300
rect 8067 29260 8116 29288
rect 8067 29257 8079 29260
rect 8021 29251 8079 29257
rect 8110 29248 8116 29260
rect 8168 29248 8174 29300
rect 8938 29248 8944 29300
rect 8996 29248 9002 29300
rect 9306 29248 9312 29300
rect 9364 29288 9370 29300
rect 9401 29291 9459 29297
rect 9401 29288 9413 29291
rect 9364 29260 9413 29288
rect 9364 29248 9370 29260
rect 9401 29257 9413 29260
rect 9447 29257 9459 29291
rect 9401 29251 9459 29257
rect 9766 29248 9772 29300
rect 9824 29288 9830 29300
rect 9861 29291 9919 29297
rect 9861 29288 9873 29291
rect 9824 29260 9873 29288
rect 9824 29248 9830 29260
rect 9861 29257 9873 29260
rect 9907 29257 9919 29291
rect 9861 29251 9919 29257
rect 11333 29291 11391 29297
rect 11333 29257 11345 29291
rect 11379 29288 11391 29291
rect 11514 29288 11520 29300
rect 11379 29260 11520 29288
rect 11379 29257 11391 29260
rect 11333 29251 11391 29257
rect 11514 29248 11520 29260
rect 11572 29248 11578 29300
rect 11790 29248 11796 29300
rect 11848 29248 11854 29300
rect 13354 29288 13360 29300
rect 12406 29260 13360 29288
rect 8846 29220 8852 29232
rect 6564 29192 7420 29220
rect 1394 29112 1400 29164
rect 1452 29112 1458 29164
rect 1578 29112 1584 29164
rect 1636 29152 1642 29164
rect 6564 29161 6592 29192
rect 7392 29164 7420 29192
rect 8220 29192 8852 29220
rect 5997 29155 6055 29161
rect 5997 29152 6009 29155
rect 1636 29124 6009 29152
rect 1636 29112 1642 29124
rect 5997 29121 6009 29124
rect 6043 29121 6055 29155
rect 5997 29115 6055 29121
rect 6549 29155 6607 29161
rect 6549 29121 6561 29155
rect 6595 29121 6607 29155
rect 6549 29115 6607 29121
rect 6638 29112 6644 29164
rect 6696 29152 6702 29164
rect 6805 29155 6863 29161
rect 6805 29152 6817 29155
rect 6696 29124 6817 29152
rect 6696 29112 6702 29124
rect 6805 29121 6817 29124
rect 6851 29121 6863 29155
rect 6805 29115 6863 29121
rect 7374 29112 7380 29164
rect 7432 29112 7438 29164
rect 8110 29112 8116 29164
rect 8168 29152 8174 29164
rect 8220 29161 8248 29192
rect 8846 29180 8852 29192
rect 8904 29180 8910 29232
rect 8205 29155 8263 29161
rect 8205 29152 8217 29155
rect 8168 29124 8217 29152
rect 8168 29112 8174 29124
rect 8205 29121 8217 29124
rect 8251 29121 8263 29155
rect 8205 29115 8263 29121
rect 8389 29155 8447 29161
rect 8389 29121 8401 29155
rect 8435 29152 8447 29155
rect 8956 29152 8984 29248
rect 9214 29180 9220 29232
rect 9272 29220 9278 29232
rect 9585 29223 9643 29229
rect 9585 29220 9597 29223
rect 9272 29192 9597 29220
rect 9272 29180 9278 29192
rect 9585 29189 9597 29192
rect 9631 29189 9643 29223
rect 9585 29183 9643 29189
rect 10873 29223 10931 29229
rect 10873 29189 10885 29223
rect 10919 29220 10931 29223
rect 11808 29220 11836 29248
rect 10919 29192 11836 29220
rect 10919 29189 10931 29192
rect 10873 29183 10931 29189
rect 12250 29180 12256 29232
rect 12308 29180 12314 29232
rect 8435 29124 8984 29152
rect 8435 29121 8447 29124
rect 8389 29115 8447 29121
rect 9490 29112 9496 29164
rect 9548 29112 9554 29164
rect 10042 29112 10048 29164
rect 10100 29112 10106 29164
rect 10137 29155 10195 29161
rect 10137 29121 10149 29155
rect 10183 29152 10195 29155
rect 10318 29152 10324 29164
rect 10183 29124 10324 29152
rect 10183 29121 10195 29124
rect 10137 29115 10195 29121
rect 10318 29112 10324 29124
rect 10376 29112 10382 29164
rect 10597 29155 10655 29161
rect 10597 29121 10609 29155
rect 10643 29152 10655 29155
rect 10778 29152 10784 29164
rect 10643 29124 10784 29152
rect 10643 29121 10655 29124
rect 10597 29115 10655 29121
rect 10778 29112 10784 29124
rect 10836 29112 10842 29164
rect 11149 29155 11207 29161
rect 11149 29121 11161 29155
rect 11195 29152 11207 29155
rect 12406 29152 12434 29260
rect 13354 29248 13360 29260
rect 13412 29248 13418 29300
rect 13909 29291 13967 29297
rect 13909 29257 13921 29291
rect 13955 29288 13967 29291
rect 13998 29288 14004 29300
rect 13955 29260 14004 29288
rect 13955 29257 13967 29260
rect 13909 29251 13967 29257
rect 13998 29248 14004 29260
rect 14056 29248 14062 29300
rect 14182 29248 14188 29300
rect 14240 29248 14246 29300
rect 14458 29248 14464 29300
rect 14516 29248 14522 29300
rect 16485 29291 16543 29297
rect 14660 29260 15792 29288
rect 13262 29220 13268 29232
rect 13096 29192 13268 29220
rect 13096 29161 13124 29192
rect 13262 29180 13268 29192
rect 13320 29180 13326 29232
rect 14660 29229 14688 29260
rect 14645 29223 14703 29229
rect 14645 29189 14657 29223
rect 14691 29189 14703 29223
rect 14645 29183 14703 29189
rect 14734 29180 14740 29232
rect 14792 29220 14798 29232
rect 14845 29223 14903 29229
rect 14845 29220 14857 29223
rect 14792 29192 14857 29220
rect 14792 29180 14798 29192
rect 14845 29189 14857 29192
rect 14891 29189 14903 29223
rect 14845 29183 14903 29189
rect 11195 29124 12434 29152
rect 13081 29155 13139 29161
rect 11195 29121 11207 29124
rect 11149 29115 11207 29121
rect 13081 29121 13093 29155
rect 13127 29121 13139 29155
rect 13081 29115 13139 29121
rect 13170 29112 13176 29164
rect 13228 29112 13234 29164
rect 14001 29155 14059 29161
rect 14001 29121 14013 29155
rect 14047 29121 14059 29155
rect 14001 29115 14059 29121
rect 14277 29155 14335 29161
rect 14277 29121 14289 29155
rect 14323 29121 14335 29155
rect 14277 29115 14335 29121
rect 5813 29087 5871 29093
rect 5813 29053 5825 29087
rect 5859 29053 5871 29087
rect 5813 29047 5871 29053
rect 5828 29016 5856 29047
rect 8478 29044 8484 29096
rect 8536 29084 8542 29096
rect 9033 29087 9091 29093
rect 9033 29084 9045 29087
rect 8536 29056 9045 29084
rect 8536 29044 8542 29056
rect 9033 29053 9045 29056
rect 9079 29084 9091 29087
rect 9217 29087 9275 29093
rect 9217 29084 9229 29087
rect 9079 29056 9229 29084
rect 9079 29053 9091 29056
rect 9033 29047 9091 29053
rect 9217 29053 9229 29056
rect 9263 29053 9275 29087
rect 10336 29084 10364 29112
rect 10870 29084 10876 29096
rect 10336 29056 10876 29084
rect 9217 29047 9275 29053
rect 10870 29044 10876 29056
rect 10928 29044 10934 29096
rect 10965 29087 11023 29093
rect 10965 29053 10977 29087
rect 11011 29053 11023 29087
rect 10965 29047 11023 29053
rect 5994 29016 6000 29028
rect 5828 28988 6000 29016
rect 5994 28976 6000 28988
rect 6052 28976 6058 29028
rect 7929 29019 7987 29025
rect 7929 28985 7941 29019
rect 7975 29016 7987 29019
rect 9306 29016 9312 29028
rect 7975 28988 9312 29016
rect 7975 28985 7987 28988
rect 7929 28979 7987 28985
rect 9306 28976 9312 28988
rect 9364 28976 9370 29028
rect 9769 29019 9827 29025
rect 9769 28985 9781 29019
rect 9815 29016 9827 29019
rect 9950 29016 9956 29028
rect 9815 28988 9956 29016
rect 9815 28985 9827 28988
rect 9769 28979 9827 28985
rect 9950 28976 9956 28988
rect 10008 28976 10014 29028
rect 10321 29019 10379 29025
rect 10321 28985 10333 29019
rect 10367 29016 10379 29019
rect 10980 29016 11008 29047
rect 11238 29044 11244 29096
rect 11296 29084 11302 29096
rect 12069 29087 12127 29093
rect 12069 29084 12081 29087
rect 11296 29056 12081 29084
rect 11296 29044 11302 29056
rect 12069 29053 12081 29056
rect 12115 29053 12127 29087
rect 12069 29047 12127 29053
rect 12342 29016 12348 29028
rect 10367 28988 10640 29016
rect 10980 28988 12348 29016
rect 10367 28985 10379 28988
rect 10321 28979 10379 28985
rect 10612 28960 10640 28988
rect 12342 28976 12348 28988
rect 12400 29016 12406 29028
rect 12529 29019 12587 29025
rect 12529 29016 12541 29019
rect 12400 28988 12541 29016
rect 12400 28976 12406 28988
rect 12529 28985 12541 28988
rect 12575 28985 12587 29019
rect 14016 29016 14044 29115
rect 14292 29084 14320 29115
rect 14366 29112 14372 29164
rect 14424 29152 14430 29164
rect 15105 29155 15163 29161
rect 15105 29152 15117 29155
rect 14424 29124 15117 29152
rect 14424 29112 14430 29124
rect 15105 29121 15117 29124
rect 15151 29121 15163 29155
rect 15105 29115 15163 29121
rect 14292 29056 14872 29084
rect 14090 29016 14096 29028
rect 14016 28988 14096 29016
rect 12529 28979 12587 28985
rect 14090 28976 14096 28988
rect 14148 29016 14154 29028
rect 14734 29016 14740 29028
rect 14148 28988 14740 29016
rect 14148 28976 14154 28988
rect 14734 28976 14740 28988
rect 14792 28976 14798 29028
rect 14844 29016 14872 29056
rect 15764 29028 15792 29260
rect 16485 29257 16497 29291
rect 16531 29288 16543 29291
rect 16758 29288 16764 29300
rect 16531 29260 16764 29288
rect 16531 29257 16543 29260
rect 16485 29251 16543 29257
rect 16758 29248 16764 29260
rect 16816 29248 16822 29300
rect 16942 29248 16948 29300
rect 17000 29288 17006 29300
rect 17957 29291 18015 29297
rect 17957 29288 17969 29291
rect 17000 29260 17969 29288
rect 17000 29248 17006 29260
rect 17957 29257 17969 29260
rect 18003 29257 18015 29291
rect 18414 29288 18420 29300
rect 17957 29251 18015 29257
rect 18064 29260 18420 29288
rect 15933 29223 15991 29229
rect 15933 29189 15945 29223
rect 15979 29220 15991 29223
rect 16574 29220 16580 29232
rect 15979 29192 16580 29220
rect 15979 29189 15991 29192
rect 15933 29183 15991 29189
rect 16574 29180 16580 29192
rect 16632 29180 16638 29232
rect 16776 29220 16804 29248
rect 18064 29232 18092 29260
rect 18414 29248 18420 29260
rect 18472 29248 18478 29300
rect 18598 29248 18604 29300
rect 18656 29248 18662 29300
rect 18874 29248 18880 29300
rect 18932 29248 18938 29300
rect 18966 29248 18972 29300
rect 19024 29288 19030 29300
rect 19150 29288 19156 29300
rect 19024 29260 19156 29288
rect 19024 29248 19030 29260
rect 19150 29248 19156 29260
rect 19208 29248 19214 29300
rect 19260 29260 19472 29288
rect 17221 29223 17279 29229
rect 16776 29192 17080 29220
rect 16022 29112 16028 29164
rect 16080 29112 16086 29164
rect 16206 29112 16212 29164
rect 16264 29152 16270 29164
rect 16301 29155 16359 29161
rect 16301 29152 16313 29155
rect 16264 29124 16313 29152
rect 16264 29112 16270 29124
rect 16301 29121 16313 29124
rect 16347 29152 16359 29155
rect 16347 29124 16804 29152
rect 16347 29121 16359 29124
rect 16301 29115 16359 29121
rect 15654 29016 15660 29028
rect 14844 28988 15660 29016
rect 6178 28908 6184 28960
rect 6236 28908 6242 28960
rect 8294 28908 8300 28960
rect 8352 28948 8358 28960
rect 8481 28951 8539 28957
rect 8481 28948 8493 28951
rect 8352 28920 8493 28948
rect 8352 28908 8358 28920
rect 8481 28917 8493 28920
rect 8527 28917 8539 28951
rect 8481 28911 8539 28917
rect 10226 28908 10232 28960
rect 10284 28948 10290 28960
rect 10413 28951 10471 28957
rect 10413 28948 10425 28951
rect 10284 28920 10425 28948
rect 10284 28908 10290 28920
rect 10413 28917 10425 28920
rect 10459 28917 10471 28951
rect 10413 28911 10471 28917
rect 10502 28908 10508 28960
rect 10560 28908 10566 28960
rect 10594 28908 10600 28960
rect 10652 28908 10658 28960
rect 11517 28951 11575 28957
rect 11517 28917 11529 28951
rect 11563 28948 11575 28951
rect 11790 28948 11796 28960
rect 11563 28920 11796 28948
rect 11563 28917 11575 28920
rect 11517 28911 11575 28917
rect 11790 28908 11796 28920
rect 11848 28908 11854 28960
rect 12710 28908 12716 28960
rect 12768 28908 12774 28960
rect 12894 28908 12900 28960
rect 12952 28908 12958 28960
rect 14844 28957 14872 28988
rect 15654 28976 15660 28988
rect 15712 28976 15718 29028
rect 15746 28976 15752 29028
rect 15804 28976 15810 29028
rect 16040 29016 16068 29112
rect 16117 29087 16175 29093
rect 16117 29053 16129 29087
rect 16163 29084 16175 29087
rect 16666 29084 16672 29096
rect 16163 29056 16672 29084
rect 16163 29053 16175 29056
rect 16117 29047 16175 29053
rect 16666 29044 16672 29056
rect 16724 29044 16730 29096
rect 16776 29084 16804 29124
rect 16850 29112 16856 29164
rect 16908 29112 16914 29164
rect 17052 29161 17080 29192
rect 17221 29189 17233 29223
rect 17267 29189 17279 29223
rect 17221 29183 17279 29189
rect 17437 29223 17495 29229
rect 17437 29189 17449 29223
rect 17483 29220 17495 29223
rect 17483 29192 17816 29220
rect 17483 29189 17495 29192
rect 17437 29183 17495 29189
rect 17037 29155 17095 29161
rect 17037 29121 17049 29155
rect 17083 29121 17095 29155
rect 17037 29115 17095 29121
rect 17129 29087 17187 29093
rect 16776 29056 17080 29084
rect 17052 29016 17080 29056
rect 17129 29053 17141 29087
rect 17175 29084 17187 29087
rect 17236 29084 17264 29183
rect 17678 29112 17684 29164
rect 17736 29112 17742 29164
rect 17586 29084 17592 29096
rect 17175 29056 17592 29084
rect 17175 29053 17187 29056
rect 17129 29047 17187 29053
rect 17586 29044 17592 29056
rect 17644 29044 17650 29096
rect 17788 29025 17816 29192
rect 18046 29180 18052 29232
rect 18104 29180 18110 29232
rect 18506 29220 18512 29232
rect 18156 29192 18512 29220
rect 18156 29152 18184 29192
rect 18506 29180 18512 29192
rect 18564 29180 18570 29232
rect 17972 29124 18184 29152
rect 18325 29155 18383 29161
rect 17972 29093 18000 29124
rect 18325 29121 18337 29155
rect 18371 29152 18383 29155
rect 18616 29152 18644 29248
rect 18371 29124 18644 29152
rect 18785 29155 18843 29161
rect 18371 29121 18383 29124
rect 18325 29115 18383 29121
rect 18785 29121 18797 29155
rect 18831 29152 18843 29155
rect 18892 29152 18920 29248
rect 19260 29164 19288 29260
rect 19242 29152 19248 29164
rect 18831 29124 18920 29152
rect 18984 29124 19248 29152
rect 18831 29121 18843 29124
rect 18785 29115 18843 29121
rect 17957 29087 18015 29093
rect 17957 29053 17969 29087
rect 18003 29053 18015 29087
rect 17957 29047 18015 29053
rect 18049 29087 18107 29093
rect 18049 29053 18061 29087
rect 18095 29084 18107 29087
rect 18984 29084 19012 29124
rect 19242 29112 19248 29124
rect 19300 29112 19306 29164
rect 19334 29112 19340 29164
rect 19392 29112 19398 29164
rect 19444 29161 19472 29260
rect 20990 29248 20996 29300
rect 21048 29248 21054 29300
rect 23290 29248 23296 29300
rect 23348 29248 23354 29300
rect 24026 29248 24032 29300
rect 24084 29288 24090 29300
rect 24121 29291 24179 29297
rect 24121 29288 24133 29291
rect 24084 29260 24133 29288
rect 24084 29248 24090 29260
rect 24121 29257 24133 29260
rect 24167 29257 24179 29291
rect 24121 29251 24179 29257
rect 21266 29220 21272 29232
rect 19628 29192 21272 29220
rect 19429 29155 19487 29161
rect 19429 29121 19441 29155
rect 19475 29121 19487 29155
rect 19429 29115 19487 29121
rect 19518 29112 19524 29164
rect 19576 29152 19582 29164
rect 19628 29161 19656 29192
rect 21266 29180 21272 29192
rect 21324 29220 21330 29232
rect 23308 29220 23336 29248
rect 21324 29192 21864 29220
rect 21324 29180 21330 29192
rect 19613 29155 19671 29161
rect 19613 29152 19625 29155
rect 19576 29124 19625 29152
rect 19576 29112 19582 29124
rect 19613 29121 19625 29124
rect 19659 29121 19671 29155
rect 19613 29115 19671 29121
rect 19702 29112 19708 29164
rect 19760 29112 19766 29164
rect 19886 29161 19892 29164
rect 19880 29152 19892 29161
rect 19847 29124 19892 29152
rect 19880 29115 19892 29124
rect 19886 29112 19892 29115
rect 19944 29112 19950 29164
rect 21085 29155 21143 29161
rect 21085 29121 21097 29155
rect 21131 29152 21143 29155
rect 21174 29152 21180 29164
rect 21131 29124 21180 29152
rect 21131 29121 21143 29124
rect 21085 29115 21143 29121
rect 21174 29112 21180 29124
rect 21232 29112 21238 29164
rect 21836 29161 21864 29192
rect 23308 29192 24256 29220
rect 21821 29155 21879 29161
rect 21821 29121 21833 29155
rect 21867 29121 21879 29155
rect 22077 29155 22135 29161
rect 22077 29152 22089 29155
rect 21821 29115 21879 29121
rect 21928 29124 22089 29152
rect 18095 29056 19012 29084
rect 19061 29087 19119 29093
rect 18095 29053 18107 29056
rect 18049 29047 18107 29053
rect 19061 29053 19073 29087
rect 19107 29084 19119 29087
rect 19720 29084 19748 29112
rect 21928 29084 21956 29124
rect 22077 29121 22089 29124
rect 22123 29121 22135 29155
rect 23308 29152 23336 29192
rect 23477 29155 23535 29161
rect 23477 29152 23489 29155
rect 23308 29124 23489 29152
rect 22077 29115 22135 29121
rect 23477 29121 23489 29124
rect 23523 29121 23535 29155
rect 23477 29115 23535 29121
rect 23750 29112 23756 29164
rect 23808 29112 23814 29164
rect 23934 29112 23940 29164
rect 23992 29112 23998 29164
rect 24228 29161 24256 29192
rect 24213 29155 24271 29161
rect 24213 29121 24225 29155
rect 24259 29121 24271 29155
rect 24213 29115 24271 29121
rect 24397 29155 24455 29161
rect 24397 29121 24409 29155
rect 24443 29121 24455 29155
rect 24397 29115 24455 29121
rect 23661 29087 23719 29093
rect 23661 29084 23673 29087
rect 19107 29056 19748 29084
rect 21284 29056 21956 29084
rect 23216 29056 23673 29084
rect 19107 29053 19119 29056
rect 19061 29047 19119 29053
rect 17773 29019 17831 29025
rect 17773 29016 17785 29019
rect 16040 28988 16896 29016
rect 17052 28988 17785 29016
rect 14829 28951 14887 28957
rect 14829 28917 14841 28951
rect 14875 28917 14887 28951
rect 14829 28911 14887 28917
rect 15013 28951 15071 28957
rect 15013 28917 15025 28951
rect 15059 28948 15071 28951
rect 16206 28948 16212 28960
rect 15059 28920 16212 28948
rect 15059 28917 15071 28920
rect 15013 28911 15071 28917
rect 16206 28908 16212 28920
rect 16264 28908 16270 28960
rect 16669 28951 16727 28957
rect 16669 28917 16681 28951
rect 16715 28948 16727 28951
rect 16758 28948 16764 28960
rect 16715 28920 16764 28948
rect 16715 28917 16727 28920
rect 16669 28911 16727 28917
rect 16758 28908 16764 28920
rect 16816 28908 16822 28960
rect 16868 28948 16896 28988
rect 17773 28985 17785 28988
rect 17819 28985 17831 29019
rect 18141 29019 18199 29025
rect 18141 29016 18153 29019
rect 17773 28979 17831 28985
rect 17880 28988 18153 29016
rect 17405 28951 17463 28957
rect 17405 28948 17417 28951
rect 16868 28920 17417 28948
rect 17405 28917 17417 28920
rect 17451 28917 17463 28951
rect 17405 28911 17463 28917
rect 17494 28908 17500 28960
rect 17552 28948 17558 28960
rect 17589 28951 17647 28957
rect 17589 28948 17601 28951
rect 17552 28920 17601 28948
rect 17552 28908 17558 28920
rect 17589 28917 17601 28920
rect 17635 28948 17647 28951
rect 17880 28948 17908 28988
rect 18141 28985 18153 28988
rect 18187 28985 18199 29019
rect 18141 28979 18199 28985
rect 18509 29019 18567 29025
rect 18509 28985 18521 29019
rect 18555 29016 18567 29019
rect 18969 29019 19027 29025
rect 18555 28988 18920 29016
rect 18555 28985 18567 28988
rect 18509 28979 18567 28985
rect 17635 28920 17908 28948
rect 17635 28917 17647 28920
rect 17589 28911 17647 28917
rect 18598 28908 18604 28960
rect 18656 28908 18662 28960
rect 18892 28948 18920 28988
rect 18969 28985 18981 29019
rect 19015 29016 19027 29019
rect 19150 29016 19156 29028
rect 19015 28988 19156 29016
rect 19015 28985 19027 28988
rect 18969 28979 19027 28985
rect 19150 28976 19156 28988
rect 19208 28976 19214 29028
rect 21284 29025 21312 29056
rect 23216 29025 23244 29056
rect 23661 29053 23673 29056
rect 23707 29084 23719 29087
rect 24412 29084 24440 29115
rect 23707 29056 24440 29084
rect 23707 29053 23719 29056
rect 23661 29047 23719 29053
rect 21269 29019 21327 29025
rect 21269 28985 21281 29019
rect 21315 28985 21327 29019
rect 21269 28979 21327 28985
rect 23201 29019 23259 29025
rect 23201 28985 23213 29019
rect 23247 28985 23259 29019
rect 23201 28979 23259 28985
rect 20346 28948 20352 28960
rect 18892 28920 20352 28948
rect 20346 28908 20352 28920
rect 20404 28908 20410 28960
rect 23290 28908 23296 28960
rect 23348 28908 23354 28960
rect 24210 28908 24216 28960
rect 24268 28908 24274 28960
rect 1104 28858 34868 28880
rect 1104 28806 5170 28858
rect 5222 28806 5234 28858
rect 5286 28806 5298 28858
rect 5350 28806 5362 28858
rect 5414 28806 5426 28858
rect 5478 28806 13611 28858
rect 13663 28806 13675 28858
rect 13727 28806 13739 28858
rect 13791 28806 13803 28858
rect 13855 28806 13867 28858
rect 13919 28806 22052 28858
rect 22104 28806 22116 28858
rect 22168 28806 22180 28858
rect 22232 28806 22244 28858
rect 22296 28806 22308 28858
rect 22360 28806 30493 28858
rect 30545 28806 30557 28858
rect 30609 28806 30621 28858
rect 30673 28806 30685 28858
rect 30737 28806 30749 28858
rect 30801 28806 34868 28858
rect 1104 28784 34868 28806
rect 6549 28747 6607 28753
rect 6549 28713 6561 28747
rect 6595 28744 6607 28747
rect 6638 28744 6644 28756
rect 6595 28716 6644 28744
rect 6595 28713 6607 28716
rect 6549 28707 6607 28713
rect 6638 28704 6644 28716
rect 6696 28704 6702 28756
rect 8297 28747 8355 28753
rect 8297 28713 8309 28747
rect 8343 28713 8355 28747
rect 8297 28707 8355 28713
rect 8757 28747 8815 28753
rect 8757 28713 8769 28747
rect 8803 28744 8815 28747
rect 9306 28744 9312 28756
rect 8803 28716 9312 28744
rect 8803 28713 8815 28716
rect 8757 28707 8815 28713
rect 8312 28676 8340 28707
rect 9306 28704 9312 28716
rect 9364 28704 9370 28756
rect 10502 28704 10508 28756
rect 10560 28704 10566 28756
rect 10686 28704 10692 28756
rect 10744 28704 10750 28756
rect 10781 28747 10839 28753
rect 10781 28713 10793 28747
rect 10827 28744 10839 28747
rect 11606 28744 11612 28756
rect 10827 28716 11612 28744
rect 10827 28713 10839 28716
rect 10781 28707 10839 28713
rect 11606 28704 11612 28716
rect 11664 28704 11670 28756
rect 12158 28744 12164 28756
rect 11808 28716 12164 28744
rect 10520 28676 10548 28704
rect 8312 28648 10548 28676
rect 10704 28676 10732 28704
rect 10873 28679 10931 28685
rect 10873 28676 10885 28679
rect 10704 28648 10885 28676
rect 10873 28645 10885 28648
rect 10919 28645 10931 28679
rect 10873 28639 10931 28645
rect 7745 28611 7803 28617
rect 7745 28577 7757 28611
rect 7791 28608 7803 28611
rect 8294 28608 8300 28620
rect 7791 28580 8300 28608
rect 7791 28577 7803 28580
rect 7745 28571 7803 28577
rect 8294 28568 8300 28580
rect 8352 28568 8358 28620
rect 8665 28611 8723 28617
rect 8665 28577 8677 28611
rect 8711 28608 8723 28611
rect 8938 28608 8944 28620
rect 8711 28580 8944 28608
rect 8711 28577 8723 28580
rect 8665 28571 8723 28577
rect 8938 28568 8944 28580
rect 8996 28608 9002 28620
rect 9490 28608 9496 28620
rect 8996 28580 9496 28608
rect 8996 28568 9002 28580
rect 9490 28568 9496 28580
rect 9548 28608 9554 28620
rect 9585 28611 9643 28617
rect 9585 28608 9597 28611
rect 9548 28580 9597 28608
rect 9548 28568 9554 28580
rect 9585 28577 9597 28580
rect 9631 28577 9643 28611
rect 9585 28571 9643 28577
rect 9858 28568 9864 28620
rect 9916 28608 9922 28620
rect 11808 28617 11836 28716
rect 12158 28704 12164 28716
rect 12216 28704 12222 28756
rect 13170 28704 13176 28756
rect 13228 28704 13234 28756
rect 14277 28747 14335 28753
rect 14277 28713 14289 28747
rect 14323 28744 14335 28747
rect 14366 28744 14372 28756
rect 14323 28716 14372 28744
rect 14323 28713 14335 28716
rect 14277 28707 14335 28713
rect 14366 28704 14372 28716
rect 14424 28704 14430 28756
rect 15933 28747 15991 28753
rect 15933 28713 15945 28747
rect 15979 28744 15991 28747
rect 16850 28744 16856 28756
rect 15979 28716 16856 28744
rect 15979 28713 15991 28716
rect 15933 28707 15991 28713
rect 16850 28704 16856 28716
rect 16908 28704 16914 28756
rect 17586 28704 17592 28756
rect 17644 28704 17650 28756
rect 17678 28704 17684 28756
rect 17736 28704 17742 28756
rect 19429 28747 19487 28753
rect 19429 28713 19441 28747
rect 19475 28744 19487 28747
rect 19702 28744 19708 28756
rect 19475 28716 19708 28744
rect 19475 28713 19487 28716
rect 19429 28707 19487 28713
rect 19702 28704 19708 28716
rect 19760 28704 19766 28756
rect 20165 28747 20223 28753
rect 20165 28713 20177 28747
rect 20211 28744 20223 28747
rect 20438 28744 20444 28756
rect 20211 28716 20444 28744
rect 20211 28713 20223 28716
rect 20165 28707 20223 28713
rect 20438 28704 20444 28716
rect 20496 28704 20502 28756
rect 20530 28704 20536 28756
rect 20588 28704 20594 28756
rect 22738 28704 22744 28756
rect 22796 28704 22802 28756
rect 23017 28747 23075 28753
rect 23017 28713 23029 28747
rect 23063 28744 23075 28747
rect 23290 28744 23296 28756
rect 23063 28716 23296 28744
rect 23063 28713 23075 28716
rect 23017 28707 23075 28713
rect 12912 28648 13584 28676
rect 12912 28620 12940 28648
rect 11793 28611 11851 28617
rect 11793 28608 11805 28611
rect 9916 28580 11805 28608
rect 9916 28568 9922 28580
rect 11793 28577 11805 28580
rect 11839 28577 11851 28611
rect 11793 28571 11851 28577
rect 6178 28500 6184 28552
rect 6236 28540 6242 28552
rect 6365 28543 6423 28549
rect 6365 28540 6377 28543
rect 6236 28512 6377 28540
rect 6236 28500 6242 28512
rect 6365 28509 6377 28512
rect 6411 28509 6423 28543
rect 6365 28503 6423 28509
rect 7561 28543 7619 28549
rect 7561 28509 7573 28543
rect 7607 28540 7619 28543
rect 8021 28543 8079 28549
rect 8021 28540 8033 28543
rect 7607 28512 8033 28540
rect 7607 28509 7619 28512
rect 7561 28503 7619 28509
rect 8021 28509 8033 28512
rect 8067 28540 8079 28543
rect 8110 28540 8116 28552
rect 8067 28512 8116 28540
rect 8067 28509 8079 28512
rect 8021 28503 8079 28509
rect 8110 28500 8116 28512
rect 8168 28500 8174 28552
rect 8202 28500 8208 28552
rect 8260 28500 8266 28552
rect 8478 28500 8484 28552
rect 8536 28500 8542 28552
rect 9769 28543 9827 28549
rect 9769 28509 9781 28543
rect 9815 28509 9827 28543
rect 9769 28503 9827 28509
rect 8757 28475 8815 28481
rect 8757 28441 8769 28475
rect 8803 28472 8815 28475
rect 9214 28472 9220 28484
rect 8803 28444 9220 28472
rect 8803 28441 8815 28444
rect 8757 28435 8815 28441
rect 9214 28432 9220 28444
rect 9272 28432 9278 28484
rect 9784 28472 9812 28503
rect 9950 28500 9956 28552
rect 10008 28540 10014 28552
rect 10137 28543 10195 28549
rect 10137 28540 10149 28543
rect 10008 28512 10149 28540
rect 10008 28500 10014 28512
rect 10137 28509 10149 28512
rect 10183 28509 10195 28543
rect 10137 28503 10195 28509
rect 10226 28500 10232 28552
rect 10284 28500 10290 28552
rect 10318 28500 10324 28552
rect 10376 28540 10382 28552
rect 10505 28543 10563 28549
rect 10505 28540 10517 28543
rect 10376 28512 10517 28540
rect 10376 28500 10382 28512
rect 10505 28509 10517 28512
rect 10551 28509 10563 28543
rect 10505 28503 10563 28509
rect 10597 28543 10655 28549
rect 10597 28509 10609 28543
rect 10643 28540 10655 28543
rect 10778 28540 10784 28552
rect 10643 28512 10784 28540
rect 10643 28509 10655 28512
rect 10597 28503 10655 28509
rect 10778 28500 10784 28512
rect 10836 28500 10842 28552
rect 10870 28500 10876 28552
rect 10928 28540 10934 28552
rect 11425 28543 11483 28549
rect 11425 28540 11437 28543
rect 10928 28512 11437 28540
rect 10928 28500 10934 28512
rect 11425 28509 11437 28512
rect 11471 28509 11483 28543
rect 11425 28503 11483 28509
rect 11698 28500 11704 28552
rect 11756 28500 11762 28552
rect 11808 28540 11836 28571
rect 12894 28568 12900 28620
rect 12952 28568 12958 28620
rect 13354 28568 13360 28620
rect 13412 28568 13418 28620
rect 13556 28608 13584 28648
rect 16666 28636 16672 28688
rect 16724 28676 16730 28688
rect 17696 28676 17724 28704
rect 20622 28676 20628 28688
rect 16724 28648 17724 28676
rect 20088 28648 20628 28676
rect 16724 28636 16730 28648
rect 20088 28620 20116 28648
rect 20622 28636 20628 28648
rect 20680 28636 20686 28688
rect 23032 28676 23060 28707
rect 23290 28704 23296 28716
rect 23348 28704 23354 28756
rect 22572 28648 23060 28676
rect 15657 28611 15715 28617
rect 13556 28580 13676 28608
rect 11808 28512 12434 28540
rect 11514 28472 11520 28484
rect 9784 28444 11520 28472
rect 11514 28432 11520 28444
rect 11572 28432 11578 28484
rect 11716 28472 11744 28500
rect 12038 28475 12096 28481
rect 12038 28472 12050 28475
rect 11716 28444 12050 28472
rect 12038 28441 12050 28444
rect 12084 28441 12096 28475
rect 12406 28472 12434 28512
rect 12802 28500 12808 28552
rect 12860 28540 12866 28552
rect 13265 28543 13323 28549
rect 13265 28540 13277 28543
rect 12860 28512 13277 28540
rect 12860 28500 12866 28512
rect 13265 28509 13277 28512
rect 13311 28509 13323 28543
rect 13265 28503 13323 28509
rect 13538 28500 13544 28552
rect 13596 28500 13602 28552
rect 13648 28549 13676 28580
rect 15657 28577 15669 28611
rect 15703 28608 15715 28611
rect 15703 28580 16712 28608
rect 15703 28577 15715 28580
rect 15657 28571 15715 28577
rect 16684 28552 16712 28580
rect 17310 28568 17316 28620
rect 17368 28608 17374 28620
rect 18046 28608 18052 28620
rect 17368 28580 18052 28608
rect 17368 28568 17374 28580
rect 18046 28568 18052 28580
rect 18104 28568 18110 28620
rect 18230 28568 18236 28620
rect 18288 28568 18294 28620
rect 18598 28568 18604 28620
rect 18656 28608 18662 28620
rect 18969 28611 19027 28617
rect 18969 28608 18981 28611
rect 18656 28580 18981 28608
rect 18656 28568 18662 28580
rect 18969 28577 18981 28580
rect 19015 28577 19027 28611
rect 18969 28571 19027 28577
rect 20070 28568 20076 28620
rect 20128 28568 20134 28620
rect 20162 28568 20168 28620
rect 20220 28608 20226 28620
rect 20717 28611 20775 28617
rect 20717 28608 20729 28611
rect 20220 28580 20729 28608
rect 20220 28568 20226 28580
rect 13633 28543 13691 28549
rect 13633 28509 13645 28543
rect 13679 28509 13691 28543
rect 15749 28543 15807 28549
rect 15749 28540 15761 28543
rect 13633 28503 13691 28509
rect 15212 28512 15761 28540
rect 15212 28484 15240 28512
rect 15749 28509 15761 28512
rect 15795 28509 15807 28543
rect 15749 28503 15807 28509
rect 15933 28543 15991 28549
rect 15933 28509 15945 28543
rect 15979 28509 15991 28543
rect 15933 28503 15991 28509
rect 13906 28472 13912 28484
rect 12406 28444 13912 28472
rect 12038 28435 12096 28441
rect 13906 28432 13912 28444
rect 13964 28432 13970 28484
rect 15194 28432 15200 28484
rect 15252 28432 15258 28484
rect 15378 28432 15384 28484
rect 15436 28481 15442 28484
rect 15436 28435 15448 28481
rect 15436 28432 15442 28435
rect 7190 28364 7196 28416
rect 7248 28404 7254 28416
rect 7377 28407 7435 28413
rect 7377 28404 7389 28407
rect 7248 28376 7389 28404
rect 7248 28364 7254 28376
rect 7377 28373 7389 28376
rect 7423 28373 7435 28407
rect 7377 28367 7435 28373
rect 7466 28364 7472 28416
rect 7524 28404 7530 28416
rect 7837 28407 7895 28413
rect 7837 28404 7849 28407
rect 7524 28376 7849 28404
rect 7524 28364 7530 28376
rect 7837 28373 7849 28376
rect 7883 28373 7895 28407
rect 7837 28367 7895 28373
rect 9030 28364 9036 28416
rect 9088 28364 9094 28416
rect 9950 28364 9956 28416
rect 10008 28364 10014 28416
rect 10413 28407 10471 28413
rect 10413 28373 10425 28407
rect 10459 28404 10471 28407
rect 10594 28404 10600 28416
rect 10459 28376 10600 28404
rect 10459 28373 10471 28376
rect 10413 28367 10471 28373
rect 10594 28364 10600 28376
rect 10652 28364 10658 28416
rect 11698 28364 11704 28416
rect 11756 28404 11762 28416
rect 13817 28407 13875 28413
rect 13817 28404 13829 28407
rect 11756 28376 13829 28404
rect 11756 28364 11762 28376
rect 13817 28373 13829 28376
rect 13863 28404 13875 28407
rect 14274 28404 14280 28416
rect 13863 28376 14280 28404
rect 13863 28373 13875 28376
rect 13817 28367 13875 28373
rect 14274 28364 14280 28376
rect 14332 28364 14338 28416
rect 15764 28404 15792 28503
rect 15948 28472 15976 28503
rect 16022 28500 16028 28552
rect 16080 28500 16086 28552
rect 16666 28500 16672 28552
rect 16724 28500 16730 28552
rect 16758 28500 16764 28552
rect 16816 28500 16822 28552
rect 20254 28500 20260 28552
rect 20312 28540 20318 28552
rect 20640 28549 20668 28580
rect 20717 28577 20729 28580
rect 20763 28577 20775 28611
rect 20717 28571 20775 28577
rect 20990 28568 20996 28620
rect 21048 28608 21054 28620
rect 21269 28611 21327 28617
rect 21269 28608 21281 28611
rect 21048 28580 21281 28608
rect 21048 28568 21054 28580
rect 21269 28577 21281 28580
rect 21315 28577 21327 28611
rect 22572 28608 22600 28648
rect 21269 28571 21327 28577
rect 22480 28580 22600 28608
rect 22480 28549 22508 28580
rect 22738 28568 22744 28620
rect 22796 28608 22802 28620
rect 22796 28580 23244 28608
rect 22796 28568 22802 28580
rect 20349 28543 20407 28549
rect 20349 28540 20361 28543
rect 20312 28512 20361 28540
rect 20312 28500 20318 28512
rect 20349 28509 20361 28512
rect 20395 28509 20407 28543
rect 20349 28503 20407 28509
rect 20625 28543 20683 28549
rect 20625 28509 20637 28543
rect 20671 28540 20683 28543
rect 22465 28543 22523 28549
rect 20671 28512 20705 28540
rect 20671 28509 20683 28512
rect 20625 28503 20683 28509
rect 22465 28509 22477 28543
rect 22511 28509 22523 28543
rect 22465 28503 22523 28509
rect 22557 28543 22615 28549
rect 22557 28509 22569 28543
rect 22603 28509 22615 28543
rect 22557 28503 22615 28509
rect 17494 28472 17500 28484
rect 15948 28444 17500 28472
rect 17494 28432 17500 28444
rect 17552 28432 17558 28484
rect 22572 28472 22600 28503
rect 22646 28500 22652 28552
rect 22704 28540 22710 28552
rect 23216 28549 23244 28580
rect 22833 28543 22891 28549
rect 22833 28540 22845 28543
rect 22704 28512 22845 28540
rect 22704 28500 22710 28512
rect 22833 28509 22845 28512
rect 22879 28540 22891 28543
rect 22925 28543 22983 28549
rect 22925 28540 22937 28543
rect 22879 28512 22937 28540
rect 22879 28509 22891 28512
rect 22833 28503 22891 28509
rect 22925 28509 22937 28512
rect 22971 28509 22983 28543
rect 22925 28503 22983 28509
rect 23201 28543 23259 28549
rect 23201 28509 23213 28543
rect 23247 28509 23259 28543
rect 23201 28503 23259 28509
rect 23293 28543 23351 28549
rect 23293 28509 23305 28543
rect 23339 28540 23351 28543
rect 24210 28540 24216 28552
rect 23339 28512 24216 28540
rect 23339 28509 23351 28512
rect 23293 28503 23351 28509
rect 23308 28472 23336 28503
rect 24210 28500 24216 28512
rect 24268 28500 24274 28552
rect 22572 28444 23336 28472
rect 17310 28404 17316 28416
rect 15764 28376 17316 28404
rect 17310 28364 17316 28376
rect 17368 28364 17374 28416
rect 17402 28364 17408 28416
rect 17460 28364 17466 28416
rect 18414 28364 18420 28416
rect 18472 28364 18478 28416
rect 22278 28364 22284 28416
rect 22336 28364 22342 28416
rect 22554 28364 22560 28416
rect 22612 28404 22618 28416
rect 23477 28407 23535 28413
rect 23477 28404 23489 28407
rect 22612 28376 23489 28404
rect 22612 28364 22618 28376
rect 23477 28373 23489 28376
rect 23523 28373 23535 28407
rect 23477 28367 23535 28373
rect 1104 28314 35027 28336
rect 1104 28262 9390 28314
rect 9442 28262 9454 28314
rect 9506 28262 9518 28314
rect 9570 28262 9582 28314
rect 9634 28262 9646 28314
rect 9698 28262 17831 28314
rect 17883 28262 17895 28314
rect 17947 28262 17959 28314
rect 18011 28262 18023 28314
rect 18075 28262 18087 28314
rect 18139 28262 26272 28314
rect 26324 28262 26336 28314
rect 26388 28262 26400 28314
rect 26452 28262 26464 28314
rect 26516 28262 26528 28314
rect 26580 28262 34713 28314
rect 34765 28262 34777 28314
rect 34829 28262 34841 28314
rect 34893 28262 34905 28314
rect 34957 28262 34969 28314
rect 35021 28262 35027 28314
rect 1104 28240 35027 28262
rect 7190 28160 7196 28212
rect 7248 28160 7254 28212
rect 7469 28203 7527 28209
rect 7469 28169 7481 28203
rect 7515 28169 7527 28203
rect 7469 28163 7527 28169
rect 7009 28067 7067 28073
rect 7009 28033 7021 28067
rect 7055 28064 7067 28067
rect 7208 28064 7236 28160
rect 7484 28132 7512 28163
rect 8202 28160 8208 28212
rect 8260 28200 8266 28212
rect 9033 28203 9091 28209
rect 9033 28200 9045 28203
rect 8260 28172 9045 28200
rect 8260 28160 8266 28172
rect 9033 28169 9045 28172
rect 9079 28169 9091 28203
rect 9033 28163 9091 28169
rect 9950 28160 9956 28212
rect 10008 28160 10014 28212
rect 10594 28160 10600 28212
rect 10652 28200 10658 28212
rect 11241 28203 11299 28209
rect 11241 28200 11253 28203
rect 10652 28172 11253 28200
rect 10652 28160 10658 28172
rect 11241 28169 11253 28172
rect 11287 28169 11299 28203
rect 11241 28163 11299 28169
rect 11514 28160 11520 28212
rect 11572 28160 11578 28212
rect 11882 28160 11888 28212
rect 11940 28160 11946 28212
rect 12621 28203 12679 28209
rect 12621 28169 12633 28203
rect 12667 28200 12679 28203
rect 13354 28200 13360 28212
rect 12667 28172 13360 28200
rect 12667 28169 12679 28172
rect 12621 28163 12679 28169
rect 7806 28135 7864 28141
rect 7806 28132 7818 28135
rect 7484 28104 7818 28132
rect 7806 28101 7818 28104
rect 7852 28101 7864 28135
rect 9968 28132 9996 28160
rect 10106 28135 10164 28141
rect 10106 28132 10118 28135
rect 9968 28104 10118 28132
rect 7806 28095 7864 28101
rect 10106 28101 10118 28104
rect 10152 28101 10164 28135
rect 11900 28132 11928 28160
rect 10106 28095 10164 28101
rect 11716 28104 11928 28132
rect 12161 28135 12219 28141
rect 7055 28036 7236 28064
rect 7285 28067 7343 28073
rect 7055 28033 7067 28036
rect 7009 28027 7067 28033
rect 7285 28033 7297 28067
rect 7331 28064 7343 28067
rect 7466 28064 7472 28076
rect 7331 28036 7472 28064
rect 7331 28033 7343 28036
rect 7285 28027 7343 28033
rect 7466 28024 7472 28036
rect 7524 28024 7530 28076
rect 9214 28024 9220 28076
rect 9272 28064 9278 28076
rect 11716 28073 11744 28104
rect 12161 28101 12173 28135
rect 12207 28132 12219 28135
rect 12342 28132 12348 28144
rect 12207 28104 12348 28132
rect 12207 28101 12219 28104
rect 12161 28095 12219 28101
rect 12342 28092 12348 28104
rect 12400 28092 12406 28144
rect 9585 28067 9643 28073
rect 9585 28064 9597 28067
rect 9272 28036 9597 28064
rect 9272 28024 9278 28036
rect 9585 28033 9597 28036
rect 9631 28033 9643 28067
rect 9585 28027 9643 28033
rect 11701 28067 11759 28073
rect 11701 28033 11713 28067
rect 11747 28033 11759 28067
rect 11701 28027 11759 28033
rect 11790 28024 11796 28076
rect 11848 28024 11854 28076
rect 12710 28024 12716 28076
rect 12768 28024 12774 28076
rect 13004 28073 13032 28172
rect 13354 28160 13360 28172
rect 13412 28160 13418 28212
rect 13449 28203 13507 28209
rect 13449 28169 13461 28203
rect 13495 28200 13507 28203
rect 13538 28200 13544 28212
rect 13495 28172 13544 28200
rect 13495 28169 13507 28172
rect 13449 28163 13507 28169
rect 13464 28132 13492 28163
rect 13538 28160 13544 28172
rect 13596 28160 13602 28212
rect 15378 28160 15384 28212
rect 15436 28200 15442 28212
rect 15473 28203 15531 28209
rect 15473 28200 15485 28203
rect 15436 28172 15485 28200
rect 15436 28160 15442 28172
rect 15473 28169 15485 28172
rect 15519 28169 15531 28203
rect 15473 28163 15531 28169
rect 16206 28160 16212 28212
rect 16264 28160 16270 28212
rect 18049 28203 18107 28209
rect 18049 28169 18061 28203
rect 18095 28200 18107 28203
rect 18230 28200 18236 28212
rect 18095 28172 18236 28200
rect 18095 28169 18107 28172
rect 18049 28163 18107 28169
rect 18230 28160 18236 28172
rect 18288 28160 18294 28212
rect 19518 28200 19524 28212
rect 19306 28172 19524 28200
rect 13096 28104 13492 28132
rect 16224 28132 16252 28160
rect 19306 28132 19334 28172
rect 19518 28160 19524 28172
rect 19576 28160 19582 28212
rect 19705 28203 19763 28209
rect 19705 28169 19717 28203
rect 19751 28200 19763 28203
rect 20070 28200 20076 28212
rect 19751 28172 20076 28200
rect 19751 28169 19763 28172
rect 19705 28163 19763 28169
rect 20070 28160 20076 28172
rect 20128 28160 20134 28212
rect 16224 28104 16344 28132
rect 13096 28073 13124 28104
rect 12989 28067 13047 28073
rect 12989 28033 13001 28067
rect 13035 28033 13047 28067
rect 12989 28027 13047 28033
rect 13081 28067 13139 28073
rect 13081 28033 13093 28067
rect 13127 28033 13139 28067
rect 13081 28027 13139 28033
rect 13170 28024 13176 28076
rect 13228 28064 13234 28076
rect 13357 28067 13415 28073
rect 13357 28064 13369 28067
rect 13228 28036 13369 28064
rect 13228 28024 13234 28036
rect 13357 28033 13369 28036
rect 13403 28033 13415 28067
rect 13357 28027 13415 28033
rect 13541 28067 13599 28073
rect 13541 28033 13553 28067
rect 13587 28033 13599 28067
rect 13541 28027 13599 28033
rect 7374 27956 7380 28008
rect 7432 27996 7438 28008
rect 7561 27999 7619 28005
rect 7561 27996 7573 27999
rect 7432 27968 7573 27996
rect 7432 27956 7438 27968
rect 7561 27965 7573 27968
rect 7607 27965 7619 27999
rect 7561 27959 7619 27965
rect 9858 27956 9864 28008
rect 9916 27956 9922 28008
rect 12805 27999 12863 28005
rect 12805 27965 12817 27999
rect 12851 27996 12863 27999
rect 12894 27996 12900 28008
rect 12851 27968 12900 27996
rect 12851 27965 12863 27968
rect 12805 27959 12863 27965
rect 12894 27956 12900 27968
rect 12952 27956 12958 28008
rect 13262 27956 13268 28008
rect 13320 27996 13326 28008
rect 13556 27996 13584 28027
rect 13906 28024 13912 28076
rect 13964 28024 13970 28076
rect 14182 28073 14188 28076
rect 14176 28027 14188 28073
rect 14182 28024 14188 28027
rect 14240 28024 14246 28076
rect 15930 28024 15936 28076
rect 15988 28064 15994 28076
rect 16316 28073 16344 28104
rect 16868 28104 17816 28132
rect 16209 28067 16267 28073
rect 16209 28064 16221 28067
rect 15988 28036 16221 28064
rect 15988 28024 15994 28036
rect 16209 28033 16221 28036
rect 16255 28033 16267 28067
rect 16209 28027 16267 28033
rect 16301 28067 16359 28073
rect 16301 28033 16313 28067
rect 16347 28033 16359 28067
rect 16868 28064 16896 28104
rect 17788 28076 17816 28104
rect 18340 28104 19334 28132
rect 21253 28135 21311 28141
rect 16301 28027 16359 28033
rect 16785 28036 16896 28064
rect 16936 28067 16994 28073
rect 13320 27968 13584 27996
rect 16117 27999 16175 28005
rect 13320 27956 13326 27968
rect 16117 27965 16129 27999
rect 16163 27996 16175 27999
rect 16163 27968 16252 27996
rect 16163 27965 16175 27968
rect 16117 27959 16175 27965
rect 8938 27888 8944 27940
rect 8996 27888 9002 27940
rect 12250 27888 12256 27940
rect 12308 27928 12314 27940
rect 16224 27937 16252 27968
rect 16482 27956 16488 28008
rect 16540 27956 16546 28008
rect 16666 27956 16672 28008
rect 16724 27996 16730 28008
rect 16785 27996 16813 28036
rect 16936 28033 16948 28067
rect 16982 28064 16994 28067
rect 17402 28064 17408 28076
rect 16982 28036 17408 28064
rect 16982 28033 16994 28036
rect 16936 28027 16994 28033
rect 17402 28024 17408 28036
rect 17460 28024 17466 28076
rect 17770 28024 17776 28076
rect 17828 28064 17834 28076
rect 18340 28073 18368 28104
rect 21253 28101 21265 28135
rect 21299 28132 21311 28135
rect 21358 28132 21364 28144
rect 21299 28104 21364 28132
rect 21299 28101 21311 28104
rect 21253 28095 21311 28101
rect 21358 28092 21364 28104
rect 21416 28092 21422 28144
rect 21453 28135 21511 28141
rect 21453 28101 21465 28135
rect 21499 28132 21511 28135
rect 21542 28132 21548 28144
rect 21499 28104 21548 28132
rect 21499 28101 21511 28104
rect 21453 28095 21511 28101
rect 21542 28092 21548 28104
rect 21600 28092 21606 28144
rect 22189 28135 22247 28141
rect 22189 28101 22201 28135
rect 22235 28132 22247 28135
rect 22554 28132 22560 28144
rect 22235 28104 22560 28132
rect 22235 28101 22247 28104
rect 22189 28095 22247 28101
rect 22554 28092 22560 28104
rect 22612 28092 22618 28144
rect 18325 28067 18383 28073
rect 18325 28064 18337 28067
rect 17828 28036 18337 28064
rect 17828 28024 17834 28036
rect 18325 28033 18337 28036
rect 18371 28033 18383 28067
rect 18325 28027 18383 28033
rect 18414 28024 18420 28076
rect 18472 28064 18478 28076
rect 18581 28067 18639 28073
rect 18581 28064 18593 28067
rect 18472 28036 18593 28064
rect 18472 28024 18478 28036
rect 18581 28033 18593 28036
rect 18627 28033 18639 28067
rect 18581 28027 18639 28033
rect 20346 28024 20352 28076
rect 20404 28024 20410 28076
rect 21910 28024 21916 28076
rect 21968 28064 21974 28076
rect 22005 28067 22063 28073
rect 22005 28064 22017 28067
rect 21968 28036 22017 28064
rect 21968 28024 21974 28036
rect 22005 28033 22017 28036
rect 22051 28033 22063 28067
rect 22005 28027 22063 28033
rect 16724 27968 16813 27996
rect 16724 27956 16730 27968
rect 12437 27931 12495 27937
rect 12437 27928 12449 27931
rect 12308 27900 12449 27928
rect 12308 27888 12314 27900
rect 12437 27897 12449 27900
rect 12483 27897 12495 27931
rect 12437 27891 12495 27897
rect 16209 27931 16267 27937
rect 16209 27897 16221 27931
rect 16255 27897 16267 27931
rect 16209 27891 16267 27897
rect 7190 27820 7196 27872
rect 7248 27820 7254 27872
rect 13265 27863 13323 27869
rect 13265 27829 13277 27863
rect 13311 27860 13323 27863
rect 13446 27860 13452 27872
rect 13311 27832 13452 27860
rect 13311 27829 13323 27832
rect 13265 27823 13323 27829
rect 13446 27820 13452 27832
rect 13504 27820 13510 27872
rect 15286 27820 15292 27872
rect 15344 27820 15350 27872
rect 19794 27820 19800 27872
rect 19852 27820 19858 27872
rect 21082 27820 21088 27872
rect 21140 27820 21146 27872
rect 21269 27863 21327 27869
rect 21269 27829 21281 27863
rect 21315 27860 21327 27863
rect 21450 27860 21456 27872
rect 21315 27832 21456 27860
rect 21315 27829 21327 27832
rect 21269 27823 21327 27829
rect 21450 27820 21456 27832
rect 21508 27860 21514 27872
rect 21821 27863 21879 27869
rect 21821 27860 21833 27863
rect 21508 27832 21833 27860
rect 21508 27820 21514 27832
rect 21821 27829 21833 27832
rect 21867 27829 21879 27863
rect 21821 27823 21879 27829
rect 22278 27820 22284 27872
rect 22336 27860 22342 27872
rect 23842 27860 23848 27872
rect 22336 27832 23848 27860
rect 22336 27820 22342 27832
rect 23842 27820 23848 27832
rect 23900 27820 23906 27872
rect 1104 27770 34868 27792
rect 1104 27718 5170 27770
rect 5222 27718 5234 27770
rect 5286 27718 5298 27770
rect 5350 27718 5362 27770
rect 5414 27718 5426 27770
rect 5478 27718 13611 27770
rect 13663 27718 13675 27770
rect 13727 27718 13739 27770
rect 13791 27718 13803 27770
rect 13855 27718 13867 27770
rect 13919 27718 22052 27770
rect 22104 27718 22116 27770
rect 22168 27718 22180 27770
rect 22232 27718 22244 27770
rect 22296 27718 22308 27770
rect 22360 27718 30493 27770
rect 30545 27718 30557 27770
rect 30609 27718 30621 27770
rect 30673 27718 30685 27770
rect 30737 27718 30749 27770
rect 30801 27718 34868 27770
rect 1104 27696 34868 27718
rect 8757 27659 8815 27665
rect 8757 27625 8769 27659
rect 8803 27656 8815 27659
rect 9214 27656 9220 27668
rect 8803 27628 9220 27656
rect 8803 27625 8815 27628
rect 8757 27619 8815 27625
rect 9214 27616 9220 27628
rect 9272 27616 9278 27668
rect 10597 27659 10655 27665
rect 10597 27625 10609 27659
rect 10643 27656 10655 27659
rect 10870 27656 10876 27668
rect 10643 27628 10876 27656
rect 10643 27625 10655 27628
rect 10597 27619 10655 27625
rect 10870 27616 10876 27628
rect 10928 27616 10934 27668
rect 14182 27616 14188 27668
rect 14240 27616 14246 27668
rect 15930 27616 15936 27668
rect 15988 27616 15994 27668
rect 16022 27616 16028 27668
rect 16080 27616 16086 27668
rect 21266 27616 21272 27668
rect 21324 27656 21330 27668
rect 23014 27656 23020 27668
rect 21324 27628 23020 27656
rect 21324 27616 21330 27628
rect 23014 27616 23020 27628
rect 23072 27616 23078 27668
rect 19242 27548 19248 27600
rect 19300 27548 19306 27600
rect 19794 27548 19800 27600
rect 19852 27548 19858 27600
rect 20714 27548 20720 27600
rect 20772 27588 20778 27600
rect 20772 27560 21588 27588
rect 20772 27548 20778 27560
rect 12434 27480 12440 27532
rect 12492 27520 12498 27532
rect 13078 27520 13084 27532
rect 12492 27492 13084 27520
rect 12492 27480 12498 27492
rect 13078 27480 13084 27492
rect 13136 27480 13142 27532
rect 13817 27523 13875 27529
rect 13817 27489 13829 27523
rect 13863 27520 13875 27523
rect 14737 27523 14795 27529
rect 14737 27520 14749 27523
rect 13863 27492 14749 27520
rect 13863 27489 13875 27492
rect 13817 27483 13875 27489
rect 14737 27489 14749 27492
rect 14783 27489 14795 27523
rect 19812 27520 19840 27548
rect 14737 27483 14795 27489
rect 18892 27492 19840 27520
rect 20349 27523 20407 27529
rect 7190 27412 7196 27464
rect 7248 27412 7254 27464
rect 7374 27412 7380 27464
rect 7432 27452 7438 27464
rect 9217 27455 9275 27461
rect 9217 27452 9229 27455
rect 7432 27424 9229 27452
rect 7432 27412 7438 27424
rect 9217 27421 9229 27424
rect 9263 27452 9275 27455
rect 9858 27452 9864 27464
rect 9263 27424 9864 27452
rect 9263 27421 9275 27424
rect 9217 27415 9275 27421
rect 9858 27412 9864 27424
rect 9916 27412 9922 27464
rect 12161 27455 12219 27461
rect 12161 27421 12173 27455
rect 12207 27452 12219 27455
rect 12250 27452 12256 27464
rect 12207 27424 12256 27452
rect 12207 27421 12219 27424
rect 12161 27415 12219 27421
rect 12250 27412 12256 27424
rect 12308 27412 12314 27464
rect 12345 27455 12403 27461
rect 12345 27421 12357 27455
rect 12391 27452 12403 27455
rect 12526 27452 12532 27464
rect 12391 27424 12532 27452
rect 12391 27421 12403 27424
rect 12345 27415 12403 27421
rect 12526 27412 12532 27424
rect 12584 27412 12590 27464
rect 12894 27412 12900 27464
rect 12952 27412 12958 27464
rect 13725 27455 13783 27461
rect 13725 27421 13737 27455
rect 13771 27421 13783 27455
rect 13725 27415 13783 27421
rect 13909 27455 13967 27461
rect 13909 27421 13921 27455
rect 13955 27452 13967 27455
rect 14090 27452 14096 27464
rect 13955 27424 14096 27452
rect 13955 27421 13967 27424
rect 13909 27415 13967 27421
rect 7208 27384 7236 27412
rect 7622 27387 7680 27393
rect 7622 27384 7634 27387
rect 7208 27356 7634 27384
rect 7622 27353 7634 27356
rect 7668 27353 7680 27387
rect 7622 27347 7680 27353
rect 9484 27387 9542 27393
rect 9484 27353 9496 27387
rect 9530 27384 9542 27387
rect 9766 27384 9772 27396
rect 9530 27356 9772 27384
rect 9530 27353 9542 27356
rect 9484 27347 9542 27353
rect 9766 27344 9772 27356
rect 9824 27344 9830 27396
rect 13740 27384 13768 27415
rect 14090 27412 14096 27424
rect 14148 27412 14154 27464
rect 15286 27412 15292 27464
rect 15344 27452 15350 27464
rect 15381 27455 15439 27461
rect 15381 27452 15393 27455
rect 15344 27424 15393 27452
rect 15344 27412 15350 27424
rect 15381 27421 15393 27424
rect 15427 27421 15439 27455
rect 15657 27455 15715 27461
rect 15657 27452 15669 27455
rect 15381 27415 15439 27421
rect 15580 27424 15669 27452
rect 13740 27356 13952 27384
rect 13924 27328 13952 27356
rect 12253 27319 12311 27325
rect 12253 27285 12265 27319
rect 12299 27316 12311 27319
rect 12618 27316 12624 27328
rect 12299 27288 12624 27316
rect 12299 27285 12311 27288
rect 12253 27279 12311 27285
rect 12618 27276 12624 27288
rect 12676 27276 12682 27328
rect 13538 27276 13544 27328
rect 13596 27276 13602 27328
rect 13906 27276 13912 27328
rect 13964 27276 13970 27328
rect 14108 27316 14136 27412
rect 15580 27325 15608 27424
rect 15657 27421 15669 27424
rect 15703 27421 15715 27455
rect 15657 27415 15715 27421
rect 15746 27412 15752 27464
rect 15804 27452 15810 27464
rect 15933 27455 15991 27461
rect 15933 27452 15945 27455
rect 15804 27424 15945 27452
rect 15804 27412 15810 27424
rect 15933 27421 15945 27424
rect 15979 27421 15991 27455
rect 15933 27415 15991 27421
rect 17126 27412 17132 27464
rect 17184 27461 17190 27464
rect 17184 27452 17196 27461
rect 17405 27455 17463 27461
rect 17184 27424 17229 27452
rect 17184 27415 17196 27424
rect 17405 27421 17417 27455
rect 17451 27452 17463 27455
rect 17681 27455 17739 27461
rect 17681 27452 17693 27455
rect 17451 27424 17693 27452
rect 17451 27421 17463 27424
rect 17405 27415 17463 27421
rect 17681 27421 17693 27424
rect 17727 27452 17739 27455
rect 17770 27452 17776 27464
rect 17727 27424 17776 27452
rect 17727 27421 17739 27424
rect 17681 27415 17739 27421
rect 17184 27412 17190 27415
rect 17770 27412 17776 27424
rect 17828 27412 17834 27464
rect 17948 27455 18006 27461
rect 17948 27421 17960 27455
rect 17994 27452 18006 27455
rect 18892 27452 18920 27492
rect 20349 27489 20361 27523
rect 20395 27520 20407 27523
rect 20993 27523 21051 27529
rect 20993 27520 21005 27523
rect 20395 27492 21005 27520
rect 20395 27489 20407 27492
rect 20349 27483 20407 27489
rect 20993 27489 21005 27492
rect 21039 27489 21051 27523
rect 20993 27483 21051 27489
rect 21100 27492 21404 27520
rect 17994 27424 18920 27452
rect 19797 27455 19855 27461
rect 17994 27421 18006 27424
rect 17948 27415 18006 27421
rect 19797 27421 19809 27455
rect 19843 27421 19855 27455
rect 21100 27452 21128 27492
rect 19797 27415 19855 27421
rect 21008 27424 21128 27452
rect 15565 27319 15623 27325
rect 15565 27316 15577 27319
rect 14108 27288 15577 27316
rect 15565 27285 15577 27288
rect 15611 27285 15623 27319
rect 15565 27279 15623 27285
rect 15654 27276 15660 27328
rect 15712 27316 15718 27328
rect 15749 27319 15807 27325
rect 15749 27316 15761 27319
rect 15712 27288 15761 27316
rect 15712 27276 15718 27288
rect 15749 27285 15761 27288
rect 15795 27285 15807 27319
rect 15749 27279 15807 27285
rect 19058 27276 19064 27328
rect 19116 27316 19122 27328
rect 19812 27316 19840 27415
rect 21008 27328 21036 27424
rect 21174 27412 21180 27464
rect 21232 27452 21238 27464
rect 21376 27461 21404 27492
rect 21269 27455 21327 27461
rect 21269 27452 21281 27455
rect 21232 27424 21281 27452
rect 21232 27412 21238 27424
rect 21269 27421 21281 27424
rect 21315 27421 21327 27455
rect 21269 27415 21327 27421
rect 21361 27455 21419 27461
rect 21361 27421 21373 27455
rect 21407 27421 21419 27455
rect 21361 27415 21419 27421
rect 21474 27452 21532 27458
rect 21474 27418 21486 27452
rect 21520 27449 21532 27452
rect 21560 27449 21588 27560
rect 21726 27480 21732 27532
rect 21784 27480 21790 27532
rect 21520 27421 21588 27449
rect 21520 27418 21532 27421
rect 21474 27412 21532 27418
rect 21634 27412 21640 27464
rect 21692 27412 21698 27464
rect 22738 27412 22744 27464
rect 22796 27452 22802 27464
rect 22925 27455 22983 27461
rect 22925 27452 22937 27455
rect 22796 27424 22937 27452
rect 22796 27412 22802 27424
rect 22925 27421 22937 27424
rect 22971 27421 22983 27455
rect 22925 27415 22983 27421
rect 23109 27455 23167 27461
rect 23109 27421 23121 27455
rect 23155 27421 23167 27455
rect 23109 27415 23167 27421
rect 22646 27344 22652 27396
rect 22704 27384 22710 27396
rect 23124 27384 23152 27415
rect 23290 27412 23296 27464
rect 23348 27412 23354 27464
rect 25041 27455 25099 27461
rect 25041 27452 25053 27455
rect 24596 27424 25053 27452
rect 22704 27356 23152 27384
rect 22704 27344 22710 27356
rect 24596 27328 24624 27424
rect 25041 27421 25053 27424
rect 25087 27421 25099 27455
rect 25041 27415 25099 27421
rect 34514 27412 34520 27464
rect 34572 27412 34578 27464
rect 19116 27288 19840 27316
rect 19116 27276 19122 27288
rect 20898 27276 20904 27328
rect 20956 27276 20962 27328
rect 20990 27276 20996 27328
rect 21048 27276 21054 27328
rect 21174 27276 21180 27328
rect 21232 27316 21238 27328
rect 21910 27316 21916 27328
rect 21232 27288 21916 27316
rect 21232 27276 21238 27288
rect 21910 27276 21916 27288
rect 21968 27316 21974 27328
rect 22373 27319 22431 27325
rect 22373 27316 22385 27319
rect 21968 27288 22385 27316
rect 21968 27276 21974 27288
rect 22373 27285 22385 27288
rect 22419 27285 22431 27319
rect 22373 27279 22431 27285
rect 22922 27276 22928 27328
rect 22980 27276 22986 27328
rect 23934 27276 23940 27328
rect 23992 27276 23998 27328
rect 24578 27276 24584 27328
rect 24636 27276 24642 27328
rect 24854 27276 24860 27328
rect 24912 27276 24918 27328
rect 1104 27226 35027 27248
rect 1104 27174 9390 27226
rect 9442 27174 9454 27226
rect 9506 27174 9518 27226
rect 9570 27174 9582 27226
rect 9634 27174 9646 27226
rect 9698 27174 17831 27226
rect 17883 27174 17895 27226
rect 17947 27174 17959 27226
rect 18011 27174 18023 27226
rect 18075 27174 18087 27226
rect 18139 27174 26272 27226
rect 26324 27174 26336 27226
rect 26388 27174 26400 27226
rect 26452 27174 26464 27226
rect 26516 27174 26528 27226
rect 26580 27174 34713 27226
rect 34765 27174 34777 27226
rect 34829 27174 34841 27226
rect 34893 27174 34905 27226
rect 34957 27174 34969 27226
rect 35021 27174 35027 27226
rect 1104 27152 35027 27174
rect 8846 27072 8852 27124
rect 8904 27072 8910 27124
rect 9401 27115 9459 27121
rect 9401 27081 9413 27115
rect 9447 27112 9459 27115
rect 10042 27112 10048 27124
rect 9447 27084 10048 27112
rect 9447 27081 9459 27084
rect 9401 27075 9459 27081
rect 10042 27072 10048 27084
rect 10100 27072 10106 27124
rect 11974 27072 11980 27124
rect 12032 27112 12038 27124
rect 12434 27112 12440 27124
rect 12032 27084 12440 27112
rect 12032 27072 12038 27084
rect 12434 27072 12440 27084
rect 12492 27072 12498 27124
rect 12526 27072 12532 27124
rect 12584 27072 12590 27124
rect 13538 27072 13544 27124
rect 13596 27072 13602 27124
rect 13906 27072 13912 27124
rect 13964 27112 13970 27124
rect 16482 27112 16488 27124
rect 13964 27084 16488 27112
rect 13964 27072 13970 27084
rect 8864 27044 8892 27072
rect 8864 27016 9260 27044
rect 9030 26936 9036 26988
rect 9088 26936 9094 26988
rect 9232 26985 9260 27016
rect 11698 27004 11704 27056
rect 11756 27004 11762 27056
rect 12802 27004 12808 27056
rect 12860 27044 12866 27056
rect 13556 27044 13584 27072
rect 13826 27047 13884 27053
rect 13826 27044 13838 27047
rect 12860 27016 13492 27044
rect 13556 27016 13838 27044
rect 12860 27004 12866 27016
rect 9217 26979 9275 26985
rect 9217 26945 9229 26979
rect 9263 26945 9275 26979
rect 9217 26939 9275 26945
rect 11146 26936 11152 26988
rect 11204 26976 11210 26988
rect 11517 26979 11575 26985
rect 11517 26976 11529 26979
rect 11204 26948 11529 26976
rect 11204 26936 11210 26948
rect 11517 26945 11529 26948
rect 11563 26976 11575 26979
rect 11716 26976 11744 27004
rect 11563 26948 11744 26976
rect 11977 26979 12035 26985
rect 11563 26945 11575 26948
rect 11517 26939 11575 26945
rect 11977 26945 11989 26979
rect 12023 26976 12035 26979
rect 12158 26976 12164 26988
rect 12023 26948 12164 26976
rect 12023 26945 12035 26948
rect 11977 26939 12035 26945
rect 12158 26936 12164 26948
rect 12216 26936 12222 26988
rect 12345 26979 12403 26985
rect 12345 26945 12357 26979
rect 12391 26945 12403 26979
rect 13354 26976 13360 26988
rect 12345 26939 12403 26945
rect 13087 26948 13360 26976
rect 11701 26843 11759 26849
rect 11701 26809 11713 26843
rect 11747 26840 11759 26843
rect 12066 26840 12072 26852
rect 11747 26812 12072 26840
rect 11747 26809 11759 26812
rect 11701 26803 11759 26809
rect 12066 26800 12072 26812
rect 12124 26800 12130 26852
rect 12360 26840 12388 26939
rect 13087 26840 13115 26948
rect 13354 26936 13360 26948
rect 13412 26936 13418 26988
rect 13464 26976 13492 27016
rect 13826 27013 13838 27016
rect 13872 27013 13884 27047
rect 13826 27007 13884 27013
rect 13924 27016 14872 27044
rect 13924 26976 13952 27016
rect 13464 26948 13952 26976
rect 13998 26936 14004 26988
rect 14056 26976 14062 26988
rect 14844 26985 14872 27016
rect 15212 26985 15240 27084
rect 16482 27072 16488 27084
rect 16540 27072 16546 27124
rect 19794 27072 19800 27124
rect 19852 27112 19858 27124
rect 19889 27115 19947 27121
rect 19889 27112 19901 27115
rect 19852 27084 19901 27112
rect 19852 27072 19858 27084
rect 19889 27081 19901 27084
rect 19935 27081 19947 27115
rect 19889 27075 19947 27081
rect 20898 27072 20904 27124
rect 20956 27072 20962 27124
rect 21450 27072 21456 27124
rect 21508 27072 21514 27124
rect 21634 27072 21640 27124
rect 21692 27072 21698 27124
rect 22373 27115 22431 27121
rect 22373 27081 22385 27115
rect 22419 27112 22431 27115
rect 22646 27112 22652 27124
rect 22419 27084 22652 27112
rect 22419 27081 22431 27084
rect 22373 27075 22431 27081
rect 22646 27072 22652 27084
rect 22704 27072 22710 27124
rect 22922 27072 22928 27124
rect 22980 27072 22986 27124
rect 23109 27115 23167 27121
rect 23109 27081 23121 27115
rect 23155 27112 23167 27115
rect 23290 27112 23296 27124
rect 23155 27084 23296 27112
rect 23155 27081 23167 27084
rect 23109 27075 23167 27081
rect 23290 27072 23296 27084
rect 23348 27072 23354 27124
rect 23934 27072 23940 27124
rect 23992 27072 23998 27124
rect 15470 27004 15476 27056
rect 15528 27004 15534 27056
rect 16853 27047 16911 27053
rect 16853 27044 16865 27047
rect 15764 27016 16865 27044
rect 14093 26979 14151 26985
rect 14093 26976 14105 26979
rect 14056 26948 14105 26976
rect 14056 26936 14062 26948
rect 14093 26945 14105 26948
rect 14139 26945 14151 26979
rect 14093 26939 14151 26945
rect 14829 26979 14887 26985
rect 14829 26945 14841 26979
rect 14875 26945 14887 26979
rect 15105 26979 15163 26985
rect 15105 26976 15117 26979
rect 14829 26939 14887 26945
rect 15028 26948 15117 26976
rect 15028 26852 15056 26948
rect 15105 26945 15117 26948
rect 15151 26945 15163 26979
rect 15105 26939 15163 26945
rect 15197 26979 15255 26985
rect 15197 26945 15209 26979
rect 15243 26945 15255 26979
rect 15197 26939 15255 26945
rect 15381 26979 15439 26985
rect 15381 26945 15393 26979
rect 15427 26945 15439 26979
rect 15381 26939 15439 26945
rect 12360 26812 13115 26840
rect 15010 26800 15016 26852
rect 15068 26800 15074 26852
rect 15396 26840 15424 26939
rect 15488 26917 15516 27004
rect 15654 26936 15660 26988
rect 15712 26976 15718 26988
rect 15764 26985 15792 27016
rect 16853 27013 16865 27016
rect 16899 27044 16911 27047
rect 17402 27044 17408 27056
rect 16899 27016 17408 27044
rect 16899 27013 16911 27016
rect 16853 27007 16911 27013
rect 17402 27004 17408 27016
rect 17460 27004 17466 27056
rect 15749 26979 15807 26985
rect 15749 26976 15761 26979
rect 15712 26948 15761 26976
rect 15712 26936 15718 26948
rect 15749 26945 15761 26948
rect 15795 26945 15807 26979
rect 15749 26939 15807 26945
rect 16761 26979 16819 26985
rect 16761 26945 16773 26979
rect 16807 26945 16819 26979
rect 16761 26939 16819 26945
rect 17037 26979 17095 26985
rect 17037 26945 17049 26979
rect 17083 26976 17095 26979
rect 18782 26976 18788 26988
rect 17083 26948 18788 26976
rect 17083 26945 17095 26948
rect 17037 26939 17095 26945
rect 15473 26911 15531 26917
rect 15473 26877 15485 26911
rect 15519 26877 15531 26911
rect 15473 26871 15531 26877
rect 15930 26868 15936 26920
rect 15988 26908 15994 26920
rect 16393 26911 16451 26917
rect 16393 26908 16405 26911
rect 15988 26880 16405 26908
rect 15988 26868 15994 26880
rect 16393 26877 16405 26880
rect 16439 26877 16451 26911
rect 16393 26871 16451 26877
rect 16776 26840 16804 26939
rect 18782 26936 18788 26948
rect 18840 26936 18846 26988
rect 19812 26985 19840 27072
rect 20916 27044 20944 27072
rect 21002 27047 21060 27053
rect 21002 27044 21014 27047
rect 20916 27016 21014 27044
rect 21002 27013 21014 27016
rect 21048 27013 21060 27047
rect 21002 27007 21060 27013
rect 21358 27004 21364 27056
rect 21416 27004 21422 27056
rect 21652 27044 21680 27072
rect 22940 27044 22968 27072
rect 21652 27016 22508 27044
rect 21364 27001 21422 27004
rect 19797 26979 19855 26985
rect 19797 26945 19809 26979
rect 19843 26945 19855 26979
rect 19797 26939 19855 26945
rect 21266 26936 21272 26988
rect 21324 26936 21330 26988
rect 21364 26967 21376 27001
rect 21410 26967 21422 27001
rect 21364 26961 21422 26967
rect 21542 26936 21548 26988
rect 21600 26976 21606 26988
rect 22480 26985 22508 27016
rect 22664 27016 22968 27044
rect 22664 26985 22692 27016
rect 23198 27004 23204 27056
rect 23256 27004 23262 27056
rect 23468 27047 23526 27053
rect 23468 27013 23480 27047
rect 23514 27044 23526 27047
rect 23952 27044 23980 27072
rect 23514 27016 23980 27044
rect 23514 27013 23526 27016
rect 23468 27007 23526 27013
rect 21637 26979 21695 26985
rect 22083 26979 22141 26985
rect 21637 26976 21649 26979
rect 21600 26948 21649 26976
rect 21600 26936 21606 26948
rect 21637 26945 21649 26948
rect 21683 26945 21695 26979
rect 21928 26976 22095 26979
rect 21637 26939 21695 26945
rect 21836 26951 22095 26976
rect 21836 26948 21956 26951
rect 17126 26868 17132 26920
rect 17184 26868 17190 26920
rect 18414 26868 18420 26920
rect 18472 26868 18478 26920
rect 19429 26911 19487 26917
rect 19429 26877 19441 26911
rect 19475 26908 19487 26911
rect 19610 26908 19616 26920
rect 19475 26880 19616 26908
rect 19475 26877 19487 26880
rect 19429 26871 19487 26877
rect 19610 26868 19616 26880
rect 19668 26868 19674 26920
rect 15396 26812 16804 26840
rect 15764 26784 15792 26812
rect 17586 26800 17592 26852
rect 17644 26840 17650 26852
rect 17865 26843 17923 26849
rect 17865 26840 17877 26843
rect 17644 26812 17877 26840
rect 17644 26800 17650 26812
rect 17865 26809 17877 26812
rect 17911 26809 17923 26843
rect 17865 26803 17923 26809
rect 21836 26784 21864 26948
rect 22083 26945 22095 26951
rect 22129 26945 22141 26979
rect 22083 26939 22141 26945
rect 22465 26979 22523 26985
rect 22465 26945 22477 26979
rect 22511 26976 22523 26979
rect 22649 26979 22707 26985
rect 22511 26948 22600 26976
rect 22511 26945 22523 26948
rect 22465 26939 22523 26945
rect 22005 26911 22063 26917
rect 22005 26877 22017 26911
rect 22051 26908 22063 26911
rect 22051 26880 22140 26908
rect 22051 26877 22063 26880
rect 22005 26871 22063 26877
rect 22112 26840 22140 26880
rect 22278 26840 22284 26852
rect 22112 26812 22284 26840
rect 22278 26800 22284 26812
rect 22336 26800 22342 26852
rect 11606 26732 11612 26784
rect 11664 26732 11670 26784
rect 11839 26775 11897 26781
rect 11839 26741 11851 26775
rect 11885 26772 11897 26775
rect 12618 26772 12624 26784
rect 11885 26744 12624 26772
rect 11885 26741 11897 26744
rect 11839 26735 11897 26741
rect 12618 26732 12624 26744
rect 12676 26732 12682 26784
rect 12713 26775 12771 26781
rect 12713 26741 12725 26775
rect 12759 26772 12771 26775
rect 12802 26772 12808 26784
rect 12759 26744 12808 26772
rect 12759 26741 12771 26744
rect 12713 26735 12771 26741
rect 12802 26732 12808 26744
rect 12860 26732 12866 26784
rect 12986 26732 12992 26784
rect 13044 26772 13050 26784
rect 14645 26775 14703 26781
rect 14645 26772 14657 26775
rect 13044 26744 14657 26772
rect 13044 26732 13050 26744
rect 14645 26741 14657 26744
rect 14691 26741 14703 26775
rect 14645 26735 14703 26741
rect 14921 26775 14979 26781
rect 14921 26741 14933 26775
rect 14967 26772 14979 26775
rect 15102 26772 15108 26784
rect 14967 26744 15108 26772
rect 14967 26741 14979 26744
rect 14921 26735 14979 26741
rect 15102 26732 15108 26744
rect 15160 26732 15166 26784
rect 15378 26732 15384 26784
rect 15436 26732 15442 26784
rect 15562 26732 15568 26784
rect 15620 26732 15626 26784
rect 15657 26775 15715 26781
rect 15657 26741 15669 26775
rect 15703 26772 15715 26775
rect 15746 26772 15752 26784
rect 15703 26744 15752 26772
rect 15703 26741 15715 26744
rect 15657 26735 15715 26741
rect 15746 26732 15752 26744
rect 15804 26732 15810 26784
rect 15838 26732 15844 26784
rect 15896 26732 15902 26784
rect 17034 26732 17040 26784
rect 17092 26732 17098 26784
rect 17770 26732 17776 26784
rect 17828 26732 17834 26784
rect 19702 26732 19708 26784
rect 19760 26732 19766 26784
rect 21634 26732 21640 26784
rect 21692 26732 21698 26784
rect 21818 26732 21824 26784
rect 21876 26732 21882 26784
rect 22462 26732 22468 26784
rect 22520 26772 22526 26784
rect 22572 26772 22600 26948
rect 22649 26945 22661 26979
rect 22695 26945 22707 26979
rect 22649 26939 22707 26945
rect 22738 26936 22744 26988
rect 22796 26936 22802 26988
rect 22833 26979 22891 26985
rect 22833 26945 22845 26979
rect 22879 26976 22891 26979
rect 23216 26976 23244 27004
rect 24854 26976 24860 26988
rect 22879 26948 24860 26976
rect 22879 26945 22891 26948
rect 22833 26939 22891 26945
rect 24854 26936 24860 26948
rect 24912 26936 24918 26988
rect 23014 26868 23020 26920
rect 23072 26908 23078 26920
rect 23201 26911 23259 26917
rect 23201 26908 23213 26911
rect 23072 26880 23213 26908
rect 23072 26868 23078 26880
rect 23201 26877 23213 26880
rect 23247 26877 23259 26911
rect 23201 26871 23259 26877
rect 22520 26744 22600 26772
rect 22520 26732 22526 26744
rect 24578 26732 24584 26784
rect 24636 26732 24642 26784
rect 1104 26682 34868 26704
rect 1104 26630 5170 26682
rect 5222 26630 5234 26682
rect 5286 26630 5298 26682
rect 5350 26630 5362 26682
rect 5414 26630 5426 26682
rect 5478 26630 13611 26682
rect 13663 26630 13675 26682
rect 13727 26630 13739 26682
rect 13791 26630 13803 26682
rect 13855 26630 13867 26682
rect 13919 26630 22052 26682
rect 22104 26630 22116 26682
rect 22168 26630 22180 26682
rect 22232 26630 22244 26682
rect 22296 26630 22308 26682
rect 22360 26630 30493 26682
rect 30545 26630 30557 26682
rect 30609 26630 30621 26682
rect 30673 26630 30685 26682
rect 30737 26630 30749 26682
rect 30801 26630 34868 26682
rect 1104 26608 34868 26630
rect 11606 26528 11612 26580
rect 11664 26528 11670 26580
rect 12713 26571 12771 26577
rect 12713 26537 12725 26571
rect 12759 26568 12771 26571
rect 12894 26568 12900 26580
rect 12759 26540 12900 26568
rect 12759 26537 12771 26540
rect 12713 26531 12771 26537
rect 12894 26528 12900 26540
rect 12952 26528 12958 26580
rect 13541 26571 13599 26577
rect 13541 26568 13553 26571
rect 13004 26540 13553 26568
rect 11624 26432 11652 26528
rect 11701 26435 11759 26441
rect 11701 26432 11713 26435
rect 11624 26404 11713 26432
rect 11701 26401 11713 26404
rect 11747 26401 11759 26435
rect 11701 26395 11759 26401
rect 12066 26392 12072 26444
rect 12124 26392 12130 26444
rect 12158 26392 12164 26444
rect 12216 26432 12222 26444
rect 12529 26435 12587 26441
rect 12529 26432 12541 26435
rect 12216 26404 12541 26432
rect 12216 26392 12222 26404
rect 8294 26324 8300 26376
rect 8352 26364 8358 26376
rect 9769 26367 9827 26373
rect 9769 26364 9781 26367
rect 8352 26336 9781 26364
rect 8352 26324 8358 26336
rect 9769 26333 9781 26336
rect 9815 26364 9827 26367
rect 9858 26364 9864 26376
rect 9815 26336 9864 26364
rect 9815 26333 9827 26336
rect 9769 26327 9827 26333
rect 9858 26324 9864 26336
rect 9916 26324 9922 26376
rect 11330 26324 11336 26376
rect 11388 26364 11394 26376
rect 11425 26367 11483 26373
rect 11425 26364 11437 26367
rect 11388 26336 11437 26364
rect 11388 26324 11394 26336
rect 11425 26333 11437 26336
rect 11471 26333 11483 26367
rect 11425 26327 11483 26333
rect 11609 26367 11667 26373
rect 11609 26333 11621 26367
rect 11655 26333 11667 26367
rect 11609 26327 11667 26333
rect 11793 26367 11851 26373
rect 11793 26333 11805 26367
rect 11839 26333 11851 26367
rect 11793 26327 11851 26333
rect 10036 26299 10094 26305
rect 10036 26265 10048 26299
rect 10082 26296 10094 26299
rect 10686 26296 10692 26308
rect 10082 26268 10692 26296
rect 10082 26265 10094 26268
rect 10036 26259 10094 26265
rect 10686 26256 10692 26268
rect 10744 26256 10750 26308
rect 11624 26296 11652 26327
rect 11808 26296 11836 26327
rect 11974 26324 11980 26376
rect 12032 26324 12038 26376
rect 12084 26364 12112 26392
rect 12360 26376 12388 26404
rect 12529 26401 12541 26404
rect 12575 26401 12587 26435
rect 12529 26395 12587 26401
rect 12618 26392 12624 26444
rect 12676 26432 12682 26444
rect 13004 26432 13032 26540
rect 13541 26537 13553 26540
rect 13587 26537 13599 26571
rect 13541 26531 13599 26537
rect 17126 26528 17132 26580
rect 17184 26528 17190 26580
rect 19702 26528 19708 26580
rect 19760 26528 19766 26580
rect 20533 26571 20591 26577
rect 20533 26537 20545 26571
rect 20579 26568 20591 26571
rect 21082 26568 21088 26580
rect 20579 26540 21088 26568
rect 20579 26537 20591 26540
rect 20533 26531 20591 26537
rect 21082 26528 21088 26540
rect 21140 26528 21146 26580
rect 21634 26528 21640 26580
rect 21692 26528 21698 26580
rect 22370 26528 22376 26580
rect 22428 26568 22434 26580
rect 22741 26571 22799 26577
rect 22741 26568 22753 26571
rect 22428 26540 22753 26568
rect 22428 26528 22434 26540
rect 22741 26537 22753 26540
rect 22787 26568 22799 26571
rect 23385 26571 23443 26577
rect 23385 26568 23397 26571
rect 22787 26540 23397 26568
rect 22787 26537 22799 26540
rect 22741 26531 22799 26537
rect 23385 26537 23397 26540
rect 23431 26537 23443 26571
rect 23385 26531 23443 26537
rect 14737 26503 14795 26509
rect 12676 26404 13032 26432
rect 13372 26472 13952 26500
rect 12676 26392 12682 26404
rect 12253 26367 12311 26373
rect 12253 26364 12265 26367
rect 12084 26336 12265 26364
rect 12253 26333 12265 26336
rect 12299 26333 12311 26367
rect 12253 26327 12311 26333
rect 12342 26324 12348 26376
rect 12400 26324 12406 26376
rect 12437 26367 12495 26373
rect 12437 26333 12449 26367
rect 12483 26364 12495 26367
rect 12728 26364 12756 26404
rect 12483 26336 12756 26364
rect 12483 26333 12495 26336
rect 12437 26327 12495 26333
rect 12986 26324 12992 26376
rect 13044 26324 13050 26376
rect 13372 26373 13400 26472
rect 13725 26435 13783 26441
rect 13725 26401 13737 26435
rect 13771 26432 13783 26435
rect 13924 26432 13952 26472
rect 14737 26469 14749 26503
rect 14783 26500 14795 26503
rect 15010 26500 15016 26512
rect 14783 26472 15016 26500
rect 14783 26469 14795 26472
rect 14737 26463 14795 26469
rect 15010 26460 15016 26472
rect 15068 26460 15074 26512
rect 19061 26503 19119 26509
rect 19061 26469 19073 26503
rect 19107 26500 19119 26503
rect 19337 26503 19395 26509
rect 19337 26500 19349 26503
rect 19107 26472 19349 26500
rect 19107 26469 19119 26472
rect 19061 26463 19119 26469
rect 19337 26469 19349 26472
rect 19383 26500 19395 26503
rect 19610 26500 19616 26512
rect 19383 26472 19616 26500
rect 19383 26469 19395 26472
rect 19337 26463 19395 26469
rect 19610 26460 19616 26472
rect 19668 26460 19674 26512
rect 16117 26435 16175 26441
rect 13771 26404 13860 26432
rect 13924 26404 14872 26432
rect 13771 26401 13783 26404
rect 13725 26395 13783 26401
rect 13081 26367 13139 26373
rect 13081 26333 13093 26367
rect 13127 26333 13139 26367
rect 13081 26327 13139 26333
rect 13173 26367 13231 26373
rect 13173 26333 13185 26367
rect 13219 26364 13231 26367
rect 13357 26367 13415 26373
rect 13219 26336 13308 26364
rect 13219 26333 13231 26336
rect 13173 26327 13231 26333
rect 12069 26299 12127 26305
rect 12069 26296 12081 26299
rect 11164 26268 11468 26296
rect 11624 26268 11744 26296
rect 11808 26268 12081 26296
rect 11164 26237 11192 26268
rect 11149 26231 11207 26237
rect 11149 26197 11161 26231
rect 11195 26197 11207 26231
rect 11149 26191 11207 26197
rect 11238 26188 11244 26240
rect 11296 26188 11302 26240
rect 11440 26228 11468 26268
rect 11606 26228 11612 26240
rect 11440 26200 11612 26228
rect 11606 26188 11612 26200
rect 11664 26188 11670 26240
rect 11716 26228 11744 26268
rect 12069 26265 12081 26268
rect 12115 26265 12127 26299
rect 12069 26259 12127 26265
rect 11790 26228 11796 26240
rect 11716 26200 11796 26228
rect 11790 26188 11796 26200
rect 11848 26228 11854 26240
rect 13096 26228 13124 26327
rect 13280 26296 13308 26336
rect 13357 26333 13369 26367
rect 13403 26333 13415 26367
rect 13357 26327 13415 26333
rect 13446 26324 13452 26376
rect 13504 26324 13510 26376
rect 13725 26299 13783 26305
rect 13725 26296 13737 26299
rect 13280 26268 13737 26296
rect 13725 26265 13737 26268
rect 13771 26265 13783 26299
rect 13725 26259 13783 26265
rect 13832 26228 13860 26404
rect 14274 26324 14280 26376
rect 14332 26364 14338 26376
rect 14642 26364 14648 26376
rect 14332 26336 14648 26364
rect 14332 26324 14338 26336
rect 14642 26324 14648 26336
rect 14700 26324 14706 26376
rect 14844 26308 14872 26404
rect 16117 26401 16129 26435
rect 16163 26432 16175 26435
rect 16666 26432 16672 26444
rect 16163 26404 16672 26432
rect 16163 26401 16175 26404
rect 16117 26395 16175 26401
rect 16666 26392 16672 26404
rect 16724 26432 16730 26444
rect 17678 26432 17684 26444
rect 16724 26404 17684 26432
rect 16724 26392 16730 26404
rect 17678 26392 17684 26404
rect 17736 26392 17742 26444
rect 19720 26432 19748 26528
rect 21652 26500 21680 26528
rect 23198 26500 23204 26512
rect 20456 26472 21680 26500
rect 22388 26472 23204 26500
rect 19536 26404 20024 26432
rect 15838 26324 15844 26376
rect 15896 26373 15902 26376
rect 15896 26364 15908 26373
rect 15896 26336 15941 26364
rect 15896 26327 15908 26336
rect 15896 26324 15902 26327
rect 16390 26324 16396 26376
rect 16448 26324 16454 26376
rect 17034 26324 17040 26376
rect 17092 26364 17098 26376
rect 17129 26367 17187 26373
rect 17129 26364 17141 26367
rect 17092 26336 17141 26364
rect 17092 26324 17098 26336
rect 17129 26333 17141 26336
rect 17175 26333 17187 26367
rect 17129 26327 17187 26333
rect 17221 26367 17279 26373
rect 17221 26333 17233 26367
rect 17267 26364 17279 26367
rect 17267 26336 17724 26364
rect 17267 26333 17279 26336
rect 17221 26327 17279 26333
rect 14826 26256 14832 26308
rect 14884 26296 14890 26308
rect 14884 26268 15424 26296
rect 14884 26256 14890 26268
rect 14461 26231 14519 26237
rect 14461 26228 14473 26231
rect 11848 26200 14473 26228
rect 11848 26188 11854 26200
rect 14461 26197 14473 26200
rect 14507 26228 14519 26231
rect 15194 26228 15200 26240
rect 14507 26200 15200 26228
rect 14507 26197 14519 26200
rect 14461 26191 14519 26197
rect 15194 26188 15200 26200
rect 15252 26188 15258 26240
rect 15396 26228 15424 26268
rect 16482 26256 16488 26308
rect 16540 26296 16546 26308
rect 17405 26299 17463 26305
rect 17405 26296 17417 26299
rect 16540 26268 17417 26296
rect 16540 26256 16546 26268
rect 17144 26240 17172 26268
rect 17405 26265 17417 26268
rect 17451 26265 17463 26299
rect 17696 26296 17724 26336
rect 17770 26324 17776 26376
rect 17828 26364 17834 26376
rect 17937 26367 17995 26373
rect 17937 26364 17949 26367
rect 17828 26336 17949 26364
rect 17828 26324 17834 26336
rect 17937 26333 17949 26336
rect 17983 26333 17995 26367
rect 17937 26327 17995 26333
rect 18414 26324 18420 26376
rect 18472 26324 18478 26376
rect 19245 26367 19303 26373
rect 19245 26333 19257 26367
rect 19291 26364 19303 26367
rect 19426 26364 19432 26376
rect 19291 26336 19432 26364
rect 19291 26333 19303 26336
rect 19245 26327 19303 26333
rect 19426 26324 19432 26336
rect 19484 26324 19490 26376
rect 19536 26373 19564 26404
rect 19996 26373 20024 26404
rect 20456 26373 20484 26472
rect 20717 26435 20775 26441
rect 20717 26401 20729 26435
rect 20763 26432 20775 26435
rect 20763 26404 20944 26432
rect 20763 26401 20775 26404
rect 20717 26395 20775 26401
rect 19521 26367 19579 26373
rect 19521 26333 19533 26367
rect 19567 26333 19579 26367
rect 19521 26327 19579 26333
rect 19613 26367 19671 26373
rect 19613 26333 19625 26367
rect 19659 26364 19671 26367
rect 19889 26367 19947 26373
rect 19889 26364 19901 26367
rect 19659 26336 19901 26364
rect 19659 26333 19671 26336
rect 19613 26327 19671 26333
rect 19889 26333 19901 26336
rect 19935 26333 19947 26367
rect 19889 26327 19947 26333
rect 19981 26367 20039 26373
rect 19981 26333 19993 26367
rect 20027 26333 20039 26367
rect 19981 26327 20039 26333
rect 20165 26367 20223 26373
rect 20165 26333 20177 26367
rect 20211 26333 20223 26367
rect 20165 26327 20223 26333
rect 20441 26367 20499 26373
rect 20441 26333 20453 26367
rect 20487 26333 20499 26367
rect 20441 26327 20499 26333
rect 18432 26296 18460 26324
rect 19628 26296 19656 26327
rect 17696 26268 18368 26296
rect 18432 26268 19656 26296
rect 17405 26259 17463 26265
rect 15470 26228 15476 26240
rect 15396 26200 15476 26228
rect 15470 26188 15476 26200
rect 15528 26188 15534 26240
rect 16942 26188 16948 26240
rect 17000 26228 17006 26240
rect 17037 26231 17095 26237
rect 17037 26228 17049 26231
rect 17000 26200 17049 26228
rect 17000 26188 17006 26200
rect 17037 26197 17049 26200
rect 17083 26197 17095 26231
rect 17037 26191 17095 26197
rect 17126 26188 17132 26240
rect 17184 26188 17190 26240
rect 18340 26228 18368 26268
rect 19702 26256 19708 26308
rect 19760 26296 19766 26308
rect 20180 26296 20208 26327
rect 19760 26268 20208 26296
rect 19760 26256 19766 26268
rect 20714 26256 20720 26308
rect 20772 26256 20778 26308
rect 20809 26299 20867 26305
rect 20809 26265 20821 26299
rect 20855 26265 20867 26299
rect 20916 26296 20944 26404
rect 21450 26392 21456 26444
rect 21508 26392 21514 26444
rect 22094 26392 22100 26444
rect 22152 26432 22158 26444
rect 22388 26432 22416 26472
rect 23198 26460 23204 26472
rect 23256 26460 23262 26512
rect 22925 26435 22983 26441
rect 22152 26404 22416 26432
rect 22152 26392 22158 26404
rect 21361 26367 21419 26373
rect 21361 26333 21373 26367
rect 21407 26364 21419 26367
rect 21542 26364 21548 26376
rect 21407 26336 21548 26364
rect 21407 26333 21419 26336
rect 21361 26327 21419 26333
rect 21542 26324 21548 26336
rect 21600 26324 21606 26376
rect 21726 26324 21732 26376
rect 21784 26364 21790 26376
rect 22388 26373 22416 26404
rect 22480 26404 22784 26432
rect 22005 26367 22063 26373
rect 22005 26364 22017 26367
rect 21784 26336 22017 26364
rect 21784 26324 21790 26336
rect 22005 26333 22017 26336
rect 22051 26364 22063 26367
rect 22189 26367 22247 26373
rect 22189 26364 22201 26367
rect 22051 26336 22201 26364
rect 22051 26333 22063 26336
rect 22005 26327 22063 26333
rect 22189 26333 22201 26336
rect 22235 26333 22247 26367
rect 22189 26327 22247 26333
rect 22373 26367 22431 26373
rect 22373 26333 22385 26367
rect 22419 26333 22431 26367
rect 22373 26327 22431 26333
rect 20990 26296 20996 26308
rect 20916 26268 20996 26296
rect 20809 26259 20867 26265
rect 18598 26228 18604 26240
rect 18340 26200 18604 26228
rect 18598 26188 18604 26200
rect 18656 26188 18662 26240
rect 19794 26188 19800 26240
rect 19852 26188 19858 26240
rect 20346 26188 20352 26240
rect 20404 26188 20410 26240
rect 20824 26228 20852 26259
rect 20990 26256 20996 26268
rect 21048 26256 21054 26308
rect 21085 26299 21143 26305
rect 21085 26265 21097 26299
rect 21131 26296 21143 26299
rect 21818 26296 21824 26308
rect 21131 26268 21824 26296
rect 21131 26265 21143 26268
rect 21085 26259 21143 26265
rect 21818 26256 21824 26268
rect 21876 26256 21882 26308
rect 20898 26228 20904 26240
rect 20824 26200 20904 26228
rect 20898 26188 20904 26200
rect 20956 26228 20962 26240
rect 21358 26228 21364 26240
rect 20956 26200 21364 26228
rect 20956 26188 20962 26200
rect 21358 26188 21364 26200
rect 21416 26188 21422 26240
rect 21910 26188 21916 26240
rect 21968 26228 21974 26240
rect 22480 26228 22508 26404
rect 22646 26324 22652 26376
rect 22704 26324 22710 26376
rect 22756 26364 22784 26404
rect 22925 26401 22937 26435
rect 22971 26432 22983 26435
rect 23109 26435 23167 26441
rect 23109 26432 23121 26435
rect 22971 26404 23121 26432
rect 22971 26401 22983 26404
rect 22925 26395 22983 26401
rect 23109 26401 23121 26404
rect 23155 26432 23167 26435
rect 23155 26404 23520 26432
rect 23155 26401 23167 26404
rect 23109 26395 23167 26401
rect 23017 26367 23075 26373
rect 23017 26364 23029 26367
rect 22756 26336 23029 26364
rect 23017 26333 23029 26336
rect 23063 26333 23075 26367
rect 23017 26327 23075 26333
rect 23198 26324 23204 26376
rect 23256 26324 23262 26376
rect 23492 26373 23520 26404
rect 23293 26367 23351 26373
rect 23293 26333 23305 26367
rect 23339 26333 23351 26367
rect 23293 26327 23351 26333
rect 23477 26367 23535 26373
rect 23477 26333 23489 26367
rect 23523 26333 23535 26367
rect 23477 26327 23535 26333
rect 22557 26299 22615 26305
rect 22557 26265 22569 26299
rect 22603 26296 22615 26299
rect 23308 26296 23336 26327
rect 22603 26268 23336 26296
rect 22603 26265 22615 26268
rect 22557 26259 22615 26265
rect 21968 26200 22508 26228
rect 22925 26231 22983 26237
rect 21968 26188 21974 26200
rect 22925 26197 22937 26231
rect 22971 26228 22983 26231
rect 23106 26228 23112 26240
rect 22971 26200 23112 26228
rect 22971 26197 22983 26200
rect 22925 26191 22983 26197
rect 23106 26188 23112 26200
rect 23164 26188 23170 26240
rect 1104 26138 35027 26160
rect 1104 26086 9390 26138
rect 9442 26086 9454 26138
rect 9506 26086 9518 26138
rect 9570 26086 9582 26138
rect 9634 26086 9646 26138
rect 9698 26086 17831 26138
rect 17883 26086 17895 26138
rect 17947 26086 17959 26138
rect 18011 26086 18023 26138
rect 18075 26086 18087 26138
rect 18139 26086 26272 26138
rect 26324 26086 26336 26138
rect 26388 26086 26400 26138
rect 26452 26086 26464 26138
rect 26516 26086 26528 26138
rect 26580 26086 34713 26138
rect 34765 26086 34777 26138
rect 34829 26086 34841 26138
rect 34893 26086 34905 26138
rect 34957 26086 34969 26138
rect 35021 26086 35027 26138
rect 1104 26064 35027 26086
rect 8294 25984 8300 26036
rect 8352 25984 8358 26036
rect 21266 26024 21272 26036
rect 10428 25996 18276 26024
rect 10428 25900 10456 25996
rect 10686 25916 10692 25968
rect 10744 25916 10750 25968
rect 12342 25916 12348 25968
rect 12400 25956 12406 25968
rect 12897 25959 12955 25965
rect 12897 25956 12909 25959
rect 12400 25928 12909 25956
rect 12400 25916 12406 25928
rect 12897 25925 12909 25928
rect 12943 25925 12955 25959
rect 12897 25919 12955 25925
rect 13262 25916 13268 25968
rect 13320 25956 13326 25968
rect 14826 25956 14832 25968
rect 13320 25928 14320 25956
rect 13320 25916 13326 25928
rect 9585 25891 9643 25897
rect 9585 25857 9597 25891
rect 9631 25888 9643 25891
rect 10410 25888 10416 25900
rect 9631 25860 10416 25888
rect 9631 25857 9643 25860
rect 9585 25851 9643 25857
rect 10410 25848 10416 25860
rect 10468 25848 10474 25900
rect 11238 25848 11244 25900
rect 11296 25848 11302 25900
rect 11517 25891 11575 25897
rect 11517 25857 11529 25891
rect 11563 25888 11575 25891
rect 11606 25888 11612 25900
rect 11563 25860 11612 25888
rect 11563 25857 11575 25860
rect 11517 25851 11575 25857
rect 11606 25848 11612 25860
rect 11664 25848 11670 25900
rect 12434 25848 12440 25900
rect 12492 25848 12498 25900
rect 12618 25848 12624 25900
rect 12676 25848 12682 25900
rect 12710 25848 12716 25900
rect 12768 25848 12774 25900
rect 12986 25848 12992 25900
rect 13044 25848 13050 25900
rect 13081 25891 13139 25897
rect 13081 25857 13093 25891
rect 13127 25888 13139 25891
rect 13170 25888 13176 25900
rect 13127 25860 13176 25888
rect 13127 25857 13139 25860
rect 13081 25851 13139 25857
rect 13170 25848 13176 25860
rect 13228 25848 13234 25900
rect 13538 25848 13544 25900
rect 13596 25888 13602 25900
rect 14182 25888 14188 25900
rect 13596 25860 14188 25888
rect 13596 25848 13602 25860
rect 14182 25848 14188 25860
rect 14240 25848 14246 25900
rect 14292 25897 14320 25928
rect 14752 25928 14832 25956
rect 14752 25897 14780 25928
rect 14826 25916 14832 25928
rect 14884 25916 14890 25968
rect 15194 25956 15200 25968
rect 15028 25928 15200 25956
rect 15028 25897 15056 25928
rect 15194 25916 15200 25928
rect 15252 25916 15258 25968
rect 15473 25959 15531 25965
rect 15473 25925 15485 25959
rect 15519 25956 15531 25959
rect 15562 25956 15568 25968
rect 15519 25928 15568 25956
rect 15519 25925 15531 25928
rect 15473 25919 15531 25925
rect 15562 25916 15568 25928
rect 15620 25916 15626 25968
rect 15654 25916 15660 25968
rect 15712 25916 15718 25968
rect 14277 25891 14335 25897
rect 14277 25857 14289 25891
rect 14323 25857 14335 25891
rect 14277 25851 14335 25857
rect 14737 25891 14795 25897
rect 14737 25857 14749 25891
rect 14783 25857 14795 25891
rect 14737 25851 14795 25857
rect 14921 25891 14979 25897
rect 14921 25857 14933 25891
rect 14967 25857 14979 25891
rect 14921 25851 14979 25857
rect 15013 25891 15071 25897
rect 15013 25857 15025 25891
rect 15059 25857 15071 25891
rect 15013 25851 15071 25857
rect 12529 25823 12587 25829
rect 12529 25789 12541 25823
rect 12575 25820 12587 25823
rect 12636 25820 12664 25848
rect 12575 25792 12664 25820
rect 13004 25820 13032 25848
rect 13265 25823 13323 25829
rect 13265 25820 13277 25823
rect 13004 25792 13277 25820
rect 12575 25789 12587 25792
rect 12529 25783 12587 25789
rect 13265 25789 13277 25792
rect 13311 25789 13323 25823
rect 13265 25783 13323 25789
rect 14369 25823 14427 25829
rect 14369 25789 14381 25823
rect 14415 25820 14427 25823
rect 14936 25820 14964 25851
rect 15102 25848 15108 25900
rect 15160 25848 15166 25900
rect 15378 25848 15384 25900
rect 15436 25848 15442 25900
rect 15746 25848 15752 25900
rect 15804 25888 15810 25900
rect 15804 25860 16160 25888
rect 15804 25848 15810 25860
rect 15396 25820 15424 25848
rect 16132 25832 16160 25860
rect 16666 25848 16672 25900
rect 16724 25848 16730 25900
rect 16942 25897 16948 25900
rect 16936 25888 16948 25897
rect 16903 25860 16948 25888
rect 16936 25851 16948 25860
rect 16942 25848 16948 25851
rect 17000 25848 17006 25900
rect 18248 25897 18276 25996
rect 19996 25996 21272 26024
rect 19996 25968 20024 25996
rect 21266 25984 21272 25996
rect 21324 25984 21330 26036
rect 21358 25984 21364 26036
rect 21416 26024 21422 26036
rect 21910 26024 21916 26036
rect 21416 25996 21916 26024
rect 21416 25984 21422 25996
rect 21910 25984 21916 25996
rect 21968 25984 21974 26036
rect 23017 26027 23075 26033
rect 23017 26024 23029 26027
rect 22756 25996 23029 26024
rect 19978 25916 19984 25968
rect 20036 25916 20042 25968
rect 21450 25956 21456 25968
rect 20824 25928 21456 25956
rect 18233 25891 18291 25897
rect 18233 25857 18245 25891
rect 18279 25888 18291 25891
rect 18322 25888 18328 25900
rect 18279 25860 18328 25888
rect 18279 25857 18291 25860
rect 18233 25851 18291 25857
rect 18322 25848 18328 25860
rect 18380 25888 18386 25900
rect 19334 25888 19340 25900
rect 18380 25860 19340 25888
rect 18380 25848 18386 25860
rect 19334 25848 19340 25860
rect 19392 25848 19398 25900
rect 19794 25848 19800 25900
rect 19852 25888 19858 25900
rect 20257 25891 20315 25897
rect 20257 25888 20269 25891
rect 19852 25860 20269 25888
rect 19852 25848 19858 25860
rect 20257 25857 20269 25860
rect 20303 25857 20315 25891
rect 20257 25851 20315 25857
rect 20346 25848 20352 25900
rect 20404 25888 20410 25900
rect 20824 25897 20852 25928
rect 21450 25916 21456 25928
rect 21508 25916 21514 25968
rect 21818 25916 21824 25968
rect 21876 25956 21882 25968
rect 22646 25956 22652 25968
rect 21876 25928 22652 25956
rect 21876 25916 21882 25928
rect 21637 25900 21695 25903
rect 20441 25891 20499 25897
rect 20441 25888 20453 25891
rect 20404 25860 20453 25888
rect 20404 25848 20410 25860
rect 20441 25857 20453 25860
rect 20487 25857 20499 25891
rect 20441 25851 20499 25857
rect 20809 25891 20867 25897
rect 20809 25857 20821 25891
rect 20855 25857 20867 25891
rect 20809 25851 20867 25857
rect 21082 25848 21088 25900
rect 21140 25848 21146 25900
rect 21634 25848 21640 25900
rect 21692 25894 21698 25900
rect 21692 25866 21731 25894
rect 22061 25891 22119 25897
rect 22061 25888 22073 25891
rect 21692 25848 21698 25866
rect 21836 25860 22073 25888
rect 15841 25823 15899 25829
rect 15841 25820 15853 25823
rect 14415 25792 14872 25820
rect 14936 25792 15240 25820
rect 15396 25792 15853 25820
rect 14415 25789 14427 25792
rect 14369 25783 14427 25789
rect 10594 25712 10600 25764
rect 10652 25752 10658 25764
rect 12253 25755 12311 25761
rect 12253 25752 12265 25755
rect 10652 25724 12265 25752
rect 10652 25712 10658 25724
rect 12253 25721 12265 25724
rect 12299 25721 12311 25755
rect 12253 25715 12311 25721
rect 12621 25755 12679 25761
rect 12621 25721 12633 25755
rect 12667 25721 12679 25755
rect 12621 25715 12679 25721
rect 11330 25644 11336 25696
rect 11388 25684 11394 25696
rect 11701 25687 11759 25693
rect 11701 25684 11713 25687
rect 11388 25656 11713 25684
rect 11388 25644 11394 25656
rect 11701 25653 11713 25656
rect 11747 25684 11759 25687
rect 11974 25684 11980 25696
rect 11747 25656 11980 25684
rect 11747 25653 11759 25656
rect 11701 25647 11759 25653
rect 11974 25644 11980 25656
rect 12032 25644 12038 25696
rect 12066 25644 12072 25696
rect 12124 25684 12130 25696
rect 12636 25684 12664 25715
rect 14844 25696 14872 25792
rect 15212 25696 15240 25792
rect 15841 25789 15853 25792
rect 15887 25789 15899 25823
rect 15841 25783 15899 25789
rect 16114 25780 16120 25832
rect 16172 25780 16178 25832
rect 16390 25780 16396 25832
rect 16448 25780 16454 25832
rect 20533 25823 20591 25829
rect 20533 25789 20545 25823
rect 20579 25820 20591 25823
rect 20717 25823 20775 25829
rect 20717 25820 20729 25823
rect 20579 25792 20729 25820
rect 20579 25789 20591 25792
rect 20533 25783 20591 25789
rect 20717 25789 20729 25792
rect 20763 25789 20775 25823
rect 20717 25783 20775 25789
rect 21358 25780 21364 25832
rect 21416 25780 21422 25832
rect 15473 25755 15531 25761
rect 15473 25721 15485 25755
rect 15519 25752 15531 25755
rect 16408 25752 16436 25780
rect 15519 25724 16436 25752
rect 18049 25755 18107 25761
rect 15519 25721 15531 25724
rect 15473 25715 15531 25721
rect 18049 25721 18061 25755
rect 18095 25752 18107 25755
rect 18414 25752 18420 25764
rect 18095 25724 18420 25752
rect 18095 25721 18107 25724
rect 18049 25715 18107 25721
rect 18414 25712 18420 25724
rect 18472 25712 18478 25764
rect 19518 25712 19524 25764
rect 19576 25752 19582 25764
rect 20993 25755 21051 25761
rect 20993 25752 21005 25755
rect 19576 25724 21005 25752
rect 19576 25712 19582 25724
rect 20993 25721 21005 25724
rect 21039 25721 21051 25755
rect 20993 25715 21051 25721
rect 21453 25755 21511 25761
rect 21453 25721 21465 25755
rect 21499 25752 21511 25755
rect 21836 25752 21864 25860
rect 22061 25857 22073 25860
rect 22107 25857 22119 25891
rect 22061 25851 22119 25857
rect 22278 25848 22284 25900
rect 22336 25848 22342 25900
rect 22388 25897 22416 25928
rect 22646 25916 22652 25928
rect 22704 25916 22710 25968
rect 22373 25891 22431 25897
rect 22373 25857 22385 25891
rect 22419 25857 22431 25891
rect 22373 25851 22431 25857
rect 21499 25724 21864 25752
rect 22189 25755 22247 25761
rect 21499 25721 21511 25724
rect 21453 25715 21511 25721
rect 22189 25721 22201 25755
rect 22235 25721 22247 25755
rect 22756 25752 22784 25996
rect 23017 25993 23029 25996
rect 23063 26024 23075 26027
rect 23063 25996 24256 26024
rect 23063 25993 23075 25996
rect 23017 25987 23075 25993
rect 23937 25959 23995 25965
rect 23937 25956 23949 25959
rect 22848 25928 23949 25956
rect 22848 25897 22876 25928
rect 23937 25925 23949 25928
rect 23983 25925 23995 25959
rect 23937 25919 23995 25925
rect 22833 25891 22891 25897
rect 22833 25857 22845 25891
rect 22879 25857 22891 25891
rect 22833 25851 22891 25857
rect 23106 25848 23112 25900
rect 23164 25888 23170 25900
rect 24228 25897 24256 25996
rect 24121 25891 24179 25897
rect 24121 25888 24133 25891
rect 23164 25860 24133 25888
rect 23164 25848 23170 25860
rect 24121 25857 24133 25860
rect 24167 25857 24179 25891
rect 24121 25851 24179 25857
rect 24213 25891 24271 25897
rect 24213 25857 24225 25891
rect 24259 25857 24271 25891
rect 24213 25851 24271 25857
rect 23750 25780 23756 25832
rect 23808 25780 23814 25832
rect 23842 25780 23848 25832
rect 23900 25820 23906 25832
rect 23937 25823 23995 25829
rect 23937 25820 23949 25823
rect 23900 25792 23949 25820
rect 23900 25780 23906 25792
rect 23937 25789 23949 25792
rect 23983 25789 23995 25823
rect 23937 25783 23995 25789
rect 22189 25715 22247 25721
rect 22388 25724 22784 25752
rect 12124 25656 12664 25684
rect 12124 25644 12130 25656
rect 13170 25644 13176 25696
rect 13228 25684 13234 25696
rect 13633 25687 13691 25693
rect 13633 25684 13645 25687
rect 13228 25656 13645 25684
rect 13228 25644 13234 25656
rect 13633 25653 13645 25656
rect 13679 25653 13691 25687
rect 13633 25647 13691 25653
rect 14550 25644 14556 25696
rect 14608 25644 14614 25696
rect 14826 25644 14832 25696
rect 14884 25644 14890 25696
rect 15194 25644 15200 25696
rect 15252 25644 15258 25696
rect 15381 25687 15439 25693
rect 15381 25653 15393 25687
rect 15427 25684 15439 25687
rect 15930 25684 15936 25696
rect 15427 25656 15936 25684
rect 15427 25653 15439 25656
rect 15381 25647 15439 25653
rect 15930 25644 15936 25656
rect 15988 25644 15994 25696
rect 16482 25644 16488 25696
rect 16540 25644 16546 25696
rect 20070 25644 20076 25696
rect 20128 25644 20134 25696
rect 21545 25687 21603 25693
rect 21545 25653 21557 25687
rect 21591 25684 21603 25687
rect 22094 25684 22100 25696
rect 21591 25656 22100 25684
rect 21591 25653 21603 25656
rect 21545 25647 21603 25653
rect 22094 25644 22100 25656
rect 22152 25644 22158 25696
rect 22204 25684 22232 25715
rect 22388 25696 22416 25724
rect 22370 25684 22376 25696
rect 22204 25656 22376 25684
rect 22370 25644 22376 25656
rect 22428 25644 22434 25696
rect 22554 25644 22560 25696
rect 22612 25644 22618 25696
rect 22646 25644 22652 25696
rect 22704 25644 22710 25696
rect 23106 25644 23112 25696
rect 23164 25684 23170 25696
rect 23201 25687 23259 25693
rect 23201 25684 23213 25687
rect 23164 25656 23213 25684
rect 23164 25644 23170 25656
rect 23201 25653 23213 25656
rect 23247 25653 23259 25687
rect 23201 25647 23259 25653
rect 1104 25594 34868 25616
rect 1104 25542 5170 25594
rect 5222 25542 5234 25594
rect 5286 25542 5298 25594
rect 5350 25542 5362 25594
rect 5414 25542 5426 25594
rect 5478 25542 13611 25594
rect 13663 25542 13675 25594
rect 13727 25542 13739 25594
rect 13791 25542 13803 25594
rect 13855 25542 13867 25594
rect 13919 25542 22052 25594
rect 22104 25542 22116 25594
rect 22168 25542 22180 25594
rect 22232 25542 22244 25594
rect 22296 25542 22308 25594
rect 22360 25542 30493 25594
rect 30545 25542 30557 25594
rect 30609 25542 30621 25594
rect 30673 25542 30685 25594
rect 30737 25542 30749 25594
rect 30801 25542 34868 25594
rect 1104 25520 34868 25542
rect 11057 25483 11115 25489
rect 11057 25449 11069 25483
rect 11103 25480 11115 25483
rect 12066 25480 12072 25492
rect 11103 25452 12072 25480
rect 11103 25449 11115 25452
rect 11057 25443 11115 25449
rect 12066 25440 12072 25452
rect 12124 25440 12130 25492
rect 12710 25440 12716 25492
rect 12768 25480 12774 25492
rect 12897 25483 12955 25489
rect 12897 25480 12909 25483
rect 12768 25452 12909 25480
rect 12768 25440 12774 25452
rect 12897 25449 12909 25452
rect 12943 25449 12955 25483
rect 12897 25443 12955 25449
rect 13354 25440 13360 25492
rect 13412 25440 13418 25492
rect 13446 25440 13452 25492
rect 13504 25440 13510 25492
rect 13722 25440 13728 25492
rect 13780 25480 13786 25492
rect 14826 25480 14832 25492
rect 13780 25452 14832 25480
rect 13780 25440 13786 25452
rect 14826 25440 14832 25452
rect 14884 25440 14890 25492
rect 15194 25440 15200 25492
rect 15252 25480 15258 25492
rect 15565 25483 15623 25489
rect 15565 25480 15577 25483
rect 15252 25452 15577 25480
rect 15252 25440 15258 25452
rect 15565 25449 15577 25452
rect 15611 25449 15623 25483
rect 16574 25480 16580 25492
rect 15565 25443 15623 25449
rect 16224 25452 16580 25480
rect 10226 25372 10232 25424
rect 10284 25412 10290 25424
rect 10505 25415 10563 25421
rect 10505 25412 10517 25415
rect 10284 25384 10517 25412
rect 10284 25372 10290 25384
rect 10505 25381 10517 25384
rect 10551 25412 10563 25415
rect 12621 25415 12679 25421
rect 10551 25384 11652 25412
rect 10551 25381 10563 25384
rect 10505 25375 10563 25381
rect 10134 25304 10140 25356
rect 10192 25344 10198 25356
rect 10689 25347 10747 25353
rect 10689 25344 10701 25347
rect 10192 25316 10701 25344
rect 10192 25304 10198 25316
rect 10689 25313 10701 25316
rect 10735 25344 10747 25347
rect 11238 25344 11244 25356
rect 10735 25316 11244 25344
rect 10735 25313 10747 25316
rect 10689 25307 10747 25313
rect 11238 25304 11244 25316
rect 11296 25304 11302 25356
rect 11624 25353 11652 25384
rect 12621 25381 12633 25415
rect 12667 25412 12679 25415
rect 13464 25412 13492 25440
rect 12667 25384 13492 25412
rect 12667 25381 12679 25384
rect 12621 25375 12679 25381
rect 14550 25372 14556 25424
rect 14608 25372 14614 25424
rect 15286 25372 15292 25424
rect 15344 25412 15350 25424
rect 15344 25384 15700 25412
rect 15344 25372 15350 25384
rect 11609 25347 11667 25353
rect 11609 25313 11621 25347
rect 11655 25344 11667 25347
rect 11882 25344 11888 25356
rect 11655 25316 11888 25344
rect 11655 25313 11667 25316
rect 11609 25307 11667 25313
rect 11882 25304 11888 25316
rect 11940 25304 11946 25356
rect 11974 25304 11980 25356
rect 12032 25344 12038 25356
rect 12805 25347 12863 25353
rect 12032 25316 12756 25344
rect 12032 25304 12038 25316
rect 10321 25279 10379 25285
rect 10321 25245 10333 25279
rect 10367 25245 10379 25279
rect 10321 25239 10379 25245
rect 10505 25279 10563 25285
rect 10505 25245 10517 25279
rect 10551 25276 10563 25279
rect 10594 25276 10600 25288
rect 10551 25248 10600 25276
rect 10551 25245 10563 25248
rect 10505 25239 10563 25245
rect 10336 25208 10364 25239
rect 10594 25236 10600 25248
rect 10652 25236 10658 25288
rect 10781 25279 10839 25285
rect 10781 25245 10793 25279
rect 10827 25276 10839 25279
rect 11330 25276 11336 25288
rect 10827 25248 11336 25276
rect 10827 25245 10839 25248
rect 10781 25239 10839 25245
rect 11330 25236 11336 25248
rect 11388 25236 11394 25288
rect 11422 25236 11428 25288
rect 11480 25236 11486 25288
rect 11701 25279 11759 25285
rect 11701 25245 11713 25279
rect 11747 25276 11759 25279
rect 12158 25276 12164 25288
rect 11747 25248 12164 25276
rect 11747 25245 11759 25248
rect 11701 25239 11759 25245
rect 12158 25236 12164 25248
rect 12216 25236 12222 25288
rect 12250 25236 12256 25288
rect 12308 25236 12314 25288
rect 12437 25279 12495 25285
rect 12437 25245 12449 25279
rect 12483 25276 12495 25279
rect 12618 25276 12624 25288
rect 12483 25248 12624 25276
rect 12483 25245 12495 25248
rect 12437 25239 12495 25245
rect 12618 25236 12624 25248
rect 12676 25236 12682 25288
rect 12728 25285 12756 25316
rect 12805 25313 12817 25347
rect 12851 25344 12863 25347
rect 12894 25344 12900 25356
rect 12851 25316 12900 25344
rect 12851 25313 12863 25316
rect 12805 25307 12863 25313
rect 12894 25304 12900 25316
rect 12952 25304 12958 25356
rect 12989 25347 13047 25353
rect 12989 25313 13001 25347
rect 13035 25344 13047 25347
rect 13909 25347 13967 25353
rect 13035 25316 13216 25344
rect 13035 25313 13047 25316
rect 12989 25307 13047 25313
rect 12713 25279 12771 25285
rect 12713 25245 12725 25279
rect 12759 25245 12771 25279
rect 12713 25239 12771 25245
rect 10962 25208 10968 25220
rect 10336 25180 10968 25208
rect 10962 25168 10968 25180
rect 11020 25208 11026 25220
rect 11793 25211 11851 25217
rect 11793 25208 11805 25211
rect 11020 25180 11805 25208
rect 11020 25168 11026 25180
rect 11793 25177 11805 25180
rect 11839 25177 11851 25211
rect 11793 25171 11851 25177
rect 11974 25168 11980 25220
rect 12032 25168 12038 25220
rect 12912 25208 12940 25304
rect 13188 25288 13216 25316
rect 13909 25313 13921 25347
rect 13955 25313 13967 25347
rect 14568 25344 14596 25372
rect 14568 25316 15516 25344
rect 13909 25307 13967 25313
rect 13170 25236 13176 25288
rect 13228 25276 13234 25288
rect 13357 25279 13415 25285
rect 13357 25276 13369 25279
rect 13228 25248 13369 25276
rect 13228 25236 13234 25248
rect 13357 25245 13369 25248
rect 13403 25245 13415 25279
rect 13357 25239 13415 25245
rect 13541 25279 13599 25285
rect 13541 25245 13553 25279
rect 13587 25245 13599 25279
rect 13541 25239 13599 25245
rect 13633 25279 13691 25285
rect 13633 25245 13645 25279
rect 13679 25245 13691 25279
rect 13924 25276 13952 25307
rect 14645 25279 14703 25285
rect 13924 25248 14596 25276
rect 13633 25239 13691 25245
rect 13556 25208 13584 25239
rect 12912 25180 13584 25208
rect 11241 25143 11299 25149
rect 11241 25109 11253 25143
rect 11287 25140 11299 25143
rect 11514 25140 11520 25152
rect 11287 25112 11520 25140
rect 11287 25109 11299 25112
rect 11241 25103 11299 25109
rect 11514 25100 11520 25112
rect 11572 25100 11578 25152
rect 13354 25100 13360 25152
rect 13412 25140 13418 25152
rect 13648 25140 13676 25239
rect 14182 25168 14188 25220
rect 14240 25208 14246 25220
rect 14277 25211 14335 25217
rect 14277 25208 14289 25211
rect 14240 25180 14289 25208
rect 14240 25168 14246 25180
rect 14277 25177 14289 25180
rect 14323 25177 14335 25211
rect 14277 25171 14335 25177
rect 14458 25168 14464 25220
rect 14516 25168 14522 25220
rect 14568 25208 14596 25248
rect 14645 25245 14657 25279
rect 14691 25276 14703 25279
rect 14737 25279 14795 25285
rect 14737 25276 14749 25279
rect 14691 25248 14749 25276
rect 14691 25245 14703 25248
rect 14645 25239 14703 25245
rect 14737 25245 14749 25248
rect 14783 25245 14795 25279
rect 14737 25239 14795 25245
rect 14918 25236 14924 25288
rect 14976 25236 14982 25288
rect 15102 25236 15108 25288
rect 15160 25236 15166 25288
rect 15488 25285 15516 25316
rect 15672 25288 15700 25384
rect 16224 25353 16252 25452
rect 16574 25440 16580 25452
rect 16632 25440 16638 25492
rect 17402 25440 17408 25492
rect 17460 25480 17466 25492
rect 18785 25483 18843 25489
rect 18785 25480 18797 25483
rect 17460 25452 18797 25480
rect 17460 25440 17466 25452
rect 18785 25449 18797 25452
rect 18831 25449 18843 25483
rect 18785 25443 18843 25449
rect 19702 25440 19708 25492
rect 19760 25440 19766 25492
rect 20070 25440 20076 25492
rect 20128 25440 20134 25492
rect 20809 25483 20867 25489
rect 20809 25449 20821 25483
rect 20855 25480 20867 25483
rect 20898 25480 20904 25492
rect 20855 25452 20904 25480
rect 20855 25449 20867 25452
rect 20809 25443 20867 25449
rect 20898 25440 20904 25452
rect 20956 25440 20962 25492
rect 22281 25483 22339 25489
rect 22281 25449 22293 25483
rect 22327 25480 22339 25483
rect 22370 25480 22376 25492
rect 22327 25452 22376 25480
rect 22327 25449 22339 25452
rect 22281 25443 22339 25449
rect 22370 25440 22376 25452
rect 22428 25440 22434 25492
rect 17589 25415 17647 25421
rect 17589 25381 17601 25415
rect 17635 25412 17647 25415
rect 19720 25412 19748 25440
rect 17635 25384 19748 25412
rect 17635 25381 17647 25384
rect 17589 25375 17647 25381
rect 17696 25353 17724 25384
rect 16209 25347 16267 25353
rect 16209 25313 16221 25347
rect 16255 25313 16267 25347
rect 16209 25307 16267 25313
rect 17681 25347 17739 25353
rect 17681 25313 17693 25347
rect 17727 25313 17739 25347
rect 17681 25307 17739 25313
rect 18782 25304 18788 25356
rect 18840 25304 18846 25356
rect 19518 25304 19524 25356
rect 19576 25344 19582 25356
rect 19576 25316 19748 25344
rect 19576 25304 19582 25316
rect 15473 25279 15531 25285
rect 15473 25245 15485 25279
rect 15519 25245 15531 25279
rect 15473 25239 15531 25245
rect 15654 25236 15660 25288
rect 15712 25236 15718 25288
rect 16482 25285 16488 25288
rect 16476 25276 16488 25285
rect 16443 25248 16488 25276
rect 16476 25239 16488 25248
rect 16482 25236 16488 25239
rect 16540 25236 16546 25288
rect 17957 25279 18015 25285
rect 17957 25245 17969 25279
rect 18003 25276 18015 25279
rect 18800 25276 18828 25304
rect 19426 25285 19432 25288
rect 18003 25248 18736 25276
rect 18800 25248 19012 25276
rect 18003 25245 18015 25248
rect 17957 25239 18015 25245
rect 14936 25208 14964 25236
rect 14568 25180 14964 25208
rect 13412 25112 13676 25140
rect 13909 25143 13967 25149
rect 13412 25100 13418 25112
rect 13909 25109 13921 25143
rect 13955 25140 13967 25143
rect 14366 25140 14372 25152
rect 13955 25112 14372 25140
rect 13955 25109 13967 25112
rect 13909 25103 13967 25109
rect 14366 25100 14372 25112
rect 14424 25100 14430 25152
rect 14467 25140 14495 25168
rect 15120 25140 15148 25236
rect 16114 25168 16120 25220
rect 16172 25208 16178 25220
rect 17972 25208 18000 25239
rect 16172 25180 18000 25208
rect 18708 25208 18736 25248
rect 18984 25217 19012 25248
rect 19424 25239 19432 25285
rect 19426 25236 19432 25239
rect 19484 25236 19490 25288
rect 19610 25236 19616 25288
rect 19668 25236 19674 25288
rect 19720 25285 19748 25316
rect 19720 25279 19799 25285
rect 19720 25248 19753 25279
rect 19741 25245 19753 25248
rect 19787 25245 19799 25279
rect 19741 25239 19799 25245
rect 19889 25279 19947 25285
rect 19889 25245 19901 25279
rect 19935 25276 19947 25279
rect 20088 25276 20116 25440
rect 20349 25415 20407 25421
rect 20349 25381 20361 25415
rect 20395 25412 20407 25415
rect 21266 25412 21272 25424
rect 20395 25384 21272 25412
rect 20395 25381 20407 25384
rect 20349 25375 20407 25381
rect 21266 25372 21272 25384
rect 21324 25372 21330 25424
rect 21726 25344 21732 25356
rect 20732 25316 21732 25344
rect 19935 25248 20116 25276
rect 19935 25245 19947 25248
rect 19889 25239 19947 25245
rect 20162 25236 20168 25288
rect 20220 25236 20226 25288
rect 20732 25285 20760 25316
rect 21726 25304 21732 25316
rect 21784 25304 21790 25356
rect 21910 25304 21916 25356
rect 21968 25304 21974 25356
rect 22830 25304 22836 25356
rect 22888 25304 22894 25356
rect 20625 25279 20683 25285
rect 20625 25245 20637 25279
rect 20671 25245 20683 25279
rect 20625 25239 20683 25245
rect 20717 25279 20775 25285
rect 20717 25245 20729 25279
rect 20763 25245 20775 25279
rect 20717 25239 20775 25245
rect 20901 25279 20959 25285
rect 20901 25245 20913 25279
rect 20947 25276 20959 25279
rect 21174 25276 21180 25288
rect 20947 25248 21180 25276
rect 20947 25245 20959 25248
rect 20901 25239 20959 25245
rect 18969 25211 19027 25217
rect 18708 25180 18828 25208
rect 16172 25168 16178 25180
rect 14467 25112 15148 25140
rect 18598 25100 18604 25152
rect 18656 25100 18662 25152
rect 18800 25149 18828 25180
rect 18969 25177 18981 25211
rect 19015 25177 19027 25211
rect 18969 25171 19027 25177
rect 19518 25168 19524 25220
rect 19576 25168 19582 25220
rect 20180 25208 20208 25236
rect 20349 25211 20407 25217
rect 20349 25208 20361 25211
rect 20180 25180 20361 25208
rect 20349 25177 20361 25180
rect 20395 25208 20407 25211
rect 20438 25208 20444 25220
rect 20395 25180 20444 25208
rect 20395 25177 20407 25180
rect 20349 25171 20407 25177
rect 20438 25168 20444 25180
rect 20496 25168 20502 25220
rect 20640 25208 20668 25239
rect 21174 25236 21180 25248
rect 21232 25236 21238 25288
rect 21634 25236 21640 25288
rect 21692 25276 21698 25288
rect 23106 25285 23112 25288
rect 22005 25279 22063 25285
rect 22005 25276 22017 25279
rect 21692 25248 22017 25276
rect 21692 25236 21698 25248
rect 22005 25245 22017 25248
rect 22051 25276 22063 25279
rect 23100 25276 23112 25285
rect 22051 25248 22876 25276
rect 23067 25248 23112 25276
rect 22051 25245 22063 25248
rect 22005 25239 22063 25245
rect 20640 25180 20852 25208
rect 20824 25152 20852 25180
rect 21818 25168 21824 25220
rect 21876 25208 21882 25220
rect 22554 25208 22560 25220
rect 21876 25180 22560 25208
rect 21876 25168 21882 25180
rect 22554 25168 22560 25180
rect 22612 25168 22618 25220
rect 22848 25208 22876 25248
rect 23100 25239 23112 25248
rect 23106 25236 23112 25239
rect 23164 25236 23170 25288
rect 24210 25236 24216 25288
rect 24268 25276 24274 25288
rect 25041 25279 25099 25285
rect 25041 25276 25053 25279
rect 24268 25248 25053 25276
rect 24268 25236 24274 25248
rect 25041 25245 25053 25248
rect 25087 25245 25099 25279
rect 25041 25239 25099 25245
rect 23014 25208 23020 25220
rect 22848 25180 23020 25208
rect 23014 25168 23020 25180
rect 23072 25168 23078 25220
rect 18759 25143 18828 25149
rect 18759 25109 18771 25143
rect 18805 25112 18828 25143
rect 19245 25143 19303 25149
rect 18805 25109 18817 25112
rect 18759 25103 18817 25109
rect 19245 25109 19257 25143
rect 19291 25140 19303 25143
rect 20162 25140 20168 25152
rect 19291 25112 20168 25140
rect 19291 25109 19303 25112
rect 19245 25103 19303 25109
rect 20162 25100 20168 25112
rect 20220 25100 20226 25152
rect 20533 25143 20591 25149
rect 20533 25109 20545 25143
rect 20579 25140 20591 25143
rect 20714 25140 20720 25152
rect 20579 25112 20720 25140
rect 20579 25109 20591 25112
rect 20533 25103 20591 25109
rect 20714 25100 20720 25112
rect 20772 25100 20778 25152
rect 20806 25100 20812 25152
rect 20864 25140 20870 25152
rect 23842 25140 23848 25152
rect 20864 25112 23848 25140
rect 20864 25100 20870 25112
rect 23842 25100 23848 25112
rect 23900 25100 23906 25152
rect 24210 25100 24216 25152
rect 24268 25100 24274 25152
rect 24854 25100 24860 25152
rect 24912 25100 24918 25152
rect 1104 25050 35027 25072
rect 1104 24998 9390 25050
rect 9442 24998 9454 25050
rect 9506 24998 9518 25050
rect 9570 24998 9582 25050
rect 9634 24998 9646 25050
rect 9698 24998 17831 25050
rect 17883 24998 17895 25050
rect 17947 24998 17959 25050
rect 18011 24998 18023 25050
rect 18075 24998 18087 25050
rect 18139 24998 26272 25050
rect 26324 24998 26336 25050
rect 26388 24998 26400 25050
rect 26452 24998 26464 25050
rect 26516 24998 26528 25050
rect 26580 24998 34713 25050
rect 34765 24998 34777 25050
rect 34829 24998 34841 25050
rect 34893 24998 34905 25050
rect 34957 24998 34969 25050
rect 35021 24998 35027 25050
rect 1104 24976 35027 24998
rect 10594 24896 10600 24948
rect 10652 24896 10658 24948
rect 11054 24896 11060 24948
rect 11112 24936 11118 24948
rect 11974 24936 11980 24948
rect 11112 24908 11980 24936
rect 11112 24896 11118 24908
rect 11974 24896 11980 24908
rect 12032 24896 12038 24948
rect 12158 24896 12164 24948
rect 12216 24896 12222 24948
rect 12250 24896 12256 24948
rect 12308 24936 12314 24948
rect 13449 24939 13507 24945
rect 13449 24936 13461 24939
rect 12308 24908 13461 24936
rect 12308 24896 12314 24908
rect 13449 24905 13461 24908
rect 13495 24905 13507 24939
rect 13449 24899 13507 24905
rect 14277 24939 14335 24945
rect 14277 24905 14289 24939
rect 14323 24936 14335 24939
rect 14918 24936 14924 24948
rect 14323 24908 14924 24936
rect 14323 24905 14335 24908
rect 14277 24899 14335 24905
rect 14918 24896 14924 24908
rect 14976 24896 14982 24948
rect 17402 24896 17408 24948
rect 17460 24896 17466 24948
rect 19245 24939 19303 24945
rect 19245 24905 19257 24939
rect 19291 24936 19303 24939
rect 19518 24936 19524 24948
rect 19291 24908 19524 24936
rect 19291 24905 19303 24908
rect 19245 24899 19303 24905
rect 19518 24896 19524 24908
rect 19576 24936 19582 24948
rect 19576 24908 19656 24936
rect 19576 24896 19582 24908
rect 10612 24868 10640 24896
rect 12176 24868 12204 24896
rect 14458 24868 14464 24880
rect 9876 24840 10456 24868
rect 10612 24840 10916 24868
rect 9769 24803 9827 24809
rect 9769 24769 9781 24803
rect 9815 24800 9827 24803
rect 9876 24800 9904 24840
rect 9815 24772 9904 24800
rect 9953 24803 10011 24809
rect 9815 24769 9827 24772
rect 9769 24763 9827 24769
rect 9953 24769 9965 24803
rect 9999 24800 10011 24803
rect 10134 24800 10140 24812
rect 9999 24772 10140 24800
rect 9999 24769 10011 24772
rect 9953 24763 10011 24769
rect 10134 24760 10140 24772
rect 10192 24760 10198 24812
rect 10226 24760 10232 24812
rect 10284 24760 10290 24812
rect 10321 24803 10379 24809
rect 10321 24769 10333 24803
rect 10367 24769 10379 24803
rect 10428 24800 10456 24840
rect 10502 24800 10508 24812
rect 10428 24772 10508 24800
rect 10321 24763 10379 24769
rect 10336 24732 10364 24763
rect 10502 24760 10508 24772
rect 10560 24760 10566 24812
rect 10594 24760 10600 24812
rect 10652 24760 10658 24812
rect 10888 24809 10916 24840
rect 12084 24840 12204 24868
rect 14292 24840 14464 24868
rect 10873 24803 10931 24809
rect 10873 24769 10885 24803
rect 10919 24769 10931 24803
rect 10873 24763 10931 24769
rect 10962 24760 10968 24812
rect 11020 24760 11026 24812
rect 11054 24760 11060 24812
rect 11112 24760 11118 24812
rect 11146 24760 11152 24812
rect 11204 24800 11210 24812
rect 12084 24809 12112 24840
rect 11333 24803 11391 24809
rect 11333 24800 11345 24803
rect 11204 24772 11345 24800
rect 11204 24760 11210 24772
rect 11333 24769 11345 24772
rect 11379 24800 11391 24803
rect 11609 24803 11667 24809
rect 11609 24800 11621 24803
rect 11379 24772 11621 24800
rect 11379 24769 11391 24772
rect 11333 24763 11391 24769
rect 11609 24769 11621 24772
rect 11655 24769 11667 24803
rect 11609 24763 11667 24769
rect 12069 24803 12127 24809
rect 12069 24769 12081 24803
rect 12115 24769 12127 24803
rect 12069 24763 12127 24769
rect 12345 24803 12403 24809
rect 12345 24769 12357 24803
rect 12391 24769 12403 24803
rect 12345 24763 12403 24769
rect 10689 24735 10747 24741
rect 10689 24732 10701 24735
rect 10336 24704 10701 24732
rect 10689 24701 10701 24704
rect 10735 24701 10747 24735
rect 10689 24695 10747 24701
rect 9953 24667 10011 24673
rect 9953 24633 9965 24667
rect 9999 24664 10011 24667
rect 11072 24664 11100 24760
rect 9999 24636 11100 24664
rect 9999 24633 10011 24636
rect 9953 24627 10011 24633
rect 10042 24556 10048 24608
rect 10100 24556 10106 24608
rect 10505 24599 10563 24605
rect 10505 24565 10517 24599
rect 10551 24596 10563 24599
rect 11164 24596 11192 24760
rect 11238 24692 11244 24744
rect 11296 24732 11302 24744
rect 12360 24732 12388 24763
rect 12986 24760 12992 24812
rect 13044 24760 13050 24812
rect 13354 24760 13360 24812
rect 13412 24800 13418 24812
rect 13633 24803 13691 24809
rect 13633 24800 13645 24803
rect 13412 24772 13645 24800
rect 13412 24760 13418 24772
rect 13633 24769 13645 24772
rect 13679 24769 13691 24803
rect 13633 24763 13691 24769
rect 13722 24760 13728 24812
rect 13780 24760 13786 24812
rect 13909 24803 13967 24809
rect 13909 24769 13921 24803
rect 13955 24800 13967 24803
rect 13998 24800 14004 24812
rect 13955 24772 14004 24800
rect 13955 24769 13967 24772
rect 13909 24763 13967 24769
rect 13998 24760 14004 24772
rect 14056 24760 14062 24812
rect 14093 24803 14151 24809
rect 14093 24769 14105 24803
rect 14139 24769 14151 24803
rect 14093 24763 14151 24769
rect 11296 24704 12388 24732
rect 11296 24692 11302 24704
rect 12360 24664 12388 24704
rect 12526 24692 12532 24744
rect 12584 24692 12590 24744
rect 13081 24735 13139 24741
rect 13081 24701 13093 24735
rect 13127 24732 13139 24735
rect 13170 24732 13176 24744
rect 13127 24704 13176 24732
rect 13127 24701 13139 24704
rect 13081 24695 13139 24701
rect 13096 24664 13124 24695
rect 13170 24692 13176 24704
rect 13228 24732 13234 24744
rect 14108 24732 14136 24763
rect 14182 24760 14188 24812
rect 14240 24800 14246 24812
rect 14292 24809 14320 24840
rect 14458 24828 14464 24840
rect 14516 24828 14522 24880
rect 15102 24868 15108 24880
rect 14659 24840 15108 24868
rect 14277 24803 14335 24809
rect 14277 24800 14289 24803
rect 14240 24772 14289 24800
rect 14240 24760 14246 24772
rect 14277 24769 14289 24772
rect 14323 24769 14335 24803
rect 14277 24763 14335 24769
rect 14550 24760 14556 24812
rect 14608 24760 14614 24812
rect 14659 24732 14687 24840
rect 15102 24828 15108 24840
rect 15160 24828 15166 24880
rect 15488 24840 15700 24868
rect 14737 24803 14795 24809
rect 14737 24769 14749 24803
rect 14783 24769 14795 24803
rect 14737 24763 14795 24769
rect 13228 24704 14136 24732
rect 14292 24704 14687 24732
rect 14752 24732 14780 24763
rect 14826 24760 14832 24812
rect 14884 24760 14890 24812
rect 15289 24803 15347 24809
rect 15289 24769 15301 24803
rect 15335 24800 15347 24803
rect 15488 24800 15516 24840
rect 15335 24772 15516 24800
rect 15565 24803 15623 24809
rect 15335 24769 15347 24772
rect 15289 24763 15347 24769
rect 15565 24769 15577 24803
rect 15611 24769 15623 24803
rect 15672 24800 15700 24840
rect 17512 24840 17816 24868
rect 16114 24800 16120 24812
rect 15672 24772 16120 24800
rect 15565 24763 15623 24769
rect 15378 24732 15384 24744
rect 14752 24704 15384 24732
rect 13228 24692 13234 24704
rect 14292 24676 14320 24704
rect 15378 24692 15384 24704
rect 15436 24732 15442 24744
rect 15473 24735 15531 24741
rect 15473 24732 15485 24735
rect 15436 24704 15485 24732
rect 15436 24692 15442 24704
rect 15473 24701 15485 24704
rect 15519 24701 15531 24735
rect 15473 24695 15531 24701
rect 11348 24636 11836 24664
rect 12360 24636 13124 24664
rect 13357 24667 13415 24673
rect 11348 24608 11376 24636
rect 10551 24568 11192 24596
rect 10551 24565 10563 24568
rect 10505 24559 10563 24565
rect 11330 24556 11336 24608
rect 11388 24556 11394 24608
rect 11698 24556 11704 24608
rect 11756 24556 11762 24608
rect 11808 24605 11836 24636
rect 13357 24633 13369 24667
rect 13403 24664 13415 24667
rect 13817 24667 13875 24673
rect 13817 24664 13829 24667
rect 13403 24636 13829 24664
rect 13403 24633 13415 24636
rect 13357 24627 13415 24633
rect 13817 24633 13829 24636
rect 13863 24664 13875 24667
rect 14090 24664 14096 24676
rect 13863 24636 14096 24664
rect 13863 24633 13875 24636
rect 13817 24627 13875 24633
rect 14090 24624 14096 24636
rect 14148 24624 14154 24676
rect 14274 24624 14280 24676
rect 14332 24624 14338 24676
rect 14553 24667 14611 24673
rect 14553 24633 14565 24667
rect 14599 24664 14611 24667
rect 15580 24664 15608 24763
rect 16114 24760 16120 24772
rect 16172 24800 16178 24812
rect 16669 24803 16727 24809
rect 16669 24800 16681 24803
rect 16172 24772 16681 24800
rect 16172 24760 16178 24772
rect 16669 24769 16681 24772
rect 16715 24769 16727 24803
rect 16669 24763 16727 24769
rect 17310 24760 17316 24812
rect 17368 24800 17374 24812
rect 17512 24800 17540 24840
rect 17368 24772 17540 24800
rect 17368 24760 17374 24772
rect 17586 24760 17592 24812
rect 17644 24760 17650 24812
rect 17681 24803 17739 24809
rect 17681 24769 17693 24803
rect 17727 24769 17739 24803
rect 17788 24800 17816 24840
rect 19426 24828 19432 24880
rect 19484 24828 19490 24880
rect 17865 24803 17923 24809
rect 17865 24800 17877 24803
rect 17788 24772 17877 24800
rect 17681 24763 17739 24769
rect 17865 24769 17877 24772
rect 17911 24769 17923 24803
rect 17865 24763 17923 24769
rect 17957 24803 18015 24809
rect 17957 24769 17969 24803
rect 18003 24769 18015 24803
rect 17957 24763 18015 24769
rect 15654 24692 15660 24744
rect 15712 24732 15718 24744
rect 15838 24732 15844 24744
rect 15712 24704 15844 24732
rect 15712 24692 15718 24704
rect 15838 24692 15844 24704
rect 15896 24692 15902 24744
rect 15930 24692 15936 24744
rect 15988 24732 15994 24744
rect 17221 24735 17279 24741
rect 17221 24732 17233 24735
rect 15988 24704 17233 24732
rect 15988 24692 15994 24704
rect 17221 24701 17233 24704
rect 17267 24701 17279 24735
rect 17696 24732 17724 24763
rect 17972 24732 18000 24763
rect 18138 24760 18144 24812
rect 18196 24760 18202 24812
rect 18230 24760 18236 24812
rect 18288 24760 18294 24812
rect 19628 24809 19656 24908
rect 20714 24896 20720 24948
rect 20772 24936 20778 24948
rect 21542 24936 21548 24948
rect 20772 24908 21548 24936
rect 20772 24896 20778 24908
rect 21542 24896 21548 24908
rect 21600 24936 21606 24948
rect 21821 24939 21879 24945
rect 21821 24936 21833 24939
rect 21600 24908 21833 24936
rect 21600 24896 21606 24908
rect 21821 24905 21833 24908
rect 21867 24905 21879 24939
rect 21821 24899 21879 24905
rect 22646 24896 22652 24948
rect 22704 24896 22710 24948
rect 22664 24868 22692 24896
rect 22664 24840 22876 24868
rect 19337 24803 19395 24809
rect 19337 24769 19349 24803
rect 19383 24769 19395 24803
rect 19337 24763 19395 24769
rect 19613 24803 19671 24809
rect 19613 24769 19625 24803
rect 19659 24769 19671 24803
rect 19613 24763 19671 24769
rect 18248 24732 18276 24760
rect 17696 24704 17908 24732
rect 17972 24704 18276 24732
rect 17221 24695 17279 24701
rect 14599 24636 15608 24664
rect 14599 24633 14611 24636
rect 14553 24627 14611 24633
rect 17034 24624 17040 24676
rect 17092 24664 17098 24676
rect 17681 24667 17739 24673
rect 17681 24664 17693 24667
rect 17092 24636 17693 24664
rect 17092 24624 17098 24636
rect 17681 24633 17693 24636
rect 17727 24633 17739 24667
rect 17880 24664 17908 24704
rect 19352 24664 19380 24763
rect 19978 24760 19984 24812
rect 20036 24760 20042 24812
rect 20254 24809 20260 24812
rect 20248 24763 20260 24809
rect 20254 24760 20260 24763
rect 20312 24760 20318 24812
rect 22462 24760 22468 24812
rect 22520 24800 22526 24812
rect 22848 24809 22876 24840
rect 22649 24803 22707 24809
rect 22649 24800 22661 24803
rect 22520 24772 22661 24800
rect 22520 24760 22526 24772
rect 22649 24769 22661 24772
rect 22695 24769 22707 24803
rect 22649 24763 22707 24769
rect 22833 24803 22891 24809
rect 22833 24769 22845 24803
rect 22879 24769 22891 24803
rect 22833 24763 22891 24769
rect 22925 24803 22983 24809
rect 22925 24769 22937 24803
rect 22971 24769 22983 24803
rect 22925 24763 22983 24769
rect 21450 24692 21456 24744
rect 21508 24732 21514 24744
rect 22373 24735 22431 24741
rect 22373 24732 22385 24735
rect 21508 24704 22385 24732
rect 21508 24692 21514 24704
rect 22373 24701 22385 24704
rect 22419 24701 22431 24735
rect 22940 24732 22968 24763
rect 23014 24760 23020 24812
rect 23072 24800 23078 24812
rect 24854 24800 24860 24812
rect 23072 24772 24860 24800
rect 23072 24760 23078 24772
rect 24854 24760 24860 24772
rect 24912 24760 24918 24812
rect 22373 24695 22431 24701
rect 22664 24704 22968 24732
rect 23293 24735 23351 24741
rect 21361 24667 21419 24673
rect 17880 24636 19288 24664
rect 19352 24636 20024 24664
rect 17681 24627 17739 24633
rect 11793 24599 11851 24605
rect 11793 24565 11805 24599
rect 11839 24565 11851 24599
rect 11793 24559 11851 24565
rect 11882 24556 11888 24608
rect 11940 24605 11946 24608
rect 11940 24599 11989 24605
rect 11940 24565 11943 24599
rect 11977 24565 11989 24599
rect 11940 24559 11989 24565
rect 11940 24556 11946 24559
rect 15654 24556 15660 24608
rect 15712 24556 15718 24608
rect 15746 24556 15752 24608
rect 15804 24556 15810 24608
rect 18141 24599 18199 24605
rect 18141 24565 18153 24599
rect 18187 24596 18199 24599
rect 18322 24596 18328 24608
rect 18187 24568 18328 24596
rect 18187 24565 18199 24568
rect 18141 24559 18199 24565
rect 18322 24556 18328 24568
rect 18380 24556 18386 24608
rect 19260 24596 19288 24636
rect 19518 24596 19524 24608
rect 19260 24568 19524 24596
rect 19518 24556 19524 24568
rect 19576 24556 19582 24608
rect 19794 24556 19800 24608
rect 19852 24556 19858 24608
rect 19996 24596 20024 24636
rect 21361 24633 21373 24667
rect 21407 24664 21419 24667
rect 21468 24664 21496 24692
rect 22664 24676 22692 24704
rect 23293 24701 23305 24735
rect 23339 24732 23351 24735
rect 23750 24732 23756 24744
rect 23339 24704 23756 24732
rect 23339 24701 23351 24704
rect 23293 24695 23351 24701
rect 23750 24692 23756 24704
rect 23808 24692 23814 24744
rect 21407 24636 21496 24664
rect 21407 24633 21419 24636
rect 21361 24627 21419 24633
rect 22646 24624 22652 24676
rect 22704 24624 22710 24676
rect 24210 24596 24216 24608
rect 19996 24568 24216 24596
rect 24210 24556 24216 24568
rect 24268 24556 24274 24608
rect 1104 24506 34868 24528
rect 1104 24454 5170 24506
rect 5222 24454 5234 24506
rect 5286 24454 5298 24506
rect 5350 24454 5362 24506
rect 5414 24454 5426 24506
rect 5478 24454 13611 24506
rect 13663 24454 13675 24506
rect 13727 24454 13739 24506
rect 13791 24454 13803 24506
rect 13855 24454 13867 24506
rect 13919 24454 22052 24506
rect 22104 24454 22116 24506
rect 22168 24454 22180 24506
rect 22232 24454 22244 24506
rect 22296 24454 22308 24506
rect 22360 24454 30493 24506
rect 30545 24454 30557 24506
rect 30609 24454 30621 24506
rect 30673 24454 30685 24506
rect 30737 24454 30749 24506
rect 30801 24454 34868 24506
rect 1104 24432 34868 24454
rect 10042 24352 10048 24404
rect 10100 24392 10106 24404
rect 12526 24392 12532 24404
rect 10100 24364 10456 24392
rect 10100 24352 10106 24364
rect 10321 24327 10379 24333
rect 10321 24293 10333 24327
rect 10367 24293 10379 24327
rect 10321 24287 10379 24293
rect 8938 24148 8944 24200
rect 8996 24148 9002 24200
rect 10336 24188 10364 24287
rect 10428 24256 10456 24364
rect 12406 24364 12532 24392
rect 10502 24284 10508 24336
rect 10560 24324 10566 24336
rect 10686 24324 10692 24336
rect 10560 24296 10692 24324
rect 10560 24284 10566 24296
rect 10686 24284 10692 24296
rect 10744 24324 10750 24336
rect 12406 24324 12434 24364
rect 12526 24352 12532 24364
rect 12584 24352 12590 24404
rect 13170 24352 13176 24404
rect 13228 24352 13234 24404
rect 13817 24395 13875 24401
rect 13817 24361 13829 24395
rect 13863 24392 13875 24395
rect 13998 24392 14004 24404
rect 13863 24364 14004 24392
rect 13863 24361 13875 24364
rect 13817 24355 13875 24361
rect 13998 24352 14004 24364
rect 14056 24352 14062 24404
rect 14090 24352 14096 24404
rect 14148 24352 14154 24404
rect 14826 24352 14832 24404
rect 14884 24352 14890 24404
rect 15378 24352 15384 24404
rect 15436 24352 15442 24404
rect 18138 24352 18144 24404
rect 18196 24392 18202 24404
rect 18785 24395 18843 24401
rect 18785 24392 18797 24395
rect 18196 24364 18797 24392
rect 18196 24352 18202 24364
rect 18785 24361 18797 24364
rect 18831 24361 18843 24395
rect 18785 24355 18843 24361
rect 20254 24352 20260 24404
rect 20312 24392 20318 24404
rect 20349 24395 20407 24401
rect 20349 24392 20361 24395
rect 20312 24364 20361 24392
rect 20312 24352 20318 24364
rect 20349 24361 20361 24364
rect 20395 24361 20407 24395
rect 20349 24355 20407 24361
rect 20990 24352 20996 24404
rect 21048 24392 21054 24404
rect 21453 24395 21511 24401
rect 21453 24392 21465 24395
rect 21048 24364 21465 24392
rect 21048 24352 21054 24364
rect 21453 24361 21465 24364
rect 21499 24392 21511 24395
rect 22646 24392 22652 24404
rect 21499 24364 22652 24392
rect 21499 24361 21511 24364
rect 21453 24355 21511 24361
rect 22646 24352 22652 24364
rect 22704 24392 22710 24404
rect 22704 24364 22968 24392
rect 22704 24352 22710 24364
rect 10744 24296 12434 24324
rect 10744 24284 10750 24296
rect 11793 24259 11851 24265
rect 11793 24256 11805 24259
rect 10428 24228 11805 24256
rect 11793 24225 11805 24228
rect 11839 24225 11851 24259
rect 13188 24256 13216 24352
rect 13725 24327 13783 24333
rect 13725 24293 13737 24327
rect 13771 24324 13783 24327
rect 13771 24296 14044 24324
rect 13771 24293 13783 24296
rect 13725 24287 13783 24293
rect 14016 24268 14044 24296
rect 13909 24259 13967 24265
rect 13909 24256 13921 24259
rect 13188 24228 13921 24256
rect 11793 24219 11851 24225
rect 13909 24225 13921 24228
rect 13955 24225 13967 24259
rect 13909 24219 13967 24225
rect 13998 24216 14004 24268
rect 14056 24216 14062 24268
rect 10505 24191 10563 24197
rect 10505 24188 10517 24191
rect 10336 24160 10517 24188
rect 10505 24157 10517 24160
rect 10551 24157 10563 24191
rect 10505 24151 10563 24157
rect 12710 24148 12716 24200
rect 12768 24148 12774 24200
rect 12986 24148 12992 24200
rect 13044 24148 13050 24200
rect 13446 24148 13452 24200
rect 13504 24148 13510 24200
rect 13633 24191 13691 24197
rect 13633 24157 13645 24191
rect 13679 24157 13691 24191
rect 14108 24188 14136 24352
rect 14550 24284 14556 24336
rect 14608 24284 14614 24336
rect 14366 24216 14372 24268
rect 14424 24216 14430 24268
rect 14568 24256 14596 24284
rect 14844 24256 14872 24352
rect 14921 24259 14979 24265
rect 14921 24256 14933 24259
rect 14568 24228 14780 24256
rect 14844 24228 14933 24256
rect 14108 24160 14228 24188
rect 13633 24151 13691 24157
rect 9208 24123 9266 24129
rect 9208 24089 9220 24123
rect 9254 24120 9266 24123
rect 9306 24120 9312 24132
rect 9254 24092 9312 24120
rect 9254 24089 9266 24092
rect 9208 24083 9266 24089
rect 9306 24080 9312 24092
rect 9364 24080 9370 24132
rect 13004 24120 13032 24148
rect 13648 24120 13676 24151
rect 13004 24092 13676 24120
rect 13722 24080 13728 24132
rect 13780 24120 13786 24132
rect 14093 24123 14151 24129
rect 14093 24120 14105 24123
rect 13780 24092 14105 24120
rect 13780 24080 13786 24092
rect 14093 24089 14105 24092
rect 14139 24089 14151 24123
rect 14200 24120 14228 24160
rect 14274 24148 14280 24200
rect 14332 24148 14338 24200
rect 14384 24188 14412 24216
rect 14553 24191 14611 24197
rect 14553 24188 14565 24191
rect 14384 24160 14565 24188
rect 14553 24157 14565 24160
rect 14599 24157 14611 24191
rect 14752 24188 14780 24228
rect 14921 24225 14933 24228
rect 14967 24225 14979 24259
rect 15396 24256 15424 24352
rect 18598 24284 18604 24336
rect 18656 24324 18662 24336
rect 18877 24327 18935 24333
rect 18877 24324 18889 24327
rect 18656 24296 18889 24324
rect 18656 24284 18662 24296
rect 18877 24293 18889 24296
rect 18923 24324 18935 24327
rect 19150 24324 19156 24336
rect 18923 24296 19156 24324
rect 18923 24293 18935 24296
rect 18877 24287 18935 24293
rect 19150 24284 19156 24296
rect 19208 24284 19214 24336
rect 21726 24324 21732 24336
rect 19352 24296 21732 24324
rect 15565 24259 15623 24265
rect 15565 24256 15577 24259
rect 15396 24228 15577 24256
rect 14921 24219 14979 24225
rect 15565 24225 15577 24228
rect 15611 24225 15623 24259
rect 18616 24256 18644 24284
rect 15565 24219 15623 24225
rect 18432 24228 18644 24256
rect 15286 24188 15292 24200
rect 14752 24160 15292 24188
rect 14553 24151 14611 24157
rect 15286 24148 15292 24160
rect 15344 24188 15350 24200
rect 15473 24191 15531 24197
rect 15473 24188 15485 24191
rect 15344 24160 15485 24188
rect 15344 24148 15350 24160
rect 15473 24157 15485 24160
rect 15519 24157 15531 24191
rect 15473 24151 15531 24157
rect 17313 24191 17371 24197
rect 17313 24157 17325 24191
rect 17359 24188 17371 24191
rect 17678 24188 17684 24200
rect 17359 24160 17684 24188
rect 17359 24157 17371 24160
rect 17313 24151 17371 24157
rect 17678 24148 17684 24160
rect 17736 24148 17742 24200
rect 18432 24197 18460 24228
rect 18690 24216 18696 24268
rect 18748 24256 18754 24268
rect 19352 24256 19380 24296
rect 21726 24284 21732 24296
rect 21784 24284 21790 24336
rect 22554 24284 22560 24336
rect 22612 24324 22618 24336
rect 22741 24327 22799 24333
rect 22741 24324 22753 24327
rect 22612 24296 22753 24324
rect 22612 24284 22618 24296
rect 22741 24293 22753 24296
rect 22787 24293 22799 24327
rect 22741 24287 22799 24293
rect 18748 24228 19380 24256
rect 18748 24216 18754 24228
rect 19426 24216 19432 24268
rect 19484 24256 19490 24268
rect 19610 24256 19616 24268
rect 19484 24228 19616 24256
rect 19484 24216 19490 24228
rect 19610 24216 19616 24228
rect 19668 24256 19674 24268
rect 19889 24259 19947 24265
rect 19889 24256 19901 24259
rect 19668 24228 19901 24256
rect 19668 24216 19674 24228
rect 19889 24225 19901 24228
rect 19935 24225 19947 24259
rect 19889 24219 19947 24225
rect 21542 24216 21548 24268
rect 21600 24216 21606 24268
rect 22940 24265 22968 24364
rect 22925 24259 22983 24265
rect 22925 24225 22937 24259
rect 22971 24225 22983 24259
rect 22925 24219 22983 24225
rect 17957 24191 18015 24197
rect 17957 24157 17969 24191
rect 18003 24157 18015 24191
rect 17957 24151 18015 24157
rect 18417 24191 18475 24197
rect 18417 24157 18429 24191
rect 18463 24157 18475 24191
rect 18417 24151 18475 24157
rect 18601 24191 18659 24197
rect 18601 24157 18613 24191
rect 18647 24157 18659 24191
rect 18601 24151 18659 24157
rect 18969 24191 19027 24197
rect 18969 24157 18981 24191
rect 19015 24188 19027 24191
rect 20993 24191 21051 24197
rect 19015 24160 19380 24188
rect 19015 24157 19027 24160
rect 18969 24151 19027 24157
rect 14458 24120 14464 24132
rect 14200 24092 14464 24120
rect 14093 24083 14151 24089
rect 14458 24080 14464 24092
rect 14516 24080 14522 24132
rect 17068 24123 17126 24129
rect 17068 24089 17080 24123
rect 17114 24120 17126 24123
rect 17405 24123 17463 24129
rect 17405 24120 17417 24123
rect 17114 24092 17417 24120
rect 17114 24089 17126 24092
rect 17068 24083 17126 24089
rect 17405 24089 17417 24092
rect 17451 24089 17463 24123
rect 17405 24083 17463 24089
rect 17494 24080 17500 24132
rect 17552 24120 17558 24132
rect 17972 24120 18000 24151
rect 17552 24092 18000 24120
rect 18616 24120 18644 24151
rect 18984 24120 19012 24151
rect 18616 24092 19012 24120
rect 17552 24080 17558 24092
rect 11238 24012 11244 24064
rect 11296 24012 11302 24064
rect 12158 24012 12164 24064
rect 12216 24012 12222 24064
rect 12894 24012 12900 24064
rect 12952 24012 12958 24064
rect 13354 24012 13360 24064
rect 13412 24052 13418 24064
rect 15197 24055 15255 24061
rect 15197 24052 15209 24055
rect 13412 24024 15209 24052
rect 13412 24012 13418 24024
rect 15197 24021 15209 24024
rect 15243 24021 15255 24055
rect 15197 24015 15255 24021
rect 15470 24012 15476 24064
rect 15528 24052 15534 24064
rect 15930 24052 15936 24064
rect 15528 24024 15936 24052
rect 15528 24012 15534 24024
rect 15930 24012 15936 24024
rect 15988 24012 15994 24064
rect 18230 24012 18236 24064
rect 18288 24012 18294 24064
rect 19352 24061 19380 24160
rect 20993 24157 21005 24191
rect 21039 24188 21051 24191
rect 21085 24191 21143 24197
rect 21085 24188 21097 24191
rect 21039 24160 21097 24188
rect 21039 24157 21051 24160
rect 20993 24151 21051 24157
rect 21085 24157 21097 24160
rect 21131 24157 21143 24191
rect 21085 24151 21143 24157
rect 21266 24148 21272 24200
rect 21324 24148 21330 24200
rect 21818 24148 21824 24200
rect 21876 24188 21882 24200
rect 22189 24191 22247 24197
rect 22189 24188 22201 24191
rect 21876 24160 22201 24188
rect 21876 24148 21882 24160
rect 22189 24157 22201 24160
rect 22235 24157 22247 24191
rect 22373 24191 22431 24197
rect 22373 24188 22385 24191
rect 22189 24151 22247 24157
rect 22296 24160 22385 24188
rect 22296 24064 22324 24160
rect 22373 24157 22385 24160
rect 22419 24157 22431 24191
rect 22373 24151 22431 24157
rect 22557 24191 22615 24197
rect 22557 24157 22569 24191
rect 22603 24188 22615 24191
rect 22649 24191 22707 24197
rect 22649 24188 22661 24191
rect 22603 24160 22661 24188
rect 22603 24157 22615 24160
rect 22557 24151 22615 24157
rect 22649 24157 22661 24160
rect 22695 24157 22707 24191
rect 22649 24151 22707 24157
rect 23198 24148 23204 24200
rect 23256 24148 23262 24200
rect 25041 24191 25099 24197
rect 25041 24188 25053 24191
rect 24504 24160 25053 24188
rect 24504 24064 24532 24160
rect 25041 24157 25053 24160
rect 25087 24157 25099 24191
rect 25041 24151 25099 24157
rect 19337 24055 19395 24061
rect 19337 24021 19349 24055
rect 19383 24052 19395 24055
rect 19426 24052 19432 24064
rect 19383 24024 19432 24052
rect 19383 24021 19395 24024
rect 19337 24015 19395 24021
rect 19426 24012 19432 24024
rect 19484 24012 19490 24064
rect 22278 24012 22284 24064
rect 22336 24012 22342 24064
rect 22922 24012 22928 24064
rect 22980 24012 22986 24064
rect 23842 24012 23848 24064
rect 23900 24012 23906 24064
rect 24486 24012 24492 24064
rect 24544 24012 24550 24064
rect 24578 24012 24584 24064
rect 24636 24052 24642 24064
rect 24857 24055 24915 24061
rect 24857 24052 24869 24055
rect 24636 24024 24869 24052
rect 24636 24012 24642 24024
rect 24857 24021 24869 24024
rect 24903 24021 24915 24055
rect 24857 24015 24915 24021
rect 1104 23962 35027 23984
rect 1104 23910 9390 23962
rect 9442 23910 9454 23962
rect 9506 23910 9518 23962
rect 9570 23910 9582 23962
rect 9634 23910 9646 23962
rect 9698 23910 17831 23962
rect 17883 23910 17895 23962
rect 17947 23910 17959 23962
rect 18011 23910 18023 23962
rect 18075 23910 18087 23962
rect 18139 23910 26272 23962
rect 26324 23910 26336 23962
rect 26388 23910 26400 23962
rect 26452 23910 26464 23962
rect 26516 23910 26528 23962
rect 26580 23910 34713 23962
rect 34765 23910 34777 23962
rect 34829 23910 34841 23962
rect 34893 23910 34905 23962
rect 34957 23910 34969 23962
rect 35021 23910 35027 23962
rect 1104 23888 35027 23910
rect 9306 23808 9312 23860
rect 9364 23848 9370 23860
rect 9769 23851 9827 23857
rect 9769 23848 9781 23851
rect 9364 23820 9781 23848
rect 9364 23808 9370 23820
rect 9769 23817 9781 23820
rect 9815 23817 9827 23851
rect 9769 23811 9827 23817
rect 10597 23851 10655 23857
rect 10597 23817 10609 23851
rect 10643 23848 10655 23851
rect 11146 23848 11152 23860
rect 10643 23820 11152 23848
rect 10643 23817 10655 23820
rect 10597 23811 10655 23817
rect 11146 23808 11152 23820
rect 11204 23808 11210 23860
rect 11238 23808 11244 23860
rect 11296 23808 11302 23860
rect 11514 23808 11520 23860
rect 11572 23808 11578 23860
rect 11698 23808 11704 23860
rect 11756 23808 11762 23860
rect 12253 23851 12311 23857
rect 12253 23817 12265 23851
rect 12299 23848 12311 23851
rect 12710 23848 12716 23860
rect 12299 23820 12716 23848
rect 12299 23817 12311 23820
rect 12253 23811 12311 23817
rect 12710 23808 12716 23820
rect 12768 23808 12774 23860
rect 12805 23851 12863 23857
rect 12805 23817 12817 23851
rect 12851 23848 12863 23851
rect 13446 23848 13452 23860
rect 12851 23820 13452 23848
rect 12851 23817 12863 23820
rect 12805 23811 12863 23817
rect 13446 23808 13452 23820
rect 13504 23808 13510 23860
rect 13722 23808 13728 23860
rect 13780 23808 13786 23860
rect 14274 23808 14280 23860
rect 14332 23808 14338 23860
rect 14458 23808 14464 23860
rect 14516 23808 14522 23860
rect 14642 23808 14648 23860
rect 14700 23808 14706 23860
rect 14826 23808 14832 23860
rect 14884 23848 14890 23860
rect 15105 23851 15163 23857
rect 15105 23848 15117 23851
rect 14884 23820 15117 23848
rect 14884 23808 14890 23820
rect 15105 23817 15117 23820
rect 15151 23848 15163 23851
rect 15489 23851 15547 23857
rect 15489 23848 15501 23851
rect 15151 23820 15501 23848
rect 15151 23817 15163 23820
rect 15105 23811 15163 23817
rect 15489 23817 15501 23820
rect 15535 23817 15547 23851
rect 15489 23811 15547 23817
rect 15654 23808 15660 23860
rect 15712 23808 15718 23860
rect 15746 23808 15752 23860
rect 15804 23808 15810 23860
rect 15838 23808 15844 23860
rect 15896 23848 15902 23860
rect 15896 23820 16068 23848
rect 15896 23808 15902 23820
rect 11256 23780 11284 23808
rect 9692 23752 11284 23780
rect 11532 23780 11560 23808
rect 11716 23780 11744 23808
rect 13740 23780 13768 23808
rect 11532 23752 11652 23780
rect 11716 23752 11928 23780
rect 9692 23721 9720 23752
rect 9677 23715 9735 23721
rect 9677 23681 9689 23715
rect 9723 23681 9735 23715
rect 9677 23675 9735 23681
rect 9861 23715 9919 23721
rect 9861 23681 9873 23715
rect 9907 23681 9919 23715
rect 9861 23675 9919 23681
rect 10229 23715 10287 23721
rect 10229 23681 10241 23715
rect 10275 23712 10287 23715
rect 10275 23684 10732 23712
rect 10275 23681 10287 23684
rect 10229 23675 10287 23681
rect 9876 23576 9904 23675
rect 10134 23604 10140 23656
rect 10192 23604 10198 23656
rect 10704 23585 10732 23684
rect 11514 23672 11520 23724
rect 11572 23672 11578 23724
rect 11624 23712 11652 23752
rect 11701 23715 11759 23721
rect 11701 23712 11713 23715
rect 11624 23684 11713 23712
rect 11701 23681 11713 23684
rect 11747 23681 11759 23715
rect 11701 23675 11759 23681
rect 11793 23715 11851 23721
rect 11793 23681 11805 23715
rect 11839 23714 11851 23715
rect 11900 23714 11928 23752
rect 13280 23752 13768 23780
rect 14476 23780 14504 23808
rect 14660 23780 14688 23808
rect 14476 23752 14596 23780
rect 11839 23686 11928 23714
rect 12069 23715 12127 23721
rect 11839 23681 11851 23686
rect 11793 23675 11851 23681
rect 12069 23681 12081 23715
rect 12115 23712 12127 23715
rect 12115 23684 12204 23712
rect 12115 23681 12127 23684
rect 12069 23675 12127 23681
rect 11238 23604 11244 23656
rect 11296 23604 11302 23656
rect 11882 23604 11888 23656
rect 11940 23604 11946 23656
rect 10689 23579 10747 23585
rect 9876 23548 10640 23576
rect 10612 23508 10640 23548
rect 10689 23545 10701 23579
rect 10735 23576 10747 23579
rect 12176 23576 12204 23684
rect 12986 23672 12992 23724
rect 13044 23712 13050 23724
rect 13081 23715 13139 23721
rect 13081 23712 13093 23715
rect 13044 23684 13093 23712
rect 13044 23672 13050 23684
rect 13081 23681 13093 23684
rect 13127 23681 13139 23715
rect 13081 23675 13139 23681
rect 13170 23672 13176 23724
rect 13228 23672 13234 23724
rect 13280 23721 13308 23752
rect 13265 23715 13323 23721
rect 13265 23681 13277 23715
rect 13311 23681 13323 23715
rect 13265 23675 13323 23681
rect 13449 23715 13507 23721
rect 13449 23681 13461 23715
rect 13495 23712 13507 23715
rect 13722 23712 13728 23724
rect 13495 23684 13728 23712
rect 13495 23681 13507 23684
rect 13449 23675 13507 23681
rect 13722 23672 13728 23684
rect 13780 23672 13786 23724
rect 14182 23672 14188 23724
rect 14240 23672 14246 23724
rect 14366 23672 14372 23724
rect 14424 23712 14430 23724
rect 14568 23721 14596 23752
rect 14659 23752 14688 23780
rect 14659 23721 14687 23752
rect 15286 23740 15292 23792
rect 15344 23740 15350 23792
rect 15764 23780 15792 23808
rect 15764 23752 15976 23780
rect 14461 23715 14519 23721
rect 14461 23712 14473 23715
rect 14424 23684 14473 23712
rect 14424 23672 14430 23684
rect 14461 23681 14473 23684
rect 14507 23681 14519 23715
rect 14461 23675 14519 23681
rect 14553 23715 14611 23721
rect 14553 23681 14565 23715
rect 14599 23681 14611 23715
rect 14553 23675 14611 23681
rect 14645 23715 14703 23721
rect 14645 23681 14657 23715
rect 14691 23681 14703 23715
rect 14645 23675 14703 23681
rect 10735 23548 12204 23576
rect 13004 23576 13032 23672
rect 14277 23647 14335 23653
rect 14277 23613 14289 23647
rect 14323 23644 14335 23647
rect 14659 23644 14687 23675
rect 14734 23672 14740 23724
rect 14792 23672 14798 23724
rect 14918 23672 14924 23724
rect 14976 23672 14982 23724
rect 15013 23715 15071 23721
rect 15013 23681 15025 23715
rect 15059 23712 15071 23715
rect 15102 23712 15108 23724
rect 15059 23684 15108 23712
rect 15059 23681 15071 23684
rect 15013 23675 15071 23681
rect 15102 23672 15108 23684
rect 15160 23672 15166 23724
rect 15197 23715 15255 23721
rect 15197 23681 15209 23715
rect 15243 23681 15255 23715
rect 15197 23675 15255 23681
rect 14323 23616 14687 23644
rect 15212 23644 15240 23675
rect 15562 23672 15568 23724
rect 15620 23712 15626 23724
rect 15948 23721 15976 23752
rect 16040 23721 16068 23820
rect 16114 23808 16120 23860
rect 16172 23808 16178 23860
rect 16393 23851 16451 23857
rect 16393 23817 16405 23851
rect 16439 23848 16451 23851
rect 17494 23848 17500 23860
rect 16439 23820 17500 23848
rect 16439 23817 16451 23820
rect 16393 23811 16451 23817
rect 17494 23808 17500 23820
rect 17552 23808 17558 23860
rect 18322 23808 18328 23860
rect 18380 23808 18386 23860
rect 19610 23808 19616 23860
rect 19668 23808 19674 23860
rect 19794 23808 19800 23860
rect 19852 23808 19858 23860
rect 22281 23851 22339 23857
rect 22281 23817 22293 23851
rect 22327 23848 22339 23851
rect 22370 23848 22376 23860
rect 22327 23820 22376 23848
rect 22327 23817 22339 23820
rect 22281 23811 22339 23817
rect 22370 23808 22376 23820
rect 22428 23808 22434 23860
rect 22462 23808 22468 23860
rect 22520 23808 22526 23860
rect 22922 23808 22928 23860
rect 22980 23808 22986 23860
rect 23017 23851 23075 23857
rect 23017 23817 23029 23851
rect 23063 23848 23075 23851
rect 23198 23848 23204 23860
rect 23063 23820 23204 23848
rect 23063 23817 23075 23820
rect 23017 23811 23075 23817
rect 23198 23808 23204 23820
rect 23256 23808 23262 23860
rect 23842 23808 23848 23860
rect 23900 23808 23906 23860
rect 16132 23721 16160 23808
rect 18340 23780 18368 23808
rect 18478 23783 18536 23789
rect 18478 23780 18490 23783
rect 18340 23752 18490 23780
rect 18478 23749 18490 23752
rect 18524 23749 18536 23783
rect 19812 23780 19840 23808
rect 20073 23783 20131 23789
rect 20073 23780 20085 23783
rect 19812 23752 20085 23780
rect 18478 23743 18536 23749
rect 20073 23749 20085 23752
rect 20119 23749 20131 23783
rect 20073 23743 20131 23749
rect 15749 23715 15807 23721
rect 15749 23712 15761 23715
rect 15620 23684 15761 23712
rect 15620 23672 15626 23684
rect 15749 23681 15761 23684
rect 15795 23681 15807 23715
rect 15749 23675 15807 23681
rect 15933 23715 15991 23721
rect 15933 23681 15945 23715
rect 15979 23681 15991 23715
rect 15933 23675 15991 23681
rect 16025 23715 16083 23721
rect 16025 23681 16037 23715
rect 16071 23681 16083 23715
rect 16025 23675 16083 23681
rect 16117 23715 16175 23721
rect 16117 23681 16129 23715
rect 16163 23681 16175 23715
rect 16117 23675 16175 23681
rect 17028 23715 17086 23721
rect 17028 23681 17040 23715
rect 17074 23712 17086 23715
rect 17310 23712 17316 23724
rect 17074 23684 17316 23712
rect 17074 23681 17086 23684
rect 17028 23675 17086 23681
rect 16132 23644 16160 23675
rect 17310 23672 17316 23684
rect 17368 23672 17374 23724
rect 19610 23672 19616 23724
rect 19668 23712 19674 23724
rect 19889 23715 19947 23721
rect 19889 23712 19901 23715
rect 19668 23684 19901 23712
rect 19668 23672 19674 23684
rect 19889 23681 19901 23684
rect 19935 23681 19947 23715
rect 19889 23675 19947 23681
rect 19981 23715 20039 23721
rect 19981 23681 19993 23715
rect 20027 23681 20039 23715
rect 19981 23675 20039 23681
rect 15212 23616 16160 23644
rect 16761 23647 16819 23653
rect 14323 23613 14335 23616
rect 14277 23607 14335 23613
rect 16761 23613 16773 23647
rect 16807 23613 16819 23647
rect 16761 23607 16819 23613
rect 18233 23647 18291 23653
rect 18233 23613 18245 23647
rect 18279 23613 18291 23647
rect 19996 23644 20024 23675
rect 20162 23672 20168 23724
rect 20220 23712 20226 23724
rect 20257 23715 20315 23721
rect 20257 23712 20269 23715
rect 20220 23684 20269 23712
rect 20220 23672 20226 23684
rect 20257 23681 20269 23684
rect 20303 23681 20315 23715
rect 20257 23675 20315 23681
rect 22097 23715 22155 23721
rect 22097 23681 22109 23715
rect 22143 23681 22155 23715
rect 22097 23675 22155 23681
rect 22373 23715 22431 23721
rect 22373 23681 22385 23715
rect 22419 23712 22431 23715
rect 22480 23712 22508 23808
rect 22940 23780 22968 23808
rect 22572 23752 22968 23780
rect 23376 23783 23434 23789
rect 22572 23721 22600 23752
rect 23376 23749 23388 23783
rect 23422 23780 23434 23783
rect 23860 23780 23888 23808
rect 23422 23752 23888 23780
rect 23422 23749 23434 23752
rect 23376 23743 23434 23749
rect 22419 23684 22508 23712
rect 22557 23715 22615 23721
rect 22419 23681 22431 23684
rect 22373 23675 22431 23681
rect 22557 23681 22569 23715
rect 22603 23681 22615 23715
rect 22557 23675 22615 23681
rect 18233 23607 18291 23613
rect 19904 23616 20024 23644
rect 13541 23579 13599 23585
rect 13541 23576 13553 23579
rect 13004 23548 13553 23576
rect 10735 23545 10747 23548
rect 10689 23539 10747 23545
rect 13541 23545 13553 23548
rect 13587 23545 13599 23579
rect 13541 23539 13599 23545
rect 15378 23536 15384 23588
rect 15436 23576 15442 23588
rect 15436 23548 15516 23576
rect 15436 23536 15442 23548
rect 11054 23508 11060 23520
rect 10612 23480 11060 23508
rect 11054 23468 11060 23480
rect 11112 23468 11118 23520
rect 11882 23468 11888 23520
rect 11940 23508 11946 23520
rect 13170 23508 13176 23520
rect 11940 23480 13176 23508
rect 11940 23468 11946 23480
rect 13170 23468 13176 23480
rect 13228 23508 13234 23520
rect 14458 23508 14464 23520
rect 13228 23480 14464 23508
rect 13228 23468 13234 23480
rect 14458 23468 14464 23480
rect 14516 23468 14522 23520
rect 14642 23468 14648 23520
rect 14700 23508 14706 23520
rect 15488 23517 15516 23548
rect 14921 23511 14979 23517
rect 14921 23508 14933 23511
rect 14700 23480 14933 23508
rect 14700 23468 14706 23480
rect 14921 23477 14933 23480
rect 14967 23477 14979 23511
rect 14921 23471 14979 23477
rect 15464 23511 15522 23517
rect 15464 23477 15476 23511
rect 15510 23477 15522 23511
rect 16776 23508 16804 23607
rect 18248 23576 18276 23607
rect 17696 23548 18276 23576
rect 17696 23520 17724 23548
rect 19904 23520 19932 23616
rect 21634 23604 21640 23656
rect 21692 23644 21698 23656
rect 21821 23647 21879 23653
rect 21821 23644 21833 23647
rect 21692 23616 21833 23644
rect 21692 23604 21698 23616
rect 21821 23613 21833 23616
rect 21867 23613 21879 23647
rect 22112 23644 22140 23675
rect 22646 23672 22652 23724
rect 22704 23672 22710 23724
rect 22741 23715 22799 23721
rect 22741 23681 22753 23715
rect 22787 23712 22799 23715
rect 23658 23712 23664 23724
rect 22787 23684 23664 23712
rect 22787 23681 22799 23684
rect 22741 23675 22799 23681
rect 23658 23672 23664 23684
rect 23716 23712 23722 23724
rect 24578 23712 24584 23724
rect 23716 23684 24584 23712
rect 23716 23672 23722 23684
rect 24578 23672 24584 23684
rect 24636 23672 24642 23724
rect 22462 23644 22468 23656
rect 22112 23616 22468 23644
rect 21821 23607 21879 23613
rect 22462 23604 22468 23616
rect 22520 23604 22526 23656
rect 22830 23604 22836 23656
rect 22888 23644 22894 23656
rect 23109 23647 23167 23653
rect 23109 23644 23121 23647
rect 22888 23616 23121 23644
rect 22888 23604 22894 23616
rect 23109 23613 23121 23616
rect 23155 23613 23167 23647
rect 23109 23607 23167 23613
rect 21913 23579 21971 23585
rect 21913 23545 21925 23579
rect 21959 23576 21971 23579
rect 21959 23548 22094 23576
rect 21959 23545 21971 23548
rect 21913 23539 21971 23545
rect 17678 23508 17684 23520
rect 16776 23480 17684 23508
rect 15464 23471 15522 23477
rect 17678 23468 17684 23480
rect 17736 23468 17742 23520
rect 18141 23511 18199 23517
rect 18141 23477 18153 23511
rect 18187 23508 18199 23511
rect 18230 23508 18236 23520
rect 18187 23480 18236 23508
rect 18187 23477 18199 23480
rect 18141 23471 18199 23477
rect 18230 23468 18236 23480
rect 18288 23468 18294 23520
rect 19702 23468 19708 23520
rect 19760 23468 19766 23520
rect 19886 23468 19892 23520
rect 19944 23468 19950 23520
rect 22066 23508 22094 23548
rect 22554 23508 22560 23520
rect 22066 23480 22560 23508
rect 22554 23468 22560 23480
rect 22612 23468 22618 23520
rect 24486 23468 24492 23520
rect 24544 23468 24550 23520
rect 1104 23418 34868 23440
rect 1104 23366 5170 23418
rect 5222 23366 5234 23418
rect 5286 23366 5298 23418
rect 5350 23366 5362 23418
rect 5414 23366 5426 23418
rect 5478 23366 13611 23418
rect 13663 23366 13675 23418
rect 13727 23366 13739 23418
rect 13791 23366 13803 23418
rect 13855 23366 13867 23418
rect 13919 23366 22052 23418
rect 22104 23366 22116 23418
rect 22168 23366 22180 23418
rect 22232 23366 22244 23418
rect 22296 23366 22308 23418
rect 22360 23366 30493 23418
rect 30545 23366 30557 23418
rect 30609 23366 30621 23418
rect 30673 23366 30685 23418
rect 30737 23366 30749 23418
rect 30801 23366 34868 23418
rect 1104 23344 34868 23366
rect 10594 23264 10600 23316
rect 10652 23264 10658 23316
rect 11057 23307 11115 23313
rect 11057 23273 11069 23307
rect 11103 23304 11115 23307
rect 11238 23304 11244 23316
rect 11103 23276 11244 23304
rect 11103 23273 11115 23276
rect 11057 23267 11115 23273
rect 11238 23264 11244 23276
rect 11296 23264 11302 23316
rect 13909 23307 13967 23313
rect 13909 23273 13921 23307
rect 13955 23304 13967 23307
rect 14182 23304 14188 23316
rect 13955 23276 14188 23304
rect 13955 23273 13967 23276
rect 13909 23267 13967 23273
rect 14182 23264 14188 23276
rect 14240 23264 14246 23316
rect 14458 23264 14464 23316
rect 14516 23264 14522 23316
rect 17310 23264 17316 23316
rect 17368 23264 17374 23316
rect 19426 23264 19432 23316
rect 19484 23264 19490 23316
rect 19518 23264 19524 23316
rect 19576 23304 19582 23316
rect 19613 23307 19671 23313
rect 19613 23304 19625 23307
rect 19576 23276 19625 23304
rect 19576 23264 19582 23276
rect 19613 23273 19625 23276
rect 19659 23273 19671 23307
rect 19613 23267 19671 23273
rect 22186 23264 22192 23316
rect 22244 23304 22250 23316
rect 22462 23304 22468 23316
rect 22244 23276 22468 23304
rect 22244 23264 22250 23276
rect 22462 23264 22468 23276
rect 22520 23264 22526 23316
rect 22554 23264 22560 23316
rect 22612 23313 22618 23316
rect 22612 23307 22661 23313
rect 22612 23273 22615 23307
rect 22649 23304 22661 23307
rect 22649 23276 24440 23304
rect 22649 23273 22661 23276
rect 22612 23267 22661 23273
rect 22612 23264 22618 23267
rect 14090 23196 14096 23248
rect 14148 23236 14154 23248
rect 15010 23236 15016 23248
rect 14148 23208 15016 23236
rect 14148 23196 14154 23208
rect 15010 23196 15016 23208
rect 15068 23196 15074 23248
rect 17129 23239 17187 23245
rect 17129 23205 17141 23239
rect 17175 23236 17187 23239
rect 18138 23236 18144 23248
rect 17175 23208 18144 23236
rect 17175 23205 17187 23208
rect 17129 23199 17187 23205
rect 18138 23196 18144 23208
rect 18196 23196 18202 23248
rect 21545 23239 21603 23245
rect 21545 23205 21557 23239
rect 21591 23236 21603 23239
rect 21634 23236 21640 23248
rect 21591 23208 21640 23236
rect 21591 23205 21603 23208
rect 21545 23199 21603 23205
rect 21634 23196 21640 23208
rect 21692 23236 21698 23248
rect 21692 23208 22232 23236
rect 21692 23196 21698 23208
rect 14369 23171 14427 23177
rect 14369 23137 14381 23171
rect 14415 23168 14427 23171
rect 14734 23168 14740 23180
rect 14415 23140 14740 23168
rect 14415 23137 14427 23140
rect 14369 23131 14427 23137
rect 14734 23128 14740 23140
rect 14792 23168 14798 23180
rect 15749 23171 15807 23177
rect 15749 23168 15761 23171
rect 14792 23140 15761 23168
rect 14792 23128 14798 23140
rect 15749 23137 15761 23140
rect 15795 23137 15807 23171
rect 15749 23131 15807 23137
rect 16761 23171 16819 23177
rect 16761 23137 16773 23171
rect 16807 23168 16819 23171
rect 17865 23171 17923 23177
rect 17865 23168 17877 23171
rect 16807 23140 17877 23168
rect 16807 23137 16819 23140
rect 16761 23131 16819 23137
rect 17865 23137 17877 23140
rect 17911 23137 17923 23171
rect 17865 23131 17923 23137
rect 18230 23128 18236 23180
rect 18288 23168 18294 23180
rect 19610 23168 19616 23180
rect 18288 23140 19616 23168
rect 18288 23128 18294 23140
rect 19610 23128 19616 23140
rect 19668 23128 19674 23180
rect 21177 23171 21235 23177
rect 21177 23137 21189 23171
rect 21223 23168 21235 23171
rect 21223 23140 21588 23168
rect 21223 23137 21235 23140
rect 21177 23131 21235 23137
rect 21560 23112 21588 23140
rect 21910 23128 21916 23180
rect 21968 23128 21974 23180
rect 10686 23060 10692 23112
rect 10744 23060 10750 23112
rect 12158 23060 12164 23112
rect 12216 23109 12222 23112
rect 12216 23100 12228 23109
rect 12437 23103 12495 23109
rect 12216 23072 12261 23100
rect 12216 23063 12228 23072
rect 12437 23069 12449 23103
rect 12483 23100 12495 23103
rect 12526 23100 12532 23112
rect 12483 23072 12532 23100
rect 12483 23069 12495 23072
rect 12437 23063 12495 23069
rect 12216 23060 12222 23063
rect 12526 23060 12532 23072
rect 12584 23100 12590 23112
rect 13538 23100 13544 23112
rect 12584 23072 13544 23100
rect 12584 23060 12590 23072
rect 13538 23060 13544 23072
rect 13596 23060 13602 23112
rect 14642 23060 14648 23112
rect 14700 23060 14706 23112
rect 14829 23103 14887 23109
rect 14829 23069 14841 23103
rect 14875 23100 14887 23103
rect 14921 23103 14979 23109
rect 14921 23100 14933 23103
rect 14875 23072 14933 23100
rect 14875 23069 14887 23072
rect 14829 23063 14887 23069
rect 14921 23069 14933 23072
rect 14967 23069 14979 23103
rect 14921 23063 14979 23069
rect 15286 23060 15292 23112
rect 15344 23100 15350 23112
rect 16114 23100 16120 23112
rect 15344 23072 16120 23100
rect 15344 23060 15350 23072
rect 16114 23060 16120 23072
rect 16172 23100 16178 23112
rect 16301 23103 16359 23109
rect 16301 23100 16313 23103
rect 16172 23072 16313 23100
rect 16172 23060 16178 23072
rect 16301 23069 16313 23072
rect 16347 23069 16359 23103
rect 16301 23063 16359 23069
rect 16945 23103 17003 23109
rect 16945 23069 16957 23103
rect 16991 23100 17003 23103
rect 17034 23100 17040 23112
rect 16991 23072 17040 23100
rect 16991 23069 17003 23072
rect 16945 23063 17003 23069
rect 17034 23060 17040 23072
rect 17092 23060 17098 23112
rect 17221 23103 17279 23109
rect 17221 23069 17233 23103
rect 17267 23069 17279 23103
rect 17221 23063 17279 23069
rect 12796 23035 12854 23041
rect 12796 23001 12808 23035
rect 12842 23032 12854 23035
rect 12894 23032 12900 23044
rect 12842 23004 12900 23032
rect 12842 23001 12854 23004
rect 12796 22995 12854 23001
rect 12894 22992 12900 23004
rect 12952 22992 12958 23044
rect 17236 23032 17264 23063
rect 17402 23060 17408 23112
rect 17460 23100 17466 23112
rect 18877 23103 18935 23109
rect 18877 23100 18889 23103
rect 17460 23072 18889 23100
rect 17460 23060 17466 23072
rect 18877 23069 18889 23072
rect 18923 23069 18935 23103
rect 18877 23063 18935 23069
rect 19058 23060 19064 23112
rect 19116 23060 19122 23112
rect 19150 23060 19156 23112
rect 19208 23100 19214 23112
rect 19208 23072 19380 23100
rect 19208 23060 19214 23072
rect 18785 23035 18843 23041
rect 18785 23032 18797 23035
rect 17236 23004 18797 23032
rect 18785 23001 18797 23004
rect 18831 23032 18843 23035
rect 19245 23035 19303 23041
rect 19245 23032 19257 23035
rect 18831 23004 19257 23032
rect 18831 23001 18843 23004
rect 18785 22995 18843 23001
rect 19245 23001 19257 23004
rect 19291 23001 19303 23035
rect 19352 23032 19380 23072
rect 20530 23060 20536 23112
rect 20588 23060 20594 23112
rect 21358 23060 21364 23112
rect 21416 23060 21422 23112
rect 21542 23060 21548 23112
rect 21600 23060 21606 23112
rect 21818 23060 21824 23112
rect 21876 23060 21882 23112
rect 22002 23060 22008 23112
rect 22060 23060 22066 23112
rect 22097 23103 22155 23109
rect 22097 23069 22109 23103
rect 22143 23069 22155 23103
rect 22097 23063 22155 23069
rect 19445 23035 19503 23041
rect 19445 23032 19457 23035
rect 19352 23004 19457 23032
rect 19245 22995 19303 23001
rect 19445 23001 19457 23004
rect 19491 23001 19503 23035
rect 19445 22995 19503 23001
rect 15562 22924 15568 22976
rect 15620 22924 15626 22976
rect 18230 22924 18236 22976
rect 18288 22964 18294 22976
rect 18969 22967 19027 22973
rect 18969 22964 18981 22967
rect 18288 22936 18981 22964
rect 18288 22924 18294 22936
rect 18969 22933 18981 22936
rect 19015 22933 19027 22967
rect 18969 22927 19027 22933
rect 19886 22924 19892 22976
rect 19944 22964 19950 22976
rect 20441 22967 20499 22973
rect 20441 22964 20453 22967
rect 19944 22936 20453 22964
rect 19944 22924 19950 22936
rect 20441 22933 20453 22936
rect 20487 22933 20499 22967
rect 20441 22927 20499 22933
rect 21634 22924 21640 22976
rect 21692 22924 21698 22976
rect 21836 22964 21864 23060
rect 21910 22992 21916 23044
rect 21968 23032 21974 23044
rect 22112 23032 22140 23063
rect 21968 23004 22140 23032
rect 22204 23032 22232 23208
rect 24412 23180 24440 23276
rect 23014 23128 23020 23180
rect 23072 23168 23078 23180
rect 23072 23140 24072 23168
rect 23072 23128 23078 23140
rect 22281 23103 22339 23109
rect 22281 23069 22293 23103
rect 22327 23102 22339 23103
rect 22327 23100 22416 23102
rect 22462 23100 22468 23112
rect 22327 23074 22468 23100
rect 22327 23072 22347 23074
rect 22388 23072 22468 23074
rect 22327 23069 22339 23072
rect 22281 23063 22339 23069
rect 22462 23060 22468 23072
rect 22520 23060 22526 23112
rect 22741 23103 22799 23109
rect 22741 23100 22753 23103
rect 22572 23072 22753 23100
rect 22572 23032 22600 23072
rect 22741 23069 22753 23072
rect 22787 23100 22799 23103
rect 22787 23072 22876 23100
rect 22787 23069 22799 23072
rect 22741 23063 22799 23069
rect 22204 23004 22600 23032
rect 22848 23032 22876 23072
rect 22922 23060 22928 23112
rect 22980 23060 22986 23112
rect 23661 23035 23719 23041
rect 23661 23032 23673 23035
rect 22848 23004 23673 23032
rect 21968 22992 21974 23004
rect 23661 23001 23673 23004
rect 23707 23001 23719 23035
rect 23661 22995 23719 23001
rect 23842 22992 23848 23044
rect 23900 22992 23906 23044
rect 22278 22964 22284 22976
rect 21836 22936 22284 22964
rect 22278 22924 22284 22936
rect 22336 22924 22342 22976
rect 22373 22967 22431 22973
rect 22373 22933 22385 22967
rect 22419 22964 22431 22967
rect 22554 22964 22560 22976
rect 22419 22936 22560 22964
rect 22419 22933 22431 22936
rect 22373 22927 22431 22933
rect 22554 22924 22560 22936
rect 22612 22924 22618 22976
rect 23290 22924 23296 22976
rect 23348 22964 23354 22976
rect 24044 22973 24072 23140
rect 24394 23128 24400 23180
rect 24452 23128 24458 23180
rect 25041 23103 25099 23109
rect 25041 23100 25053 23103
rect 24228 23072 25053 23100
rect 24228 22976 24256 23072
rect 25041 23069 25053 23072
rect 25087 23069 25099 23103
rect 25041 23063 25099 23069
rect 23569 22967 23627 22973
rect 23569 22964 23581 22967
rect 23348 22936 23581 22964
rect 23348 22924 23354 22936
rect 23569 22933 23581 22936
rect 23615 22933 23627 22967
rect 23569 22927 23627 22933
rect 24029 22967 24087 22973
rect 24029 22933 24041 22967
rect 24075 22964 24087 22967
rect 24118 22964 24124 22976
rect 24075 22936 24124 22964
rect 24075 22933 24087 22936
rect 24029 22927 24087 22933
rect 24118 22924 24124 22936
rect 24176 22924 24182 22976
rect 24210 22924 24216 22976
rect 24268 22924 24274 22976
rect 24302 22924 24308 22976
rect 24360 22964 24366 22976
rect 24857 22967 24915 22973
rect 24857 22964 24869 22967
rect 24360 22936 24869 22964
rect 24360 22924 24366 22936
rect 24857 22933 24869 22936
rect 24903 22933 24915 22967
rect 24857 22927 24915 22933
rect 1104 22874 35027 22896
rect 1104 22822 9390 22874
rect 9442 22822 9454 22874
rect 9506 22822 9518 22874
rect 9570 22822 9582 22874
rect 9634 22822 9646 22874
rect 9698 22822 17831 22874
rect 17883 22822 17895 22874
rect 17947 22822 17959 22874
rect 18011 22822 18023 22874
rect 18075 22822 18087 22874
rect 18139 22822 26272 22874
rect 26324 22822 26336 22874
rect 26388 22822 26400 22874
rect 26452 22822 26464 22874
rect 26516 22822 26528 22874
rect 26580 22822 34713 22874
rect 34765 22822 34777 22874
rect 34829 22822 34841 22874
rect 34893 22822 34905 22874
rect 34957 22822 34969 22874
rect 35021 22822 35027 22874
rect 1104 22800 35027 22822
rect 11238 22720 11244 22772
rect 11296 22720 11302 22772
rect 14182 22760 14188 22772
rect 13372 22732 14188 22760
rect 9030 22652 9036 22704
rect 9088 22692 9094 22704
rect 9088 22664 10180 22692
rect 9088 22652 9094 22664
rect 9858 22584 9864 22636
rect 9916 22584 9922 22636
rect 10152 22633 10180 22664
rect 11256 22633 11284 22720
rect 10045 22627 10103 22633
rect 10045 22593 10057 22627
rect 10091 22593 10103 22627
rect 10045 22587 10103 22593
rect 10137 22627 10195 22633
rect 10137 22593 10149 22627
rect 10183 22593 10195 22627
rect 10137 22587 10195 22593
rect 11241 22627 11299 22633
rect 11241 22593 11253 22627
rect 11287 22593 11299 22627
rect 11241 22587 11299 22593
rect 12621 22627 12679 22633
rect 12621 22593 12633 22627
rect 12667 22624 12679 22627
rect 12802 22624 12808 22636
rect 12667 22596 12808 22624
rect 12667 22593 12679 22596
rect 12621 22587 12679 22593
rect 10060 22556 10088 22587
rect 12802 22584 12808 22596
rect 12860 22584 12866 22636
rect 13078 22584 13084 22636
rect 13136 22584 13142 22636
rect 13372 22633 13400 22732
rect 14182 22720 14188 22732
rect 14240 22720 14246 22772
rect 14550 22720 14556 22772
rect 14608 22720 14614 22772
rect 15470 22760 15476 22772
rect 14660 22732 15476 22760
rect 13446 22652 13452 22704
rect 13504 22692 13510 22704
rect 13504 22664 13768 22692
rect 13504 22652 13510 22664
rect 13740 22633 13768 22664
rect 13357 22627 13415 22633
rect 13357 22593 13369 22627
rect 13403 22593 13415 22627
rect 13357 22587 13415 22593
rect 13725 22627 13783 22633
rect 13725 22593 13737 22627
rect 13771 22593 13783 22627
rect 13725 22587 13783 22593
rect 14090 22584 14096 22636
rect 14148 22584 14154 22636
rect 14369 22627 14427 22633
rect 14369 22593 14381 22627
rect 14415 22624 14427 22627
rect 14568 22624 14596 22720
rect 14660 22633 14688 22732
rect 15470 22720 15476 22732
rect 15528 22720 15534 22772
rect 15562 22720 15568 22772
rect 15620 22720 15626 22772
rect 16114 22720 16120 22772
rect 16172 22720 16178 22772
rect 17405 22763 17463 22769
rect 17405 22729 17417 22763
rect 17451 22729 17463 22763
rect 17405 22723 17463 22729
rect 15004 22695 15062 22701
rect 15004 22661 15016 22695
rect 15050 22692 15062 22695
rect 15580 22692 15608 22720
rect 15050 22664 15608 22692
rect 16209 22695 16267 22701
rect 15050 22661 15062 22664
rect 15004 22655 15062 22661
rect 16209 22661 16221 22695
rect 16255 22661 16267 22695
rect 17420 22692 17448 22723
rect 19702 22720 19708 22772
rect 19760 22720 19766 22772
rect 21545 22763 21603 22769
rect 21545 22729 21557 22763
rect 21591 22760 21603 22763
rect 22002 22760 22008 22772
rect 21591 22732 22008 22760
rect 21591 22729 21603 22732
rect 21545 22723 21603 22729
rect 22002 22720 22008 22732
rect 22060 22720 22066 22772
rect 22186 22720 22192 22772
rect 22244 22720 22250 22772
rect 22554 22760 22560 22772
rect 22296 22732 22560 22760
rect 19720 22692 19748 22720
rect 17420 22664 18552 22692
rect 16209 22655 16267 22661
rect 14415 22596 14596 22624
rect 14645 22627 14703 22633
rect 14415 22593 14427 22596
rect 14369 22587 14427 22593
rect 14645 22593 14657 22627
rect 14691 22593 14703 22627
rect 14645 22587 14703 22593
rect 14826 22584 14832 22636
rect 14884 22624 14890 22636
rect 16224 22624 16252 22655
rect 14884 22596 16252 22624
rect 14884 22584 14890 22596
rect 16482 22584 16488 22636
rect 16540 22584 16546 22636
rect 16666 22584 16672 22636
rect 16724 22624 16730 22636
rect 16853 22627 16911 22633
rect 16853 22624 16865 22627
rect 16724 22596 16865 22624
rect 16724 22584 16730 22596
rect 16853 22593 16865 22596
rect 16899 22624 16911 22627
rect 17402 22624 17408 22636
rect 16899 22596 17408 22624
rect 16899 22593 16911 22596
rect 16853 22587 16911 22593
rect 17402 22584 17408 22596
rect 17460 22584 17466 22636
rect 17589 22627 17647 22633
rect 17589 22593 17601 22627
rect 17635 22624 17647 22627
rect 18230 22624 18236 22636
rect 17635 22596 18236 22624
rect 17635 22593 17647 22596
rect 17589 22587 17647 22593
rect 18230 22584 18236 22596
rect 18288 22584 18294 22636
rect 10060 22528 10272 22556
rect 10244 22432 10272 22528
rect 10778 22516 10784 22568
rect 10836 22516 10842 22568
rect 11514 22516 11520 22568
rect 11572 22556 11578 22568
rect 13096 22556 13124 22584
rect 13449 22559 13507 22565
rect 13449 22556 13461 22559
rect 11572 22528 13461 22556
rect 11572 22516 11578 22528
rect 13449 22525 13461 22528
rect 13495 22525 13507 22559
rect 13449 22519 13507 22525
rect 13538 22516 13544 22568
rect 13596 22556 13602 22568
rect 14737 22559 14795 22565
rect 14737 22556 14749 22559
rect 13596 22528 14749 22556
rect 13596 22516 13602 22528
rect 14737 22525 14749 22528
rect 14783 22525 14795 22559
rect 16209 22559 16267 22565
rect 16209 22556 16221 22559
rect 14737 22519 14795 22525
rect 16132 22528 16221 22556
rect 13170 22448 13176 22500
rect 13228 22488 13234 22500
rect 14642 22488 14648 22500
rect 13228 22460 13676 22488
rect 13228 22448 13234 22460
rect 9858 22380 9864 22432
rect 9916 22380 9922 22432
rect 10226 22380 10232 22432
rect 10284 22380 10290 22432
rect 11146 22380 11152 22432
rect 11204 22380 11210 22432
rect 12434 22380 12440 22432
rect 12492 22420 12498 22432
rect 12529 22423 12587 22429
rect 12529 22420 12541 22423
rect 12492 22392 12541 22420
rect 12492 22380 12498 22392
rect 12529 22389 12541 22392
rect 12575 22389 12587 22423
rect 12529 22383 12587 22389
rect 13262 22380 13268 22432
rect 13320 22380 13326 22432
rect 13354 22380 13360 22432
rect 13412 22420 13418 22432
rect 13648 22429 13676 22460
rect 14016 22460 14648 22488
rect 14016 22429 14044 22460
rect 14642 22448 14648 22460
rect 14700 22448 14706 22500
rect 16132 22432 16160 22528
rect 16209 22525 16221 22528
rect 16255 22525 16267 22559
rect 16209 22519 16267 22525
rect 17126 22516 17132 22568
rect 17184 22516 17190 22568
rect 18524 22565 18552 22664
rect 19444 22664 19748 22692
rect 20824 22664 21680 22692
rect 19444 22633 19472 22664
rect 19429 22627 19487 22633
rect 19429 22593 19441 22627
rect 19475 22593 19487 22627
rect 19429 22587 19487 22593
rect 19610 22584 19616 22636
rect 19668 22584 19674 22636
rect 19705 22627 19763 22633
rect 19705 22593 19717 22627
rect 19751 22624 19763 22627
rect 19886 22624 19892 22636
rect 19751 22596 19892 22624
rect 19751 22593 19763 22596
rect 19705 22587 19763 22593
rect 19886 22584 19892 22596
rect 19944 22584 19950 22636
rect 19981 22627 20039 22633
rect 19981 22593 19993 22627
rect 20027 22624 20039 22627
rect 20254 22624 20260 22636
rect 20027 22596 20260 22624
rect 20027 22593 20039 22596
rect 19981 22587 20039 22593
rect 20254 22584 20260 22596
rect 20312 22624 20318 22636
rect 20441 22627 20499 22633
rect 20441 22624 20453 22627
rect 20312 22596 20453 22624
rect 20312 22584 20318 22596
rect 20441 22593 20453 22596
rect 20487 22593 20499 22627
rect 20441 22587 20499 22593
rect 20533 22627 20591 22633
rect 20533 22593 20545 22627
rect 20579 22593 20591 22627
rect 20533 22587 20591 22593
rect 17865 22559 17923 22565
rect 17865 22525 17877 22559
rect 17911 22525 17923 22559
rect 17865 22519 17923 22525
rect 18509 22559 18567 22565
rect 18509 22525 18521 22559
rect 18555 22525 18567 22559
rect 18509 22519 18567 22525
rect 19337 22559 19395 22565
rect 19337 22525 19349 22559
rect 19383 22525 19395 22559
rect 19337 22519 19395 22525
rect 19797 22559 19855 22565
rect 19797 22525 19809 22559
rect 19843 22556 19855 22559
rect 20162 22556 20168 22568
rect 19843 22528 20168 22556
rect 19843 22525 19855 22528
rect 19797 22519 19855 22525
rect 17880 22488 17908 22519
rect 19352 22488 19380 22519
rect 20162 22516 20168 22528
rect 20220 22516 20226 22568
rect 19426 22488 19432 22500
rect 17880 22460 18736 22488
rect 19352 22460 19432 22488
rect 13541 22423 13599 22429
rect 13541 22420 13553 22423
rect 13412 22392 13553 22420
rect 13412 22380 13418 22392
rect 13541 22389 13553 22392
rect 13587 22389 13599 22423
rect 13541 22383 13599 22389
rect 13633 22423 13691 22429
rect 13633 22389 13645 22423
rect 13679 22389 13691 22423
rect 13633 22383 13691 22389
rect 14001 22423 14059 22429
rect 14001 22389 14013 22423
rect 14047 22389 14059 22423
rect 14001 22383 14059 22389
rect 14274 22380 14280 22432
rect 14332 22380 14338 22432
rect 14553 22423 14611 22429
rect 14553 22389 14565 22423
rect 14599 22420 14611 22423
rect 15102 22420 15108 22432
rect 14599 22392 15108 22420
rect 14599 22389 14611 22392
rect 14553 22383 14611 22389
rect 15102 22380 15108 22392
rect 15160 22380 15166 22432
rect 16114 22380 16120 22432
rect 16172 22380 16178 22432
rect 16390 22380 16396 22432
rect 16448 22380 16454 22432
rect 17494 22380 17500 22432
rect 17552 22420 17558 22432
rect 17773 22423 17831 22429
rect 17773 22420 17785 22423
rect 17552 22392 17785 22420
rect 17552 22380 17558 22392
rect 17773 22389 17785 22392
rect 17819 22389 17831 22423
rect 17773 22383 17831 22389
rect 17954 22380 17960 22432
rect 18012 22380 18018 22432
rect 18708 22429 18736 22460
rect 19426 22448 19432 22460
rect 19484 22448 19490 22500
rect 18693 22423 18751 22429
rect 18693 22389 18705 22423
rect 18739 22420 18751 22423
rect 19610 22420 19616 22432
rect 18739 22392 19616 22420
rect 18739 22389 18751 22392
rect 18693 22383 18751 22389
rect 19610 22380 19616 22392
rect 19668 22380 19674 22432
rect 20165 22423 20223 22429
rect 20165 22389 20177 22423
rect 20211 22420 20223 22423
rect 20346 22420 20352 22432
rect 20211 22392 20352 22420
rect 20211 22389 20223 22392
rect 20165 22383 20223 22389
rect 20346 22380 20352 22392
rect 20404 22380 20410 22432
rect 20548 22420 20576 22587
rect 20824 22565 20852 22664
rect 21376 22636 21404 22664
rect 20901 22627 20959 22633
rect 20901 22593 20913 22627
rect 20947 22593 20959 22627
rect 20901 22587 20959 22593
rect 20809 22559 20867 22565
rect 20809 22525 20821 22559
rect 20855 22525 20867 22559
rect 20916 22556 20944 22587
rect 21358 22584 21364 22636
rect 21416 22584 21422 22636
rect 21453 22627 21511 22633
rect 21453 22593 21465 22627
rect 21499 22624 21511 22627
rect 21542 22624 21548 22636
rect 21499 22596 21548 22624
rect 21499 22593 21511 22596
rect 21453 22587 21511 22593
rect 21542 22584 21548 22596
rect 21600 22584 21606 22636
rect 21652 22633 21680 22664
rect 21637 22627 21695 22633
rect 21637 22593 21649 22627
rect 21683 22593 21695 22627
rect 21637 22587 21695 22593
rect 21726 22584 21732 22636
rect 21784 22624 21790 22636
rect 22204 22633 22232 22720
rect 22296 22633 22324 22732
rect 22554 22720 22560 22732
rect 22612 22720 22618 22772
rect 22741 22763 22799 22769
rect 22741 22729 22753 22763
rect 22787 22760 22799 22763
rect 22922 22760 22928 22772
rect 22787 22732 22928 22760
rect 22787 22729 22799 22732
rect 22741 22723 22799 22729
rect 22922 22720 22928 22732
rect 22980 22720 22986 22772
rect 23032 22732 23419 22760
rect 22462 22652 22468 22704
rect 22520 22692 22526 22704
rect 23032 22692 23060 22732
rect 22520 22664 23060 22692
rect 23100 22695 23158 22701
rect 22520 22652 22526 22664
rect 23100 22661 23112 22695
rect 23146 22692 23158 22695
rect 23290 22692 23296 22704
rect 23146 22664 23296 22692
rect 23146 22661 23158 22664
rect 23100 22655 23158 22661
rect 23290 22652 23296 22664
rect 23348 22652 23354 22704
rect 23391 22692 23419 22732
rect 24394 22720 24400 22772
rect 24452 22720 24458 22772
rect 23391 22664 24532 22692
rect 22005 22627 22063 22633
rect 22005 22624 22017 22627
rect 21784 22596 22017 22624
rect 21784 22584 21790 22596
rect 22005 22593 22017 22596
rect 22051 22593 22063 22627
rect 22005 22587 22063 22593
rect 22189 22627 22247 22633
rect 22189 22593 22201 22627
rect 22235 22593 22247 22627
rect 22189 22587 22247 22593
rect 22281 22627 22339 22633
rect 22281 22593 22293 22627
rect 22327 22593 22339 22627
rect 22281 22587 22339 22593
rect 22557 22627 22615 22633
rect 22557 22593 22569 22627
rect 22603 22624 22615 22627
rect 23566 22624 23572 22636
rect 22603 22596 23572 22624
rect 22603 22593 22615 22596
rect 22557 22587 22615 22593
rect 20916 22528 22324 22556
rect 20809 22519 20867 22525
rect 21269 22491 21327 22497
rect 21269 22457 21281 22491
rect 21315 22488 21327 22491
rect 22094 22488 22100 22500
rect 21315 22460 22100 22488
rect 21315 22457 21327 22460
rect 21269 22451 21327 22457
rect 22094 22448 22100 22460
rect 22152 22448 22158 22500
rect 22296 22488 22324 22528
rect 22370 22516 22376 22568
rect 22428 22516 22434 22568
rect 22664 22488 22692 22596
rect 23566 22584 23572 22596
rect 23624 22584 23630 22636
rect 24118 22584 24124 22636
rect 24176 22624 24182 22636
rect 24504 22633 24532 22664
rect 24305 22627 24363 22633
rect 24305 22624 24317 22627
rect 24176 22596 24317 22624
rect 24176 22584 24182 22596
rect 24305 22593 24317 22596
rect 24351 22593 24363 22627
rect 24305 22587 24363 22593
rect 24489 22627 24547 22633
rect 24489 22593 24501 22627
rect 24535 22593 24547 22627
rect 24489 22587 24547 22593
rect 22830 22516 22836 22568
rect 22888 22516 22894 22568
rect 22296 22460 22692 22488
rect 24210 22420 24216 22432
rect 20548 22392 24216 22420
rect 24210 22380 24216 22392
rect 24268 22380 24274 22432
rect 1104 22330 34868 22352
rect 1104 22278 5170 22330
rect 5222 22278 5234 22330
rect 5286 22278 5298 22330
rect 5350 22278 5362 22330
rect 5414 22278 5426 22330
rect 5478 22278 13611 22330
rect 13663 22278 13675 22330
rect 13727 22278 13739 22330
rect 13791 22278 13803 22330
rect 13855 22278 13867 22330
rect 13919 22278 22052 22330
rect 22104 22278 22116 22330
rect 22168 22278 22180 22330
rect 22232 22278 22244 22330
rect 22296 22278 22308 22330
rect 22360 22278 30493 22330
rect 30545 22278 30557 22330
rect 30609 22278 30621 22330
rect 30673 22278 30685 22330
rect 30737 22278 30749 22330
rect 30801 22278 34868 22330
rect 1104 22256 34868 22278
rect 13078 22176 13084 22228
rect 13136 22216 13142 22228
rect 16114 22216 16120 22228
rect 13136 22188 16120 22216
rect 13136 22176 13142 22188
rect 16114 22176 16120 22188
rect 16172 22176 16178 22228
rect 19429 22219 19487 22225
rect 19429 22216 19441 22219
rect 18984 22188 19441 22216
rect 10321 22151 10379 22157
rect 10321 22117 10333 22151
rect 10367 22148 10379 22151
rect 10778 22148 10784 22160
rect 10367 22120 10784 22148
rect 10367 22117 10379 22120
rect 10321 22111 10379 22117
rect 8938 22040 8944 22092
rect 8996 22040 9002 22092
rect 10428 22089 10456 22120
rect 10778 22108 10784 22120
rect 10836 22108 10842 22160
rect 12434 22108 12440 22160
rect 12492 22108 12498 22160
rect 13909 22151 13967 22157
rect 13909 22117 13921 22151
rect 13955 22148 13967 22151
rect 14366 22148 14372 22160
rect 13955 22120 14372 22148
rect 13955 22117 13967 22120
rect 13909 22111 13967 22117
rect 14366 22108 14372 22120
rect 14424 22108 14430 22160
rect 15286 22148 15292 22160
rect 14568 22120 14964 22148
rect 10413 22083 10471 22089
rect 10413 22049 10425 22083
rect 10459 22049 10471 22083
rect 10413 22043 10471 22049
rect 10796 22052 11192 22080
rect 10796 22021 10824 22052
rect 11164 22024 11192 22052
rect 11974 22040 11980 22092
rect 12032 22080 12038 22092
rect 12345 22083 12403 22089
rect 12032 22052 12296 22080
rect 12032 22040 12038 22052
rect 2685 22015 2743 22021
rect 2685 21981 2697 22015
rect 2731 22012 2743 22015
rect 10781 22015 10839 22021
rect 2731 21984 9444 22012
rect 2731 21981 2743 21984
rect 2685 21975 2743 21981
rect 934 21904 940 21956
rect 992 21944 998 21956
rect 1581 21947 1639 21953
rect 1581 21944 1593 21947
rect 992 21916 1593 21944
rect 992 21904 998 21916
rect 1581 21913 1593 21916
rect 1627 21913 1639 21947
rect 1581 21907 1639 21913
rect 9208 21947 9266 21953
rect 9208 21913 9220 21947
rect 9254 21944 9266 21947
rect 9306 21944 9312 21956
rect 9254 21916 9312 21944
rect 9254 21913 9266 21916
rect 9208 21907 9266 21913
rect 9306 21904 9312 21916
rect 9364 21904 9370 21956
rect 9416 21944 9444 21984
rect 10781 21981 10793 22015
rect 10827 21981 10839 22015
rect 10781 21975 10839 21981
rect 10962 21972 10968 22024
rect 11020 21972 11026 22024
rect 11146 21972 11152 22024
rect 11204 21972 11210 22024
rect 11238 21972 11244 22024
rect 11296 21972 11302 22024
rect 11514 21972 11520 22024
rect 11572 21972 11578 22024
rect 11609 22015 11667 22021
rect 11609 21981 11621 22015
rect 11655 22012 11667 22015
rect 12066 22012 12072 22024
rect 11655 21984 12072 22012
rect 11655 21981 11667 21984
rect 11609 21975 11667 21981
rect 12066 21972 12072 21984
rect 12124 21972 12130 22024
rect 12268 22021 12296 22052
rect 12345 22049 12357 22083
rect 12391 22080 12403 22083
rect 12452 22080 12480 22108
rect 13262 22080 13268 22092
rect 12391 22052 12480 22080
rect 13188 22052 13268 22080
rect 12391 22049 12403 22052
rect 12345 22043 12403 22049
rect 12253 22015 12311 22021
rect 12253 21981 12265 22015
rect 12299 21981 12311 22015
rect 12253 21975 12311 21981
rect 12437 22015 12495 22021
rect 12437 21981 12449 22015
rect 12483 21981 12495 22015
rect 12437 21975 12495 21981
rect 10873 21947 10931 21953
rect 10873 21944 10885 21947
rect 9416 21916 10885 21944
rect 10873 21913 10885 21916
rect 10919 21913 10931 21947
rect 11256 21944 11284 21972
rect 12452 21944 12480 21975
rect 12618 21972 12624 22024
rect 12676 21972 12682 22024
rect 13188 22021 13216 22052
rect 13262 22040 13268 22052
rect 13320 22080 13326 22092
rect 14568 22080 14596 22120
rect 14936 22089 14964 22120
rect 15120 22120 15292 22148
rect 13320 22052 14412 22080
rect 13320 22040 13326 22052
rect 13173 22015 13231 22021
rect 13173 21981 13185 22015
rect 13219 21981 13231 22015
rect 13173 21975 13231 21981
rect 13633 22015 13691 22021
rect 13633 21981 13645 22015
rect 13679 22012 13691 22015
rect 13814 22012 13820 22024
rect 13679 21984 13820 22012
rect 13679 21981 13691 21984
rect 13633 21975 13691 21981
rect 13814 21972 13820 21984
rect 13872 21972 13878 22024
rect 13909 22015 13967 22021
rect 13909 21981 13921 22015
rect 13955 21981 13967 22015
rect 13909 21975 13967 21981
rect 13357 21947 13415 21953
rect 11256 21916 12388 21944
rect 12452 21916 12756 21944
rect 10873 21907 10931 21913
rect 12360 21888 12388 21916
rect 12728 21888 12756 21916
rect 13357 21913 13369 21947
rect 13403 21944 13415 21947
rect 13924 21944 13952 21975
rect 14182 21972 14188 22024
rect 14240 22021 14246 22024
rect 14384 22021 14412 22052
rect 14476 22052 14596 22080
rect 14921 22083 14979 22089
rect 14476 22021 14504 22052
rect 14921 22049 14933 22083
rect 14967 22080 14979 22083
rect 15120 22080 15148 22120
rect 15286 22108 15292 22120
rect 15344 22108 15350 22160
rect 15565 22151 15623 22157
rect 15565 22117 15577 22151
rect 15611 22148 15623 22151
rect 15611 22120 16574 22148
rect 15611 22117 15623 22120
rect 15565 22111 15623 22117
rect 16117 22083 16175 22089
rect 16117 22080 16129 22083
rect 14967 22052 15148 22080
rect 15212 22052 16129 22080
rect 14967 22049 14979 22052
rect 14921 22043 14979 22049
rect 15212 22024 15240 22052
rect 16117 22049 16129 22052
rect 16163 22049 16175 22083
rect 16546 22080 16574 22120
rect 16945 22083 17003 22089
rect 16945 22080 16957 22083
rect 16546 22052 16957 22080
rect 16117 22043 16175 22049
rect 16945 22049 16957 22052
rect 16991 22049 17003 22083
rect 16945 22043 17003 22049
rect 14240 22015 14289 22021
rect 14240 21981 14243 22015
rect 14277 21981 14289 22015
rect 14240 21975 14289 21981
rect 14369 22015 14427 22021
rect 14369 21981 14381 22015
rect 14415 21981 14427 22015
rect 14369 21975 14427 21981
rect 14461 22015 14519 22021
rect 14461 21981 14473 22015
rect 14507 21981 14519 22015
rect 14642 22012 14648 22024
rect 14603 21984 14648 22012
rect 14461 21975 14519 21981
rect 14240 21972 14246 21975
rect 14642 21972 14648 21984
rect 14700 21972 14706 22024
rect 14734 21972 14740 22024
rect 14792 21972 14798 22024
rect 14829 22015 14887 22021
rect 14829 21981 14841 22015
rect 14875 21981 14887 22015
rect 14829 21975 14887 21981
rect 14660 21944 14688 21972
rect 14844 21944 14872 21975
rect 15102 21972 15108 22024
rect 15160 21972 15166 22024
rect 15194 21972 15200 22024
rect 15252 21972 15258 22024
rect 15749 22015 15807 22021
rect 15749 21981 15761 22015
rect 15795 22012 15807 22015
rect 15838 22012 15844 22024
rect 15795 21984 15844 22012
rect 15795 21981 15807 21984
rect 15749 21975 15807 21981
rect 15838 21972 15844 21984
rect 15896 21972 15902 22024
rect 15933 22015 15991 22021
rect 15933 21981 15945 22015
rect 15979 21981 15991 22015
rect 15933 21975 15991 21981
rect 16025 22015 16083 22021
rect 16025 21981 16037 22015
rect 16071 22012 16083 22015
rect 17402 22012 17408 22024
rect 16071 21984 17408 22012
rect 16071 21981 16083 21984
rect 16025 21975 16083 21981
rect 13403 21916 13860 21944
rect 13924 21916 14596 21944
rect 14660 21916 14872 21944
rect 13403 21913 13415 21916
rect 13357 21907 13415 21913
rect 11882 21836 11888 21888
rect 11940 21836 11946 21888
rect 12342 21836 12348 21888
rect 12400 21836 12406 21888
rect 12710 21836 12716 21888
rect 12768 21836 12774 21888
rect 12986 21836 12992 21888
rect 13044 21836 13050 21888
rect 13722 21836 13728 21888
rect 13780 21836 13786 21888
rect 13832 21876 13860 21916
rect 13998 21876 14004 21888
rect 13832 21848 14004 21876
rect 13998 21836 14004 21848
rect 14056 21836 14062 21888
rect 14090 21836 14096 21888
rect 14148 21836 14154 21888
rect 14568 21876 14596 21916
rect 14826 21876 14832 21888
rect 14568 21848 14832 21876
rect 14826 21836 14832 21848
rect 14884 21836 14890 21888
rect 15378 21836 15384 21888
rect 15436 21836 15442 21888
rect 15948 21876 15976 21975
rect 17402 21972 17408 21984
rect 17460 21972 17466 22024
rect 17678 21972 17684 22024
rect 17736 21972 17742 22024
rect 17954 22021 17960 22024
rect 17948 21975 17960 22021
rect 17954 21972 17960 21975
rect 18012 21972 18018 22024
rect 18414 21972 18420 22024
rect 18472 22012 18478 22024
rect 18984 22012 19012 22188
rect 19429 22185 19441 22188
rect 19475 22185 19487 22219
rect 19429 22179 19487 22185
rect 20806 22176 20812 22228
rect 20864 22176 20870 22228
rect 21358 22176 21364 22228
rect 21416 22176 21422 22228
rect 21910 22176 21916 22228
rect 21968 22216 21974 22228
rect 23385 22219 23443 22225
rect 23385 22216 23397 22219
rect 21968 22188 23397 22216
rect 21968 22176 21974 22188
rect 23385 22185 23397 22188
rect 23431 22185 23443 22219
rect 23385 22179 23443 22185
rect 23477 22219 23535 22225
rect 23477 22185 23489 22219
rect 23523 22216 23535 22219
rect 23658 22216 23664 22228
rect 23523 22188 23664 22216
rect 23523 22185 23535 22188
rect 23477 22179 23535 22185
rect 19061 22151 19119 22157
rect 19061 22117 19073 22151
rect 19107 22117 19119 22151
rect 19061 22111 19119 22117
rect 18472 21984 19012 22012
rect 19076 22012 19104 22111
rect 20070 22040 20076 22092
rect 20128 22040 20134 22092
rect 21376 22080 21404 22176
rect 21542 22108 21548 22160
rect 21600 22148 21606 22160
rect 23492 22148 23520 22179
rect 23658 22176 23664 22188
rect 23716 22176 23722 22228
rect 21600 22120 23520 22148
rect 21600 22108 21606 22120
rect 21910 22080 21916 22092
rect 21376 22052 21916 22080
rect 21910 22040 21916 22052
rect 21968 22080 21974 22092
rect 23293 22083 23351 22089
rect 23293 22080 23305 22083
rect 21968 22052 23305 22080
rect 21968 22040 21974 22052
rect 23293 22049 23305 22052
rect 23339 22049 23351 22083
rect 23293 22043 23351 22049
rect 24302 22040 24308 22092
rect 24360 22040 24366 22092
rect 19426 22012 19432 22024
rect 19076 21984 19432 22012
rect 18472 21972 18478 21984
rect 19426 21972 19432 21984
rect 19484 22012 19490 22024
rect 19884 22015 19942 22021
rect 19884 22012 19896 22015
rect 19484 21984 19896 22012
rect 19484 21972 19490 21984
rect 19884 21981 19896 21984
rect 19930 22012 19942 22015
rect 20088 22012 20116 22040
rect 19930 21984 20116 22012
rect 19930 21981 19942 21984
rect 19884 21975 19942 21981
rect 20162 21972 20168 22024
rect 20220 21972 20226 22024
rect 20254 21972 20260 22024
rect 20312 21972 20318 22024
rect 20346 21972 20352 22024
rect 20404 21972 20410 22024
rect 20717 22015 20775 22021
rect 20717 21981 20729 22015
rect 20763 22012 20775 22015
rect 20898 22012 20904 22024
rect 20763 21984 20904 22012
rect 20763 21981 20775 21984
rect 20717 21975 20775 21981
rect 16684 21916 19380 21944
rect 16684 21876 16712 21916
rect 15948 21848 16712 21876
rect 16758 21836 16764 21888
rect 16816 21836 16822 21888
rect 17310 21836 17316 21888
rect 17368 21876 17374 21888
rect 17589 21879 17647 21885
rect 17589 21876 17601 21879
rect 17368 21848 17601 21876
rect 17368 21836 17374 21848
rect 17589 21845 17601 21848
rect 17635 21845 17647 21879
rect 17589 21839 17647 21845
rect 18782 21836 18788 21888
rect 18840 21876 18846 21888
rect 19242 21876 19248 21888
rect 18840 21848 19248 21876
rect 18840 21836 18846 21848
rect 19242 21836 19248 21848
rect 19300 21836 19306 21888
rect 19352 21876 19380 21916
rect 19610 21904 19616 21956
rect 19668 21904 19674 21956
rect 19981 21947 20039 21953
rect 19981 21913 19993 21947
rect 20027 21913 20039 21947
rect 19981 21907 20039 21913
rect 20073 21947 20131 21953
rect 20073 21913 20085 21947
rect 20119 21944 20131 21947
rect 20180 21944 20208 21972
rect 20119 21916 20208 21944
rect 20119 21913 20131 21916
rect 20073 21907 20131 21913
rect 19426 21885 19432 21888
rect 19408 21879 19432 21885
rect 19408 21876 19420 21879
rect 19352 21848 19420 21876
rect 19408 21845 19420 21848
rect 19408 21839 19432 21845
rect 19426 21836 19432 21839
rect 19484 21836 19490 21888
rect 19705 21879 19763 21885
rect 19705 21845 19717 21879
rect 19751 21876 19763 21879
rect 19886 21876 19892 21888
rect 19751 21848 19892 21876
rect 19751 21845 19763 21848
rect 19705 21839 19763 21845
rect 19886 21836 19892 21848
rect 19944 21836 19950 21888
rect 19996 21876 20024 21907
rect 20732 21876 20760 21975
rect 20898 21972 20904 21984
rect 20956 21972 20962 22024
rect 20990 21972 20996 22024
rect 21048 21972 21054 22024
rect 21085 22015 21143 22021
rect 21085 21981 21097 22015
rect 21131 22012 21143 22015
rect 22462 22012 22468 22024
rect 21131 21984 22468 22012
rect 21131 21981 21143 21984
rect 21085 21975 21143 21981
rect 22462 21972 22468 21984
rect 22520 21972 22526 22024
rect 23566 21972 23572 22024
rect 23624 22012 23630 22024
rect 24320 22012 24348 22040
rect 23624 21984 24348 22012
rect 23624 21972 23630 21984
rect 19996 21848 20760 21876
rect 21266 21836 21272 21888
rect 21324 21836 21330 21888
rect 1104 21786 35027 21808
rect 1104 21734 9390 21786
rect 9442 21734 9454 21786
rect 9506 21734 9518 21786
rect 9570 21734 9582 21786
rect 9634 21734 9646 21786
rect 9698 21734 17831 21786
rect 17883 21734 17895 21786
rect 17947 21734 17959 21786
rect 18011 21734 18023 21786
rect 18075 21734 18087 21786
rect 18139 21734 26272 21786
rect 26324 21734 26336 21786
rect 26388 21734 26400 21786
rect 26452 21734 26464 21786
rect 26516 21734 26528 21786
rect 26580 21734 34713 21786
rect 34765 21734 34777 21786
rect 34829 21734 34841 21786
rect 34893 21734 34905 21786
rect 34957 21734 34969 21786
rect 35021 21734 35027 21786
rect 1104 21712 35027 21734
rect 9306 21632 9312 21684
rect 9364 21672 9370 21684
rect 9493 21675 9551 21681
rect 9493 21672 9505 21675
rect 9364 21644 9505 21672
rect 9364 21632 9370 21644
rect 9493 21641 9505 21644
rect 9539 21641 9551 21675
rect 9493 21635 9551 21641
rect 10413 21675 10471 21681
rect 10413 21641 10425 21675
rect 10459 21672 10471 21675
rect 10962 21672 10968 21684
rect 10459 21644 10968 21672
rect 10459 21641 10471 21644
rect 10413 21635 10471 21641
rect 10962 21632 10968 21644
rect 11020 21632 11026 21684
rect 11146 21632 11152 21684
rect 11204 21632 11210 21684
rect 11517 21675 11575 21681
rect 11517 21641 11529 21675
rect 11563 21641 11575 21675
rect 11517 21635 11575 21641
rect 10226 21604 10232 21616
rect 8956 21576 10232 21604
rect 8956 21545 8984 21576
rect 10226 21564 10232 21576
rect 10284 21564 10290 21616
rect 11164 21604 11192 21632
rect 10612 21576 11192 21604
rect 8941 21539 8999 21545
rect 8941 21505 8953 21539
rect 8987 21505 8999 21539
rect 8941 21499 8999 21505
rect 9217 21539 9275 21545
rect 9217 21505 9229 21539
rect 9263 21536 9275 21539
rect 9858 21536 9864 21548
rect 9263 21508 9864 21536
rect 9263 21505 9275 21508
rect 9217 21499 9275 21505
rect 9858 21496 9864 21508
rect 9916 21496 9922 21548
rect 10612 21545 10640 21576
rect 10597 21539 10655 21545
rect 10597 21505 10609 21539
rect 10643 21505 10655 21539
rect 10597 21499 10655 21505
rect 10686 21496 10692 21548
rect 10744 21496 10750 21548
rect 10778 21496 10784 21548
rect 10836 21496 10842 21548
rect 10962 21496 10968 21548
rect 11020 21536 11026 21548
rect 11149 21539 11207 21545
rect 11020 21508 11100 21536
rect 11020 21496 11026 21508
rect 9401 21471 9459 21477
rect 9401 21437 9413 21471
rect 9447 21468 9459 21471
rect 10045 21471 10103 21477
rect 10045 21468 10057 21471
rect 9447 21440 10057 21468
rect 9447 21437 9459 21440
rect 9401 21431 9459 21437
rect 10045 21437 10057 21440
rect 10091 21437 10103 21471
rect 10704 21468 10732 21496
rect 10873 21471 10931 21477
rect 10873 21468 10885 21471
rect 10704 21440 10885 21468
rect 10045 21431 10103 21437
rect 10873 21437 10885 21440
rect 10919 21437 10931 21471
rect 11072 21468 11100 21508
rect 11149 21505 11161 21539
rect 11195 21536 11207 21539
rect 11532 21536 11560 21635
rect 11882 21632 11888 21684
rect 11940 21632 11946 21684
rect 12437 21675 12495 21681
rect 12437 21641 12449 21675
rect 12483 21672 12495 21675
rect 12618 21672 12624 21684
rect 12483 21644 12624 21672
rect 12483 21641 12495 21644
rect 12437 21635 12495 21641
rect 12618 21632 12624 21644
rect 12676 21632 12682 21684
rect 12986 21632 12992 21684
rect 13044 21632 13050 21684
rect 13188 21644 13676 21672
rect 11900 21604 11928 21632
rect 12713 21607 12771 21613
rect 12713 21604 12725 21607
rect 11900 21576 12204 21604
rect 11195 21508 11560 21536
rect 11696 21539 11754 21545
rect 11195 21505 11207 21508
rect 11149 21499 11207 21505
rect 11696 21505 11708 21539
rect 11742 21505 11754 21539
rect 11696 21499 11754 21505
rect 11793 21539 11851 21545
rect 11793 21505 11805 21539
rect 11839 21505 11851 21539
rect 11793 21499 11851 21505
rect 11716 21468 11744 21499
rect 11072 21440 11744 21468
rect 10873 21431 10931 21437
rect 10888 21400 10916 21431
rect 11808 21400 11836 21499
rect 11882 21496 11888 21548
rect 11940 21496 11946 21548
rect 12066 21536 12072 21548
rect 12027 21508 12072 21536
rect 12066 21496 12072 21508
rect 12124 21496 12130 21548
rect 12176 21545 12204 21576
rect 12544 21576 12725 21604
rect 12161 21539 12219 21545
rect 12161 21505 12173 21539
rect 12207 21505 12219 21539
rect 12161 21499 12219 21505
rect 12434 21496 12440 21548
rect 12492 21536 12498 21548
rect 12544 21536 12572 21576
rect 12713 21573 12725 21576
rect 12759 21573 12771 21607
rect 12713 21567 12771 21573
rect 12805 21607 12863 21613
rect 12805 21573 12817 21607
rect 12851 21604 12863 21607
rect 13004 21604 13032 21632
rect 12851 21576 13032 21604
rect 12851 21573 12863 21576
rect 12805 21567 12863 21573
rect 12492 21508 12572 21536
rect 12492 21496 12498 21508
rect 12618 21496 12624 21548
rect 12676 21496 12682 21548
rect 12989 21539 13047 21545
rect 12989 21505 13001 21539
rect 13035 21536 13047 21539
rect 13188 21536 13216 21644
rect 13648 21604 13676 21644
rect 13722 21632 13728 21684
rect 13780 21672 13786 21684
rect 13780 21644 14228 21672
rect 13780 21632 13786 21644
rect 14090 21604 14096 21616
rect 13648 21576 14096 21604
rect 14090 21564 14096 21576
rect 14148 21564 14154 21616
rect 14200 21604 14228 21644
rect 15102 21632 15108 21684
rect 15160 21632 15166 21684
rect 15470 21632 15476 21684
rect 15528 21672 15534 21684
rect 16482 21672 16488 21684
rect 15528 21644 16488 21672
rect 15528 21632 15534 21644
rect 16482 21632 16488 21644
rect 16540 21672 16546 21684
rect 16669 21675 16727 21681
rect 16669 21672 16681 21675
rect 16540 21644 16681 21672
rect 16540 21632 16546 21644
rect 16669 21641 16681 21644
rect 16715 21641 16727 21675
rect 16669 21635 16727 21641
rect 16758 21632 16764 21684
rect 16816 21632 16822 21684
rect 17310 21632 17316 21684
rect 17368 21632 17374 21684
rect 17402 21632 17408 21684
rect 17460 21672 17466 21684
rect 18414 21672 18420 21684
rect 17460 21644 18420 21672
rect 17460 21632 17466 21644
rect 18414 21632 18420 21644
rect 18472 21632 18478 21684
rect 19426 21672 19432 21684
rect 19352 21644 19432 21672
rect 15488 21604 15516 21632
rect 14200 21576 15516 21604
rect 13035 21508 13216 21536
rect 13035 21505 13047 21508
rect 12989 21499 13047 21505
rect 13262 21496 13268 21548
rect 13320 21496 13326 21548
rect 13538 21496 13544 21548
rect 13596 21545 13602 21548
rect 13596 21499 13605 21545
rect 13725 21539 13783 21545
rect 13725 21505 13737 21539
rect 13771 21536 13783 21539
rect 13771 21508 14872 21536
rect 13771 21505 13783 21508
rect 13725 21499 13783 21505
rect 13596 21496 13602 21499
rect 13446 21428 13452 21480
rect 13504 21468 13510 21480
rect 13817 21471 13875 21477
rect 13817 21468 13829 21471
rect 13504 21440 13829 21468
rect 13504 21428 13510 21440
rect 13817 21437 13829 21440
rect 13863 21437 13875 21471
rect 13817 21431 13875 21437
rect 13924 21400 13952 21508
rect 14182 21428 14188 21480
rect 14240 21468 14246 21480
rect 14369 21471 14427 21477
rect 14369 21468 14381 21471
rect 14240 21440 14381 21468
rect 14240 21428 14246 21440
rect 14369 21437 14381 21440
rect 14415 21437 14427 21471
rect 14844 21468 14872 21508
rect 14918 21496 14924 21548
rect 14976 21496 14982 21548
rect 15010 21496 15016 21548
rect 15068 21496 15074 21548
rect 15194 21496 15200 21548
rect 15252 21496 15258 21548
rect 15381 21539 15439 21545
rect 15381 21505 15393 21539
rect 15427 21536 15439 21539
rect 16666 21536 16672 21548
rect 15427 21508 16672 21536
rect 15427 21505 15439 21508
rect 15381 21499 15439 21505
rect 16666 21496 16672 21508
rect 16724 21496 16730 21548
rect 16776 21536 16804 21632
rect 17212 21607 17270 21613
rect 17212 21573 17224 21607
rect 17258 21604 17270 21607
rect 17328 21604 17356 21632
rect 17258 21576 17356 21604
rect 17258 21573 17270 21576
rect 17212 21567 17270 21573
rect 16853 21539 16911 21545
rect 16853 21536 16865 21539
rect 16776 21508 16865 21536
rect 16853 21505 16865 21508
rect 16899 21505 16911 21539
rect 16853 21499 16911 21505
rect 17494 21496 17500 21548
rect 17552 21536 17558 21548
rect 19352 21545 19380 21644
rect 19426 21632 19432 21644
rect 19484 21632 19490 21684
rect 20162 21632 20168 21684
rect 20220 21632 20226 21684
rect 20806 21632 20812 21684
rect 20864 21672 20870 21684
rect 21818 21672 21824 21684
rect 20864 21644 21824 21672
rect 20864 21632 20870 21644
rect 21818 21632 21824 21644
rect 21876 21632 21882 21684
rect 22462 21632 22468 21684
rect 22520 21672 22526 21684
rect 22557 21675 22615 21681
rect 22557 21672 22569 21675
rect 22520 21644 22569 21672
rect 22520 21632 22526 21644
rect 22557 21641 22569 21644
rect 22603 21641 22615 21675
rect 22557 21635 22615 21641
rect 20180 21604 20208 21632
rect 19444 21576 20208 21604
rect 19153 21539 19211 21545
rect 19153 21536 19165 21539
rect 17552 21508 19165 21536
rect 17552 21496 17558 21508
rect 19153 21505 19165 21508
rect 19199 21505 19211 21539
rect 19153 21499 19211 21505
rect 19337 21539 19395 21545
rect 19337 21505 19349 21539
rect 19383 21505 19395 21539
rect 19337 21499 19395 21505
rect 15028 21468 15056 21496
rect 14844 21440 15056 21468
rect 15212 21468 15240 21496
rect 15654 21468 15660 21480
rect 15212 21440 15660 21468
rect 14369 21431 14427 21437
rect 15654 21428 15660 21440
rect 15712 21428 15718 21480
rect 15933 21471 15991 21477
rect 15933 21437 15945 21471
rect 15979 21437 15991 21471
rect 15933 21431 15991 21437
rect 10888 21372 11836 21400
rect 12406 21372 13952 21400
rect 9030 21292 9036 21344
rect 9088 21332 9094 21344
rect 9214 21332 9220 21344
rect 9088 21304 9220 21332
rect 9088 21292 9094 21304
rect 9214 21292 9220 21304
rect 9272 21292 9278 21344
rect 9950 21292 9956 21344
rect 10008 21332 10014 21344
rect 12406 21332 12434 21372
rect 14458 21360 14464 21412
rect 14516 21400 14522 21412
rect 15948 21400 15976 21431
rect 16942 21428 16948 21480
rect 17000 21428 17006 21480
rect 19061 21471 19119 21477
rect 19061 21468 19073 21471
rect 18340 21440 19073 21468
rect 18340 21409 18368 21440
rect 19061 21437 19073 21440
rect 19107 21468 19119 21471
rect 19444 21468 19472 21576
rect 21082 21564 21088 21616
rect 21140 21604 21146 21616
rect 21542 21604 21548 21616
rect 21140 21576 21548 21604
rect 21140 21564 21146 21576
rect 21542 21564 21548 21576
rect 21600 21604 21606 21616
rect 21600 21576 22508 21604
rect 21600 21564 21606 21576
rect 19886 21496 19892 21548
rect 19944 21496 19950 21548
rect 20070 21496 20076 21548
rect 20128 21496 20134 21548
rect 20441 21539 20499 21545
rect 20441 21505 20453 21539
rect 20487 21505 20499 21539
rect 20441 21499 20499 21505
rect 19107 21440 19472 21468
rect 19521 21471 19579 21477
rect 19107 21437 19119 21440
rect 19061 21431 19119 21437
rect 19521 21437 19533 21471
rect 19567 21437 19579 21471
rect 19521 21431 19579 21437
rect 20165 21471 20223 21477
rect 20165 21437 20177 21471
rect 20211 21437 20223 21471
rect 20165 21431 20223 21437
rect 20257 21471 20315 21477
rect 20257 21437 20269 21471
rect 20303 21468 20315 21471
rect 20346 21468 20352 21480
rect 20303 21440 20352 21468
rect 20303 21437 20315 21440
rect 20257 21431 20315 21437
rect 14516 21372 15976 21400
rect 18325 21403 18383 21409
rect 14516 21360 14522 21372
rect 18325 21369 18337 21403
rect 18371 21369 18383 21403
rect 18325 21363 18383 21369
rect 18414 21360 18420 21412
rect 18472 21400 18478 21412
rect 19536 21400 19564 21431
rect 18472 21372 19564 21400
rect 20180 21400 20208 21431
rect 20346 21428 20352 21440
rect 20404 21428 20410 21480
rect 20456 21468 20484 21499
rect 21266 21496 21272 21548
rect 21324 21536 21330 21548
rect 21361 21539 21419 21545
rect 21361 21536 21373 21539
rect 21324 21508 21373 21536
rect 21324 21496 21330 21508
rect 21361 21505 21373 21508
rect 21407 21505 21419 21539
rect 21361 21499 21419 21505
rect 21818 21496 21824 21548
rect 21876 21496 21882 21548
rect 22480 21545 22508 21576
rect 22373 21539 22431 21545
rect 22373 21505 22385 21539
rect 22419 21505 22431 21539
rect 22373 21499 22431 21505
rect 22465 21539 22523 21545
rect 22465 21505 22477 21539
rect 22511 21505 22523 21539
rect 22465 21499 22523 21505
rect 20714 21468 20720 21480
rect 20456 21440 20720 21468
rect 20714 21428 20720 21440
rect 20772 21468 20778 21480
rect 22281 21471 22339 21477
rect 22281 21468 22293 21471
rect 20772 21440 22293 21468
rect 20772 21428 20778 21440
rect 22281 21437 22293 21440
rect 22327 21437 22339 21471
rect 22388 21468 22416 21499
rect 22646 21496 22652 21548
rect 22704 21496 22710 21548
rect 23474 21468 23480 21480
rect 22388 21440 23480 21468
rect 22281 21431 22339 21437
rect 23474 21428 23480 21440
rect 23532 21428 23538 21480
rect 20180 21372 20944 21400
rect 18472 21360 18478 21372
rect 20916 21344 20944 21372
rect 10008 21304 12434 21332
rect 10008 21292 10014 21304
rect 13078 21292 13084 21344
rect 13136 21292 13142 21344
rect 13170 21292 13176 21344
rect 13228 21332 13234 21344
rect 13541 21335 13599 21341
rect 13541 21332 13553 21335
rect 13228 21304 13553 21332
rect 13228 21292 13234 21304
rect 13541 21301 13553 21304
rect 13587 21301 13599 21335
rect 13541 21295 13599 21301
rect 14734 21292 14740 21344
rect 14792 21292 14798 21344
rect 15102 21292 15108 21344
rect 15160 21332 15166 21344
rect 15657 21335 15715 21341
rect 15657 21332 15669 21335
rect 15160 21304 15669 21332
rect 15160 21292 15166 21304
rect 15657 21301 15669 21304
rect 15703 21332 15715 21335
rect 15746 21332 15752 21344
rect 15703 21304 15752 21332
rect 15703 21301 15715 21304
rect 15657 21295 15715 21301
rect 15746 21292 15752 21304
rect 15804 21292 15810 21344
rect 16482 21292 16488 21344
rect 16540 21292 16546 21344
rect 20622 21292 20628 21344
rect 20680 21292 20686 21344
rect 20806 21292 20812 21344
rect 20864 21292 20870 21344
rect 20898 21292 20904 21344
rect 20956 21292 20962 21344
rect 21726 21292 21732 21344
rect 21784 21332 21790 21344
rect 22005 21335 22063 21341
rect 22005 21332 22017 21335
rect 21784 21304 22017 21332
rect 21784 21292 21790 21304
rect 22005 21301 22017 21304
rect 22051 21332 22063 21335
rect 22370 21332 22376 21344
rect 22051 21304 22376 21332
rect 22051 21301 22063 21304
rect 22005 21295 22063 21301
rect 22370 21292 22376 21304
rect 22428 21292 22434 21344
rect 22554 21292 22560 21344
rect 22612 21332 22618 21344
rect 22925 21335 22983 21341
rect 22925 21332 22937 21335
rect 22612 21304 22937 21332
rect 22612 21292 22618 21304
rect 22925 21301 22937 21304
rect 22971 21301 22983 21335
rect 22925 21295 22983 21301
rect 1104 21242 34868 21264
rect 1104 21190 5170 21242
rect 5222 21190 5234 21242
rect 5286 21190 5298 21242
rect 5350 21190 5362 21242
rect 5414 21190 5426 21242
rect 5478 21190 13611 21242
rect 13663 21190 13675 21242
rect 13727 21190 13739 21242
rect 13791 21190 13803 21242
rect 13855 21190 13867 21242
rect 13919 21190 22052 21242
rect 22104 21190 22116 21242
rect 22168 21190 22180 21242
rect 22232 21190 22244 21242
rect 22296 21190 22308 21242
rect 22360 21190 30493 21242
rect 30545 21190 30557 21242
rect 30609 21190 30621 21242
rect 30673 21190 30685 21242
rect 30737 21190 30749 21242
rect 30801 21190 34868 21242
rect 1104 21168 34868 21190
rect 8665 21131 8723 21137
rect 8665 21097 8677 21131
rect 8711 21128 8723 21131
rect 9766 21128 9772 21140
rect 8711 21100 9772 21128
rect 8711 21097 8723 21100
rect 8665 21091 8723 21097
rect 9766 21088 9772 21100
rect 9824 21088 9830 21140
rect 12621 21131 12679 21137
rect 12621 21097 12633 21131
rect 12667 21128 12679 21131
rect 13078 21128 13084 21140
rect 12667 21100 13084 21128
rect 12667 21097 12679 21100
rect 12621 21091 12679 21097
rect 13078 21088 13084 21100
rect 13136 21088 13142 21140
rect 13170 21088 13176 21140
rect 13228 21088 13234 21140
rect 13446 21088 13452 21140
rect 13504 21128 13510 21140
rect 13541 21131 13599 21137
rect 13541 21128 13553 21131
rect 13504 21100 13553 21128
rect 13504 21088 13510 21100
rect 13541 21097 13553 21100
rect 13587 21097 13599 21131
rect 13541 21091 13599 21097
rect 13725 21131 13783 21137
rect 13725 21097 13737 21131
rect 13771 21128 13783 21131
rect 14182 21128 14188 21140
rect 13771 21100 14188 21128
rect 13771 21097 13783 21100
rect 13725 21091 13783 21097
rect 14182 21088 14188 21100
rect 14240 21088 14246 21140
rect 14645 21131 14703 21137
rect 14384 21100 14596 21128
rect 13188 21060 13216 21088
rect 12452 21032 13216 21060
rect 8297 20995 8355 21001
rect 8297 20961 8309 20995
rect 8343 20992 8355 20995
rect 8941 20995 8999 21001
rect 8941 20992 8953 20995
rect 8343 20964 8953 20992
rect 8343 20961 8355 20964
rect 8297 20955 8355 20961
rect 8941 20961 8953 20964
rect 8987 20961 8999 20995
rect 8941 20955 8999 20961
rect 10321 20995 10379 21001
rect 10321 20961 10333 20995
rect 10367 20992 10379 20995
rect 10962 20992 10968 21004
rect 10367 20964 10968 20992
rect 10367 20961 10379 20964
rect 10321 20955 10379 20961
rect 10962 20952 10968 20964
rect 11020 20952 11026 21004
rect 8478 20884 8484 20936
rect 8536 20884 8542 20936
rect 8757 20927 8815 20933
rect 8757 20893 8769 20927
rect 8803 20924 8815 20927
rect 8803 20896 9720 20924
rect 8803 20893 8815 20896
rect 8757 20887 8815 20893
rect 9306 20748 9312 20800
rect 9364 20788 9370 20800
rect 9692 20797 9720 20896
rect 10410 20884 10416 20936
rect 10468 20884 10474 20936
rect 12452 20933 12480 21032
rect 14090 21020 14096 21072
rect 14148 21060 14154 21072
rect 14384 21060 14412 21100
rect 14148 21032 14412 21060
rect 14148 21020 14154 21032
rect 14458 21020 14464 21072
rect 14516 21020 14522 21072
rect 14568 21060 14596 21100
rect 14645 21097 14657 21131
rect 14691 21128 14703 21131
rect 14734 21128 14740 21140
rect 14691 21100 14740 21128
rect 14691 21097 14703 21100
rect 14645 21091 14703 21097
rect 14734 21088 14740 21100
rect 14792 21088 14798 21140
rect 14826 21088 14832 21140
rect 14884 21128 14890 21140
rect 15013 21131 15071 21137
rect 15013 21128 15025 21131
rect 14884 21100 15025 21128
rect 14884 21088 14890 21100
rect 15013 21097 15025 21100
rect 15059 21097 15071 21131
rect 15013 21091 15071 21097
rect 15289 21131 15347 21137
rect 15289 21097 15301 21131
rect 15335 21128 15347 21131
rect 15470 21128 15476 21140
rect 15335 21100 15476 21128
rect 15335 21097 15347 21100
rect 15289 21091 15347 21097
rect 15194 21060 15200 21072
rect 14568 21032 15200 21060
rect 15194 21020 15200 21032
rect 15252 21020 15258 21072
rect 12713 20995 12771 21001
rect 12713 20961 12725 20995
rect 12759 20992 12771 20995
rect 13449 20995 13507 21001
rect 13449 20992 13461 20995
rect 12759 20964 13461 20992
rect 12759 20961 12771 20964
rect 12713 20955 12771 20961
rect 13449 20961 13461 20964
rect 13495 20992 13507 20995
rect 13495 20964 13952 20992
rect 13495 20961 13507 20964
rect 13449 20955 13507 20961
rect 12437 20927 12495 20933
rect 12437 20893 12449 20927
rect 12483 20893 12495 20927
rect 12437 20887 12495 20893
rect 12802 20884 12808 20936
rect 12860 20884 12866 20936
rect 13814 20924 13820 20936
rect 13372 20896 13820 20924
rect 12526 20856 12532 20868
rect 11716 20828 12532 20856
rect 11716 20800 11744 20828
rect 12526 20816 12532 20828
rect 12584 20816 12590 20868
rect 13372 20856 13400 20896
rect 13814 20884 13820 20896
rect 13872 20884 13878 20936
rect 13924 20865 13952 20964
rect 14108 20924 14136 21020
rect 14274 20952 14280 21004
rect 14332 20992 14338 21004
rect 14553 20995 14611 21001
rect 14553 20992 14565 20995
rect 14332 20964 14565 20992
rect 14332 20952 14338 20964
rect 14553 20961 14565 20964
rect 14599 20961 14611 20995
rect 15304 20992 15332 21091
rect 15470 21088 15476 21100
rect 15528 21088 15534 21140
rect 15654 21088 15660 21140
rect 15712 21088 15718 21140
rect 15746 21088 15752 21140
rect 15804 21128 15810 21140
rect 20438 21128 20444 21140
rect 15804 21100 20444 21128
rect 15804 21088 15810 21100
rect 15378 21020 15384 21072
rect 15436 21020 15442 21072
rect 15838 21020 15844 21072
rect 15896 21020 15902 21072
rect 17494 21020 17500 21072
rect 17552 21020 17558 21072
rect 18690 21020 18696 21072
rect 18748 21020 18754 21072
rect 14553 20955 14611 20961
rect 14752 20964 15332 20992
rect 14185 20927 14243 20933
rect 14185 20924 14197 20927
rect 14108 20896 14197 20924
rect 14185 20893 14197 20896
rect 14231 20893 14243 20927
rect 14752 20924 14780 20964
rect 14185 20887 14243 20893
rect 14292 20896 14780 20924
rect 14829 20927 14887 20933
rect 14292 20865 14320 20896
rect 14829 20893 14841 20927
rect 14875 20924 14887 20927
rect 15396 20924 15424 21020
rect 14875 20896 15424 20924
rect 14875 20893 14887 20896
rect 14829 20887 14887 20893
rect 13909 20859 13967 20865
rect 12636 20828 13400 20856
rect 13464 20828 13676 20856
rect 9585 20791 9643 20797
rect 9585 20788 9597 20791
rect 9364 20760 9597 20788
rect 9364 20748 9370 20760
rect 9585 20757 9597 20760
rect 9631 20757 9643 20791
rect 9585 20751 9643 20757
rect 9677 20791 9735 20797
rect 9677 20757 9689 20791
rect 9723 20788 9735 20791
rect 11054 20788 11060 20800
rect 9723 20760 11060 20788
rect 9723 20757 9735 20760
rect 9677 20751 9735 20757
rect 11054 20748 11060 20760
rect 11112 20748 11118 20800
rect 11698 20748 11704 20800
rect 11756 20748 11762 20800
rect 12250 20748 12256 20800
rect 12308 20748 12314 20800
rect 12342 20748 12348 20800
rect 12400 20788 12406 20800
rect 12636 20788 12664 20828
rect 12400 20760 12664 20788
rect 12400 20748 12406 20760
rect 12986 20748 12992 20800
rect 13044 20788 13050 20800
rect 13464 20788 13492 20828
rect 13044 20760 13492 20788
rect 13648 20788 13676 20828
rect 13909 20825 13921 20859
rect 13955 20825 13967 20859
rect 13909 20819 13967 20825
rect 14277 20859 14335 20865
rect 14277 20825 14289 20859
rect 14323 20825 14335 20859
rect 14277 20819 14335 20825
rect 14461 20859 14519 20865
rect 14461 20825 14473 20859
rect 14507 20856 14519 20859
rect 15273 20859 15331 20865
rect 14507 20828 15240 20856
rect 14507 20825 14519 20828
rect 14461 20819 14519 20825
rect 13709 20791 13767 20797
rect 13709 20788 13721 20791
rect 13648 20760 13721 20788
rect 13044 20748 13050 20760
rect 13709 20757 13721 20760
rect 13755 20788 13767 20791
rect 14090 20788 14096 20800
rect 13755 20760 14096 20788
rect 13755 20757 13767 20760
rect 13709 20751 13767 20757
rect 14090 20748 14096 20760
rect 14148 20788 14154 20800
rect 15105 20791 15163 20797
rect 15105 20788 15117 20791
rect 14148 20760 15117 20788
rect 14148 20748 14154 20760
rect 15105 20757 15117 20760
rect 15151 20757 15163 20791
rect 15212 20788 15240 20828
rect 15273 20825 15285 20859
rect 15319 20856 15331 20859
rect 15378 20856 15384 20868
rect 15319 20828 15384 20856
rect 15319 20825 15331 20828
rect 15273 20819 15331 20825
rect 15378 20816 15384 20828
rect 15436 20816 15442 20868
rect 15473 20859 15531 20865
rect 15473 20825 15485 20859
rect 15519 20856 15531 20859
rect 15654 20856 15660 20868
rect 15519 20828 15660 20856
rect 15519 20825 15531 20828
rect 15473 20819 15531 20825
rect 15488 20788 15516 20819
rect 15654 20816 15660 20828
rect 15712 20816 15718 20868
rect 15856 20856 15884 21020
rect 17512 20992 17540 21020
rect 18800 20992 18828 21100
rect 20438 21088 20444 21100
rect 20496 21088 20502 21140
rect 20622 21088 20628 21140
rect 20680 21088 20686 21140
rect 22278 21088 22284 21140
rect 22336 21128 22342 21140
rect 22554 21128 22560 21140
rect 22336 21100 22560 21128
rect 22336 21088 22342 21100
rect 22554 21088 22560 21100
rect 22612 21088 22618 21140
rect 23474 21088 23480 21140
rect 23532 21128 23538 21140
rect 23753 21131 23811 21137
rect 23753 21128 23765 21131
rect 23532 21100 23765 21128
rect 23532 21088 23538 21100
rect 23753 21097 23765 21100
rect 23799 21097 23811 21131
rect 23753 21091 23811 21097
rect 19889 21063 19947 21069
rect 19889 21029 19901 21063
rect 19935 21060 19947 21063
rect 20162 21060 20168 21072
rect 19935 21032 20168 21060
rect 19935 21029 19947 21032
rect 19889 21023 19947 21029
rect 20162 21020 20168 21032
rect 20220 21020 20226 21072
rect 20640 20992 20668 21088
rect 21726 21020 21732 21072
rect 21784 21060 21790 21072
rect 21784 21032 21956 21060
rect 21784 21020 21790 21032
rect 21928 21001 21956 21032
rect 17512 20964 17908 20992
rect 16482 20884 16488 20936
rect 16540 20924 16546 20936
rect 16770 20927 16828 20933
rect 16770 20924 16782 20927
rect 16540 20896 16782 20924
rect 16540 20884 16546 20896
rect 16770 20893 16782 20896
rect 16816 20893 16828 20927
rect 16770 20887 16828 20893
rect 16942 20884 16948 20936
rect 17000 20924 17006 20936
rect 17037 20927 17095 20933
rect 17037 20924 17049 20927
rect 17000 20896 17049 20924
rect 17000 20884 17006 20896
rect 17037 20893 17049 20896
rect 17083 20924 17095 20927
rect 17678 20924 17684 20936
rect 17083 20896 17684 20924
rect 17083 20893 17095 20896
rect 17037 20887 17095 20893
rect 17678 20884 17684 20896
rect 17736 20884 17742 20936
rect 17880 20933 17908 20964
rect 18708 20964 18828 20992
rect 20562 20964 20668 20992
rect 21913 20995 21971 21001
rect 18708 20933 18736 20964
rect 21913 20961 21925 20995
rect 21959 20961 21971 20995
rect 21913 20955 21971 20961
rect 17865 20927 17923 20933
rect 17865 20893 17877 20927
rect 17911 20893 17923 20927
rect 17865 20887 17923 20893
rect 18049 20927 18107 20933
rect 18049 20893 18061 20927
rect 18095 20893 18107 20927
rect 18049 20887 18107 20893
rect 18693 20927 18751 20933
rect 18693 20893 18705 20927
rect 18739 20893 18751 20927
rect 18969 20927 19027 20933
rect 18969 20924 18981 20927
rect 18693 20887 18751 20893
rect 18800 20896 18981 20924
rect 15856 20828 16620 20856
rect 15212 20760 15516 20788
rect 16592 20788 16620 20828
rect 16666 20816 16672 20868
rect 16724 20856 16730 20868
rect 18064 20856 18092 20887
rect 18800 20868 18828 20896
rect 18969 20893 18981 20896
rect 19015 20893 19027 20927
rect 18969 20887 19027 20893
rect 20070 20884 20076 20936
rect 20128 20884 20134 20936
rect 20346 20884 20352 20936
rect 20404 20924 20410 20936
rect 20625 20927 20683 20933
rect 20625 20924 20637 20927
rect 20404 20896 20637 20924
rect 20404 20884 20410 20896
rect 20625 20893 20637 20896
rect 20671 20893 20683 20927
rect 20625 20887 20683 20893
rect 20714 20884 20720 20936
rect 20772 20884 20778 20936
rect 21542 20884 21548 20936
rect 21600 20884 21606 20936
rect 21726 20884 21732 20936
rect 21784 20884 21790 20936
rect 21821 20927 21879 20933
rect 21821 20893 21833 20927
rect 21867 20893 21879 20927
rect 21821 20887 21879 20893
rect 22097 20927 22155 20933
rect 22097 20893 22109 20927
rect 22143 20924 22155 20927
rect 22278 20924 22284 20936
rect 22143 20896 22284 20924
rect 22143 20893 22155 20896
rect 22097 20887 22155 20893
rect 16724 20828 18092 20856
rect 16724 20816 16730 20828
rect 18782 20816 18788 20868
rect 18840 20816 18846 20868
rect 21836 20856 21864 20887
rect 22278 20884 22284 20896
rect 22336 20884 22342 20936
rect 22370 20884 22376 20936
rect 22428 20924 22434 20936
rect 22428 20896 22876 20924
rect 22428 20884 22434 20896
rect 22848 20868 22876 20896
rect 22640 20859 22698 20865
rect 21836 20828 22600 20856
rect 17957 20791 18015 20797
rect 17957 20788 17969 20791
rect 16592 20760 17969 20788
rect 15105 20751 15163 20757
rect 17957 20757 17969 20760
rect 18003 20757 18015 20791
rect 17957 20751 18015 20757
rect 18874 20748 18880 20800
rect 18932 20748 18938 20800
rect 22278 20748 22284 20800
rect 22336 20748 22342 20800
rect 22572 20788 22600 20828
rect 22640 20825 22652 20859
rect 22686 20856 22698 20859
rect 22738 20856 22744 20868
rect 22686 20828 22744 20856
rect 22686 20825 22698 20828
rect 22640 20819 22698 20825
rect 22738 20816 22744 20828
rect 22796 20816 22802 20868
rect 22830 20816 22836 20868
rect 22888 20816 22894 20868
rect 23566 20788 23572 20800
rect 22572 20760 23572 20788
rect 23566 20748 23572 20760
rect 23624 20748 23630 20800
rect 1104 20698 35027 20720
rect 1104 20646 9390 20698
rect 9442 20646 9454 20698
rect 9506 20646 9518 20698
rect 9570 20646 9582 20698
rect 9634 20646 9646 20698
rect 9698 20646 17831 20698
rect 17883 20646 17895 20698
rect 17947 20646 17959 20698
rect 18011 20646 18023 20698
rect 18075 20646 18087 20698
rect 18139 20646 26272 20698
rect 26324 20646 26336 20698
rect 26388 20646 26400 20698
rect 26452 20646 26464 20698
rect 26516 20646 26528 20698
rect 26580 20646 34713 20698
rect 34765 20646 34777 20698
rect 34829 20646 34841 20698
rect 34893 20646 34905 20698
rect 34957 20646 34969 20698
rect 35021 20646 35027 20698
rect 1104 20624 35027 20646
rect 8478 20544 8484 20596
rect 8536 20584 8542 20596
rect 9125 20587 9183 20593
rect 9125 20584 9137 20587
rect 8536 20556 9137 20584
rect 8536 20544 8542 20556
rect 9125 20553 9137 20556
rect 9171 20553 9183 20587
rect 9125 20547 9183 20553
rect 9214 20544 9220 20596
rect 9272 20544 9278 20596
rect 10689 20587 10747 20593
rect 10689 20553 10701 20587
rect 10735 20584 10747 20587
rect 10962 20584 10968 20596
rect 10735 20556 10968 20584
rect 10735 20553 10747 20556
rect 10689 20547 10747 20553
rect 10962 20544 10968 20556
rect 11020 20544 11026 20596
rect 11054 20544 11060 20596
rect 11112 20584 11118 20596
rect 11112 20556 12020 20584
rect 11112 20544 11118 20556
rect 9232 20516 9260 20544
rect 9140 20488 9260 20516
rect 8938 20408 8944 20460
rect 8996 20408 9002 20460
rect 9033 20451 9091 20457
rect 9033 20417 9045 20451
rect 9079 20448 9091 20451
rect 9140 20448 9168 20488
rect 9306 20476 9312 20528
rect 9364 20516 9370 20528
rect 11992 20525 12020 20556
rect 13446 20544 13452 20596
rect 13504 20544 13510 20596
rect 14182 20544 14188 20596
rect 14240 20544 14246 20596
rect 14918 20544 14924 20596
rect 14976 20584 14982 20596
rect 15105 20587 15163 20593
rect 15105 20584 15117 20587
rect 14976 20556 15117 20584
rect 14976 20544 14982 20556
rect 15105 20553 15117 20556
rect 15151 20553 15163 20587
rect 15105 20547 15163 20553
rect 15194 20544 15200 20596
rect 15252 20584 15258 20596
rect 15378 20584 15384 20596
rect 15252 20556 15384 20584
rect 15252 20544 15258 20556
rect 15378 20544 15384 20556
rect 15436 20584 15442 20596
rect 16390 20584 16396 20596
rect 15436 20556 16396 20584
rect 15436 20544 15442 20556
rect 16390 20544 16396 20556
rect 16448 20544 16454 20596
rect 20714 20584 20720 20596
rect 20364 20556 20720 20584
rect 9554 20519 9612 20525
rect 9554 20516 9566 20519
rect 9364 20488 9566 20516
rect 9364 20476 9370 20488
rect 9554 20485 9566 20488
rect 9600 20485 9612 20519
rect 11977 20519 12035 20525
rect 9554 20479 9612 20485
rect 11747 20485 11805 20491
rect 9079 20420 9168 20448
rect 9217 20451 9275 20457
rect 9079 20417 9091 20420
rect 9033 20411 9091 20417
rect 9217 20417 9229 20451
rect 9263 20448 9275 20451
rect 9950 20448 9956 20460
rect 9263 20420 9956 20448
rect 9263 20417 9275 20420
rect 9217 20411 9275 20417
rect 9950 20408 9956 20420
rect 10008 20408 10014 20460
rect 10042 20408 10048 20460
rect 10100 20448 10106 20460
rect 10965 20451 11023 20457
rect 10965 20448 10977 20451
rect 10100 20420 10977 20448
rect 10100 20408 10106 20420
rect 10965 20417 10977 20420
rect 11011 20417 11023 20451
rect 10965 20411 11023 20417
rect 11149 20451 11207 20457
rect 11149 20417 11161 20451
rect 11195 20448 11207 20451
rect 11747 20451 11759 20485
rect 11793 20451 11805 20485
rect 11977 20485 11989 20519
rect 12023 20485 12035 20519
rect 12342 20516 12348 20528
rect 11977 20479 12035 20485
rect 12083 20488 12348 20516
rect 11747 20448 11805 20451
rect 12083 20448 12111 20488
rect 12342 20476 12348 20488
rect 12400 20516 12406 20528
rect 13464 20516 13492 20544
rect 12400 20488 13492 20516
rect 16240 20519 16298 20525
rect 12400 20476 12406 20488
rect 16240 20485 16252 20519
rect 16286 20516 16298 20519
rect 16669 20519 16727 20525
rect 16669 20516 16681 20519
rect 16286 20488 16681 20516
rect 16286 20485 16298 20488
rect 16240 20479 16298 20485
rect 16669 20485 16681 20488
rect 16715 20485 16727 20519
rect 16669 20479 16727 20485
rect 19334 20476 19340 20528
rect 19392 20516 19398 20528
rect 19981 20519 20039 20525
rect 19981 20516 19993 20519
rect 19392 20488 19993 20516
rect 19392 20476 19398 20488
rect 19981 20485 19993 20488
rect 20027 20485 20039 20519
rect 19981 20479 20039 20485
rect 11195 20420 12111 20448
rect 12161 20451 12219 20457
rect 11195 20417 11207 20420
rect 11149 20411 11207 20417
rect 12161 20417 12173 20451
rect 12207 20448 12219 20451
rect 12250 20448 12256 20460
rect 12207 20420 12256 20448
rect 12207 20417 12219 20420
rect 12161 20411 12219 20417
rect 12250 20408 12256 20420
rect 12308 20408 12314 20460
rect 12526 20408 12532 20460
rect 12584 20448 12590 20460
rect 13078 20457 13084 20460
rect 12805 20451 12863 20457
rect 12805 20448 12817 20451
rect 12584 20420 12817 20448
rect 12584 20408 12590 20420
rect 12805 20417 12817 20420
rect 12851 20417 12863 20451
rect 12805 20411 12863 20417
rect 13072 20411 13084 20457
rect 13078 20408 13084 20411
rect 13136 20408 13142 20460
rect 17126 20408 17132 20460
rect 17184 20448 17190 20460
rect 20070 20448 20076 20460
rect 17184 20420 20076 20448
rect 17184 20408 17190 20420
rect 20070 20408 20076 20420
rect 20128 20408 20134 20460
rect 20364 20457 20392 20556
rect 20714 20544 20720 20556
rect 20772 20584 20778 20596
rect 20993 20587 21051 20593
rect 20993 20584 21005 20587
rect 20772 20556 21005 20584
rect 20772 20544 20778 20556
rect 20993 20553 21005 20556
rect 21039 20553 21051 20587
rect 20993 20547 21051 20553
rect 21174 20544 21180 20596
rect 21232 20584 21238 20596
rect 21232 20556 26234 20584
rect 21232 20544 21238 20556
rect 20806 20516 20812 20528
rect 20456 20488 20812 20516
rect 20257 20451 20315 20457
rect 20257 20417 20269 20451
rect 20303 20417 20315 20451
rect 20257 20411 20315 20417
rect 20349 20451 20407 20457
rect 20349 20417 20361 20451
rect 20395 20417 20407 20451
rect 20349 20411 20407 20417
rect 8956 20380 8984 20408
rect 9306 20380 9312 20392
rect 8956 20352 9312 20380
rect 9306 20340 9312 20352
rect 9364 20340 9370 20392
rect 11241 20383 11299 20389
rect 11241 20349 11253 20383
rect 11287 20349 11299 20383
rect 11241 20343 11299 20349
rect 11256 20312 11284 20343
rect 14366 20340 14372 20392
rect 14424 20340 14430 20392
rect 16485 20383 16543 20389
rect 16485 20349 16497 20383
rect 16531 20349 16543 20383
rect 16485 20343 16543 20349
rect 10244 20284 11192 20312
rect 11256 20284 11836 20312
rect 9214 20204 9220 20256
rect 9272 20244 9278 20256
rect 10244 20244 10272 20284
rect 9272 20216 10272 20244
rect 10781 20247 10839 20253
rect 9272 20204 9278 20216
rect 10781 20213 10793 20247
rect 10827 20244 10839 20247
rect 11054 20244 11060 20256
rect 10827 20216 11060 20244
rect 10827 20213 10839 20216
rect 10781 20207 10839 20213
rect 11054 20204 11060 20216
rect 11112 20204 11118 20256
rect 11164 20244 11192 20284
rect 11808 20253 11836 20284
rect 13814 20272 13820 20324
rect 13872 20312 13878 20324
rect 14550 20312 14556 20324
rect 13872 20284 14556 20312
rect 13872 20272 13878 20284
rect 14550 20272 14556 20284
rect 14608 20272 14614 20324
rect 16500 20312 16528 20343
rect 17218 20340 17224 20392
rect 17276 20340 17282 20392
rect 20272 20380 20300 20411
rect 20456 20380 20484 20488
rect 20806 20476 20812 20488
rect 20864 20476 20870 20528
rect 21836 20488 22600 20516
rect 21836 20460 21864 20488
rect 20533 20451 20591 20457
rect 20533 20417 20545 20451
rect 20579 20448 20591 20451
rect 20579 20420 20760 20448
rect 20579 20417 20591 20420
rect 20533 20411 20591 20417
rect 20272 20352 20484 20380
rect 16500 20284 17816 20312
rect 17788 20256 17816 20284
rect 11609 20247 11667 20253
rect 11609 20244 11621 20247
rect 11164 20216 11621 20244
rect 11609 20213 11621 20216
rect 11655 20213 11667 20247
rect 11609 20207 11667 20213
rect 11793 20247 11851 20253
rect 11793 20213 11805 20247
rect 11839 20244 11851 20247
rect 12434 20244 12440 20256
rect 11839 20216 12440 20244
rect 11839 20213 11851 20216
rect 11793 20207 11851 20213
rect 12434 20204 12440 20216
rect 12492 20204 12498 20256
rect 12710 20204 12716 20256
rect 12768 20204 12774 20256
rect 15010 20204 15016 20256
rect 15068 20204 15074 20256
rect 17770 20204 17776 20256
rect 17828 20244 17834 20256
rect 18509 20247 18567 20253
rect 18509 20244 18521 20247
rect 17828 20216 18521 20244
rect 17828 20204 17834 20216
rect 18509 20213 18521 20216
rect 18555 20213 18567 20247
rect 18509 20207 18567 20213
rect 20254 20204 20260 20256
rect 20312 20204 20318 20256
rect 20530 20204 20536 20256
rect 20588 20204 20594 20256
rect 20732 20244 20760 20420
rect 20809 20435 20867 20441
rect 20809 20401 20821 20435
rect 20855 20401 20867 20435
rect 21818 20408 21824 20460
rect 21876 20408 21882 20460
rect 22005 20451 22063 20457
rect 22005 20417 22017 20451
rect 22051 20448 22063 20451
rect 22186 20448 22192 20460
rect 22051 20420 22192 20448
rect 22051 20417 22063 20420
rect 22005 20411 22063 20417
rect 22186 20408 22192 20420
rect 22244 20408 22250 20460
rect 22278 20408 22284 20460
rect 22336 20448 22342 20460
rect 22465 20451 22523 20457
rect 22465 20448 22477 20451
rect 22336 20420 22477 20448
rect 22336 20408 22342 20420
rect 22465 20417 22477 20420
rect 22511 20417 22523 20451
rect 22465 20411 22523 20417
rect 20809 20395 20867 20401
rect 20824 20324 20852 20395
rect 21910 20340 21916 20392
rect 21968 20340 21974 20392
rect 22572 20380 22600 20488
rect 22738 20476 22744 20528
rect 22796 20516 22802 20528
rect 23109 20519 23167 20525
rect 23109 20516 23121 20519
rect 22796 20488 23121 20516
rect 22796 20476 22802 20488
rect 23109 20485 23121 20488
rect 23155 20485 23167 20519
rect 23109 20479 23167 20485
rect 23566 20476 23572 20528
rect 23624 20476 23630 20528
rect 23198 20408 23204 20460
rect 23256 20408 23262 20460
rect 23661 20451 23719 20457
rect 23661 20417 23673 20451
rect 23707 20417 23719 20451
rect 23661 20411 23719 20417
rect 23676 20380 23704 20411
rect 22572 20352 23704 20380
rect 20806 20272 20812 20324
rect 20864 20272 20870 20324
rect 21542 20312 21548 20324
rect 21100 20284 21548 20312
rect 21100 20244 21128 20284
rect 21542 20272 21548 20284
rect 21600 20312 21606 20324
rect 21928 20312 21956 20340
rect 21600 20284 21956 20312
rect 22373 20315 22431 20321
rect 21600 20272 21606 20284
rect 22373 20281 22385 20315
rect 22419 20312 22431 20315
rect 23477 20315 23535 20321
rect 23477 20312 23489 20315
rect 22419 20284 23489 20312
rect 22419 20281 22431 20284
rect 22373 20275 22431 20281
rect 23477 20281 23489 20284
rect 23523 20281 23535 20315
rect 23477 20275 23535 20281
rect 20732 20216 21128 20244
rect 21910 20204 21916 20256
rect 21968 20244 21974 20256
rect 22388 20244 22416 20275
rect 21968 20216 22416 20244
rect 21968 20204 21974 20216
rect 22462 20204 22468 20256
rect 22520 20244 22526 20256
rect 23339 20247 23397 20253
rect 23339 20244 23351 20247
rect 22520 20216 23351 20244
rect 22520 20204 22526 20216
rect 23339 20213 23351 20216
rect 23385 20213 23397 20247
rect 26206 20244 26234 20556
rect 33134 20244 33140 20256
rect 26206 20216 33140 20244
rect 23339 20207 23397 20213
rect 33134 20204 33140 20216
rect 33192 20204 33198 20256
rect 1104 20154 34868 20176
rect 1104 20102 5170 20154
rect 5222 20102 5234 20154
rect 5286 20102 5298 20154
rect 5350 20102 5362 20154
rect 5414 20102 5426 20154
rect 5478 20102 13611 20154
rect 13663 20102 13675 20154
rect 13727 20102 13739 20154
rect 13791 20102 13803 20154
rect 13855 20102 13867 20154
rect 13919 20102 22052 20154
rect 22104 20102 22116 20154
rect 22168 20102 22180 20154
rect 22232 20102 22244 20154
rect 22296 20102 22308 20154
rect 22360 20102 30493 20154
rect 30545 20102 30557 20154
rect 30609 20102 30621 20154
rect 30673 20102 30685 20154
rect 30737 20102 30749 20154
rect 30801 20102 34868 20154
rect 1104 20080 34868 20102
rect 9769 20043 9827 20049
rect 9769 20009 9781 20043
rect 9815 20040 9827 20043
rect 10042 20040 10048 20052
rect 9815 20012 10048 20040
rect 9815 20009 9827 20012
rect 9769 20003 9827 20009
rect 10042 20000 10048 20012
rect 10100 20000 10106 20052
rect 11698 20040 11704 20052
rect 10152 20012 11704 20040
rect 9306 19864 9312 19916
rect 9364 19904 9370 19916
rect 10152 19913 10180 20012
rect 11698 20000 11704 20012
rect 11756 20040 11762 20052
rect 11756 20012 13032 20040
rect 11756 20000 11762 20012
rect 11517 19975 11575 19981
rect 11517 19941 11529 19975
rect 11563 19972 11575 19975
rect 11882 19972 11888 19984
rect 11563 19944 11888 19972
rect 11563 19941 11575 19944
rect 11517 19935 11575 19941
rect 11882 19932 11888 19944
rect 11940 19932 11946 19984
rect 13004 19913 13032 20012
rect 13078 20000 13084 20052
rect 13136 20040 13142 20052
rect 13265 20043 13323 20049
rect 13265 20040 13277 20043
rect 13136 20012 13277 20040
rect 13136 20000 13142 20012
rect 13265 20009 13277 20012
rect 13311 20009 13323 20043
rect 13265 20003 13323 20009
rect 14550 20000 14556 20052
rect 14608 20040 14614 20052
rect 14608 20012 15240 20040
rect 14608 20000 14614 20012
rect 10137 19907 10195 19913
rect 10137 19904 10149 19907
rect 9364 19876 10149 19904
rect 9364 19864 9370 19876
rect 10137 19873 10149 19876
rect 10183 19873 10195 19907
rect 10137 19867 10195 19873
rect 12989 19907 13047 19913
rect 12989 19873 13001 19907
rect 13035 19904 13047 19907
rect 14185 19907 14243 19913
rect 14185 19904 14197 19907
rect 13035 19876 14197 19904
rect 13035 19873 13047 19876
rect 12989 19867 13047 19873
rect 14185 19873 14197 19876
rect 14231 19873 14243 19907
rect 14185 19867 14243 19873
rect 9585 19839 9643 19845
rect 9585 19805 9597 19839
rect 9631 19805 9643 19839
rect 9585 19799 9643 19805
rect 9600 19768 9628 19799
rect 9766 19796 9772 19848
rect 9824 19836 9830 19848
rect 10686 19836 10692 19848
rect 9824 19808 10692 19836
rect 9824 19796 9830 19808
rect 10686 19796 10692 19808
rect 10744 19796 10750 19848
rect 12710 19796 12716 19848
rect 12768 19845 12774 19848
rect 12768 19836 12780 19845
rect 13081 19839 13139 19845
rect 12768 19808 12813 19836
rect 12768 19799 12780 19808
rect 13081 19805 13093 19839
rect 13127 19836 13139 19839
rect 13170 19836 13176 19848
rect 13127 19808 13176 19836
rect 13127 19805 13139 19808
rect 13081 19799 13139 19805
rect 12768 19796 12774 19799
rect 13170 19796 13176 19808
rect 13228 19796 13234 19848
rect 13262 19796 13268 19848
rect 13320 19796 13326 19848
rect 14452 19839 14510 19845
rect 14452 19805 14464 19839
rect 14498 19836 14510 19839
rect 15010 19836 15016 19848
rect 14498 19808 15016 19836
rect 14498 19805 14510 19808
rect 14452 19799 14510 19805
rect 15010 19796 15016 19808
rect 15068 19796 15074 19848
rect 15212 19836 15240 20012
rect 15286 20000 15292 20052
rect 15344 20000 15350 20052
rect 15654 20000 15660 20052
rect 15712 20000 15718 20052
rect 16393 20043 16451 20049
rect 16393 20009 16405 20043
rect 16439 20040 16451 20043
rect 17218 20040 17224 20052
rect 16439 20012 17224 20040
rect 16439 20009 16451 20012
rect 16393 20003 16451 20009
rect 17218 20000 17224 20012
rect 17276 20000 17282 20052
rect 19061 20043 19119 20049
rect 19061 20009 19073 20043
rect 19107 20040 19119 20043
rect 19610 20040 19616 20052
rect 19107 20012 19616 20040
rect 19107 20009 19119 20012
rect 19061 20003 19119 20009
rect 19610 20000 19616 20012
rect 19668 20040 19674 20052
rect 20346 20040 20352 20052
rect 19668 20012 20352 20040
rect 19668 20000 19674 20012
rect 20346 20000 20352 20012
rect 20404 20000 20410 20052
rect 20530 20000 20536 20052
rect 20588 20000 20594 20052
rect 20806 20000 20812 20052
rect 20864 20000 20870 20052
rect 20901 20043 20959 20049
rect 20901 20009 20913 20043
rect 20947 20040 20959 20043
rect 20990 20040 20996 20052
rect 20947 20012 20996 20040
rect 20947 20009 20959 20012
rect 20901 20003 20959 20009
rect 20990 20000 20996 20012
rect 21048 20000 21054 20052
rect 21726 20000 21732 20052
rect 21784 20000 21790 20052
rect 22097 20043 22155 20049
rect 22097 20009 22109 20043
rect 22143 20040 22155 20043
rect 22462 20040 22468 20052
rect 22143 20012 22468 20040
rect 22143 20009 22155 20012
rect 22097 20003 22155 20009
rect 22462 20000 22468 20012
rect 22520 20000 22526 20052
rect 22646 20000 22652 20052
rect 22704 20000 22710 20052
rect 23198 20000 23204 20052
rect 23256 20000 23262 20052
rect 15304 19972 15332 20000
rect 15565 19975 15623 19981
rect 15565 19972 15577 19975
rect 15304 19944 15577 19972
rect 15565 19941 15577 19944
rect 15611 19941 15623 19975
rect 20548 19972 20576 20000
rect 20548 19944 22508 19972
rect 15565 19935 15623 19941
rect 15580 19904 15608 19935
rect 16209 19907 16267 19913
rect 16209 19904 16221 19907
rect 15580 19876 16221 19904
rect 16209 19873 16221 19876
rect 16255 19873 16267 19907
rect 17126 19904 17132 19916
rect 16209 19867 16267 19873
rect 16316 19876 17132 19904
rect 16316 19836 16344 19876
rect 15212 19808 16344 19836
rect 16390 19796 16396 19848
rect 16448 19796 16454 19848
rect 16592 19845 16620 19876
rect 17126 19864 17132 19876
rect 17184 19864 17190 19916
rect 22370 19904 22376 19916
rect 20456 19876 22376 19904
rect 16577 19839 16635 19845
rect 16577 19805 16589 19839
rect 16623 19805 16635 19839
rect 16577 19799 16635 19805
rect 17681 19839 17739 19845
rect 17681 19805 17693 19839
rect 17727 19836 17739 19839
rect 17770 19836 17776 19848
rect 17727 19808 17776 19836
rect 17727 19805 17739 19808
rect 17681 19799 17739 19805
rect 17770 19796 17776 19808
rect 17828 19836 17834 19848
rect 19429 19839 19487 19845
rect 19429 19836 19441 19839
rect 17828 19808 19441 19836
rect 17828 19796 17834 19808
rect 19429 19805 19441 19808
rect 19475 19836 19487 19839
rect 20456 19836 20484 19876
rect 22370 19864 22376 19876
rect 22428 19864 22434 19916
rect 19475 19808 20484 19836
rect 19475 19805 19487 19808
rect 19429 19799 19487 19805
rect 21082 19796 21088 19848
rect 21140 19796 21146 19848
rect 21177 19839 21235 19845
rect 21177 19805 21189 19839
rect 21223 19805 21235 19839
rect 21177 19799 21235 19805
rect 21545 19839 21603 19845
rect 21545 19805 21557 19839
rect 21591 19836 21603 19839
rect 21818 19836 21824 19848
rect 21591 19808 21824 19836
rect 21591 19805 21603 19808
rect 21545 19799 21603 19805
rect 9950 19768 9956 19780
rect 9600 19740 9956 19768
rect 9950 19728 9956 19740
rect 10008 19728 10014 19780
rect 10404 19771 10462 19777
rect 10404 19737 10416 19771
rect 10450 19768 10462 19771
rect 10594 19768 10600 19780
rect 10450 19740 10600 19768
rect 10450 19737 10462 19740
rect 10404 19731 10462 19737
rect 10594 19728 10600 19740
rect 10652 19728 10658 19780
rect 17948 19771 18006 19777
rect 10704 19740 17264 19768
rect 7650 19660 7656 19712
rect 7708 19700 7714 19712
rect 10704 19700 10732 19740
rect 7708 19672 10732 19700
rect 11609 19703 11667 19709
rect 7708 19660 7714 19672
rect 11609 19669 11621 19703
rect 11655 19700 11667 19703
rect 12802 19700 12808 19712
rect 11655 19672 12808 19700
rect 11655 19669 11667 19672
rect 11609 19663 11667 19669
rect 12802 19660 12808 19672
rect 12860 19660 12866 19712
rect 17236 19700 17264 19740
rect 17948 19737 17960 19771
rect 17994 19768 18006 19771
rect 18414 19768 18420 19780
rect 17994 19740 18420 19768
rect 17994 19737 18006 19740
rect 17948 19731 18006 19737
rect 18414 19728 18420 19740
rect 18472 19728 18478 19780
rect 19696 19771 19754 19777
rect 19696 19737 19708 19771
rect 19742 19768 19754 19771
rect 20254 19768 20260 19780
rect 19742 19740 20260 19768
rect 19742 19737 19754 19740
rect 19696 19731 19754 19737
rect 20254 19728 20260 19740
rect 20312 19728 20318 19780
rect 21192 19768 21220 19799
rect 21818 19796 21824 19808
rect 21876 19796 21882 19848
rect 21910 19796 21916 19848
rect 21968 19796 21974 19848
rect 22480 19845 22508 19944
rect 22189 19839 22247 19845
rect 22189 19805 22201 19839
rect 22235 19836 22247 19839
rect 22465 19839 22523 19845
rect 22235 19808 22324 19836
rect 22235 19805 22247 19808
rect 22189 19799 22247 19805
rect 22296 19780 22324 19808
rect 22465 19805 22477 19839
rect 22511 19805 22523 19839
rect 22465 19799 22523 19805
rect 21192 19740 22094 19768
rect 21174 19700 21180 19712
rect 17236 19672 21180 19700
rect 21174 19660 21180 19672
rect 21232 19660 21238 19712
rect 22066 19700 22094 19740
rect 22278 19728 22284 19780
rect 22336 19768 22342 19780
rect 23216 19768 23244 20000
rect 33134 19796 33140 19848
rect 33192 19796 33198 19848
rect 22336 19740 23244 19768
rect 34333 19771 34391 19777
rect 22336 19728 22342 19740
rect 34333 19737 34345 19771
rect 34379 19768 34391 19771
rect 34606 19768 34612 19780
rect 34379 19740 34612 19768
rect 34379 19737 34391 19740
rect 34333 19731 34391 19737
rect 34606 19728 34612 19740
rect 34664 19728 34670 19780
rect 22646 19700 22652 19712
rect 22066 19672 22652 19700
rect 22646 19660 22652 19672
rect 22704 19660 22710 19712
rect 1104 19610 35027 19632
rect 1104 19558 9390 19610
rect 9442 19558 9454 19610
rect 9506 19558 9518 19610
rect 9570 19558 9582 19610
rect 9634 19558 9646 19610
rect 9698 19558 17831 19610
rect 17883 19558 17895 19610
rect 17947 19558 17959 19610
rect 18011 19558 18023 19610
rect 18075 19558 18087 19610
rect 18139 19558 26272 19610
rect 26324 19558 26336 19610
rect 26388 19558 26400 19610
rect 26452 19558 26464 19610
rect 26516 19558 26528 19610
rect 26580 19558 34713 19610
rect 34765 19558 34777 19610
rect 34829 19558 34841 19610
rect 34893 19558 34905 19610
rect 34957 19558 34969 19610
rect 35021 19558 35027 19610
rect 1104 19536 35027 19558
rect 10594 19456 10600 19508
rect 10652 19456 10658 19508
rect 10686 19456 10692 19508
rect 10744 19496 10750 19508
rect 12253 19499 12311 19505
rect 12253 19496 12265 19499
rect 10744 19468 12265 19496
rect 10744 19456 10750 19468
rect 12253 19465 12265 19468
rect 12299 19465 12311 19499
rect 12434 19496 12440 19508
rect 12253 19459 12311 19465
rect 12360 19468 12440 19496
rect 11517 19431 11575 19437
rect 11517 19397 11529 19431
rect 11563 19428 11575 19431
rect 12360 19428 12388 19468
rect 12434 19456 12440 19468
rect 12492 19456 12498 19508
rect 14277 19499 14335 19505
rect 14277 19465 14289 19499
rect 14323 19496 14335 19499
rect 14366 19496 14372 19508
rect 14323 19468 14372 19496
rect 14323 19465 14335 19468
rect 14277 19459 14335 19465
rect 14366 19456 14372 19468
rect 14424 19456 14430 19508
rect 14458 19456 14464 19508
rect 14516 19456 14522 19508
rect 16390 19456 16396 19508
rect 16448 19456 16454 19508
rect 18414 19456 18420 19508
rect 18472 19456 18478 19508
rect 18874 19456 18880 19508
rect 18932 19496 18938 19508
rect 18969 19499 19027 19505
rect 18969 19496 18981 19499
rect 18932 19468 18981 19496
rect 18932 19456 18938 19468
rect 18969 19465 18981 19468
rect 19015 19465 19027 19499
rect 18969 19459 19027 19465
rect 20714 19456 20720 19508
rect 20772 19456 20778 19508
rect 21542 19456 21548 19508
rect 21600 19456 21606 19508
rect 21637 19499 21695 19505
rect 21637 19465 21649 19499
rect 21683 19496 21695 19499
rect 22278 19496 22284 19508
rect 21683 19468 22284 19496
rect 21683 19465 21695 19468
rect 21637 19459 21695 19465
rect 22278 19456 22284 19468
rect 22336 19456 22342 19508
rect 11563 19400 12572 19428
rect 11563 19397 11575 19400
rect 11517 19391 11575 19397
rect 11054 19320 11060 19372
rect 11112 19360 11118 19372
rect 11112 19332 11192 19360
rect 11112 19320 11118 19332
rect 11164 19301 11192 19332
rect 11882 19320 11888 19372
rect 11940 19360 11946 19372
rect 12069 19363 12127 19369
rect 12069 19360 12081 19363
rect 11940 19332 12081 19360
rect 11940 19320 11946 19332
rect 12069 19329 12081 19332
rect 12115 19329 12127 19363
rect 12069 19323 12127 19329
rect 12342 19320 12348 19372
rect 12400 19360 12406 19372
rect 12544 19369 12572 19400
rect 12437 19363 12495 19369
rect 12437 19360 12449 19363
rect 12400 19332 12449 19360
rect 12400 19320 12406 19332
rect 12437 19329 12449 19332
rect 12483 19329 12495 19363
rect 12437 19323 12495 19329
rect 12529 19363 12587 19369
rect 12529 19329 12541 19363
rect 12575 19329 12587 19363
rect 12529 19323 12587 19329
rect 14277 19363 14335 19369
rect 14277 19329 14289 19363
rect 14323 19360 14335 19363
rect 14476 19360 14504 19456
rect 14550 19388 14556 19440
rect 14608 19388 14614 19440
rect 14323 19332 14504 19360
rect 14323 19329 14335 19332
rect 14277 19323 14335 19329
rect 14918 19320 14924 19372
rect 14976 19320 14982 19372
rect 15749 19363 15807 19369
rect 15749 19329 15761 19363
rect 15795 19360 15807 19363
rect 16408 19360 16436 19456
rect 15795 19332 16436 19360
rect 18601 19363 18659 19369
rect 15795 19329 15807 19332
rect 15749 19323 15807 19329
rect 18601 19329 18613 19363
rect 18647 19360 18659 19363
rect 18690 19360 18696 19372
rect 18647 19332 18696 19360
rect 18647 19329 18659 19332
rect 18601 19323 18659 19329
rect 18690 19320 18696 19332
rect 18748 19320 18754 19372
rect 18782 19320 18788 19372
rect 18840 19320 18846 19372
rect 18892 19369 18920 19456
rect 18877 19363 18935 19369
rect 18877 19329 18889 19363
rect 18923 19329 18935 19363
rect 18877 19323 18935 19329
rect 19610 19320 19616 19372
rect 19668 19320 19674 19372
rect 20732 19360 20760 19456
rect 20809 19363 20867 19369
rect 20809 19360 20821 19363
rect 20732 19332 20821 19360
rect 20809 19329 20821 19332
rect 20855 19360 20867 19363
rect 21269 19363 21327 19369
rect 21269 19360 21281 19363
rect 20855 19332 21281 19360
rect 20855 19329 20867 19332
rect 20809 19323 20867 19329
rect 21269 19329 21281 19332
rect 21315 19329 21327 19363
rect 21269 19323 21327 19329
rect 21453 19363 21511 19369
rect 21453 19329 21465 19363
rect 21499 19360 21511 19363
rect 21560 19360 21588 19456
rect 21499 19332 21588 19360
rect 21499 19329 21511 19332
rect 21453 19323 21511 19329
rect 11149 19295 11207 19301
rect 11149 19261 11161 19295
rect 11195 19261 11207 19295
rect 11149 19255 11207 19261
rect 14090 19252 14096 19304
rect 14148 19292 14154 19304
rect 14369 19295 14427 19301
rect 14369 19292 14381 19295
rect 14148 19264 14381 19292
rect 14148 19252 14154 19264
rect 14369 19261 14381 19264
rect 14415 19261 14427 19295
rect 14936 19292 14964 19320
rect 15473 19295 15531 19301
rect 15473 19292 15485 19295
rect 14936 19264 15485 19292
rect 14369 19255 14427 19261
rect 15473 19261 15485 19264
rect 15519 19261 15531 19295
rect 15473 19255 15531 19261
rect 20717 19295 20775 19301
rect 20717 19261 20729 19295
rect 20763 19292 20775 19295
rect 20898 19292 20904 19304
rect 20763 19264 20904 19292
rect 20763 19261 20775 19264
rect 20717 19255 20775 19261
rect 20898 19252 20904 19264
rect 20956 19252 20962 19304
rect 1104 19066 34868 19088
rect 1104 19014 5170 19066
rect 5222 19014 5234 19066
rect 5286 19014 5298 19066
rect 5350 19014 5362 19066
rect 5414 19014 5426 19066
rect 5478 19014 13611 19066
rect 13663 19014 13675 19066
rect 13727 19014 13739 19066
rect 13791 19014 13803 19066
rect 13855 19014 13867 19066
rect 13919 19014 22052 19066
rect 22104 19014 22116 19066
rect 22168 19014 22180 19066
rect 22232 19014 22244 19066
rect 22296 19014 22308 19066
rect 22360 19014 30493 19066
rect 30545 19014 30557 19066
rect 30609 19014 30621 19066
rect 30673 19014 30685 19066
rect 30737 19014 30749 19066
rect 30801 19014 34868 19066
rect 1104 18992 34868 19014
rect 1104 18522 35027 18544
rect 1104 18470 9390 18522
rect 9442 18470 9454 18522
rect 9506 18470 9518 18522
rect 9570 18470 9582 18522
rect 9634 18470 9646 18522
rect 9698 18470 17831 18522
rect 17883 18470 17895 18522
rect 17947 18470 17959 18522
rect 18011 18470 18023 18522
rect 18075 18470 18087 18522
rect 18139 18470 26272 18522
rect 26324 18470 26336 18522
rect 26388 18470 26400 18522
rect 26452 18470 26464 18522
rect 26516 18470 26528 18522
rect 26580 18470 34713 18522
rect 34765 18470 34777 18522
rect 34829 18470 34841 18522
rect 34893 18470 34905 18522
rect 34957 18470 34969 18522
rect 35021 18470 35027 18522
rect 1104 18448 35027 18470
rect 1104 17978 34868 18000
rect 1104 17926 5170 17978
rect 5222 17926 5234 17978
rect 5286 17926 5298 17978
rect 5350 17926 5362 17978
rect 5414 17926 5426 17978
rect 5478 17926 13611 17978
rect 13663 17926 13675 17978
rect 13727 17926 13739 17978
rect 13791 17926 13803 17978
rect 13855 17926 13867 17978
rect 13919 17926 22052 17978
rect 22104 17926 22116 17978
rect 22168 17926 22180 17978
rect 22232 17926 22244 17978
rect 22296 17926 22308 17978
rect 22360 17926 30493 17978
rect 30545 17926 30557 17978
rect 30609 17926 30621 17978
rect 30673 17926 30685 17978
rect 30737 17926 30749 17978
rect 30801 17926 34868 17978
rect 1104 17904 34868 17926
rect 1104 17434 35027 17456
rect 1104 17382 9390 17434
rect 9442 17382 9454 17434
rect 9506 17382 9518 17434
rect 9570 17382 9582 17434
rect 9634 17382 9646 17434
rect 9698 17382 17831 17434
rect 17883 17382 17895 17434
rect 17947 17382 17959 17434
rect 18011 17382 18023 17434
rect 18075 17382 18087 17434
rect 18139 17382 26272 17434
rect 26324 17382 26336 17434
rect 26388 17382 26400 17434
rect 26452 17382 26464 17434
rect 26516 17382 26528 17434
rect 26580 17382 34713 17434
rect 34765 17382 34777 17434
rect 34829 17382 34841 17434
rect 34893 17382 34905 17434
rect 34957 17382 34969 17434
rect 35021 17382 35027 17434
rect 1104 17360 35027 17382
rect 1104 16890 34868 16912
rect 1104 16838 5170 16890
rect 5222 16838 5234 16890
rect 5286 16838 5298 16890
rect 5350 16838 5362 16890
rect 5414 16838 5426 16890
rect 5478 16838 13611 16890
rect 13663 16838 13675 16890
rect 13727 16838 13739 16890
rect 13791 16838 13803 16890
rect 13855 16838 13867 16890
rect 13919 16838 22052 16890
rect 22104 16838 22116 16890
rect 22168 16838 22180 16890
rect 22232 16838 22244 16890
rect 22296 16838 22308 16890
rect 22360 16838 30493 16890
rect 30545 16838 30557 16890
rect 30609 16838 30621 16890
rect 30673 16838 30685 16890
rect 30737 16838 30749 16890
rect 30801 16838 34868 16890
rect 1104 16816 34868 16838
rect 1104 16346 35027 16368
rect 1104 16294 9390 16346
rect 9442 16294 9454 16346
rect 9506 16294 9518 16346
rect 9570 16294 9582 16346
rect 9634 16294 9646 16346
rect 9698 16294 17831 16346
rect 17883 16294 17895 16346
rect 17947 16294 17959 16346
rect 18011 16294 18023 16346
rect 18075 16294 18087 16346
rect 18139 16294 26272 16346
rect 26324 16294 26336 16346
rect 26388 16294 26400 16346
rect 26452 16294 26464 16346
rect 26516 16294 26528 16346
rect 26580 16294 34713 16346
rect 34765 16294 34777 16346
rect 34829 16294 34841 16346
rect 34893 16294 34905 16346
rect 34957 16294 34969 16346
rect 35021 16294 35027 16346
rect 1104 16272 35027 16294
rect 1104 15802 34868 15824
rect 1104 15750 5170 15802
rect 5222 15750 5234 15802
rect 5286 15750 5298 15802
rect 5350 15750 5362 15802
rect 5414 15750 5426 15802
rect 5478 15750 13611 15802
rect 13663 15750 13675 15802
rect 13727 15750 13739 15802
rect 13791 15750 13803 15802
rect 13855 15750 13867 15802
rect 13919 15750 22052 15802
rect 22104 15750 22116 15802
rect 22168 15750 22180 15802
rect 22232 15750 22244 15802
rect 22296 15750 22308 15802
rect 22360 15750 30493 15802
rect 30545 15750 30557 15802
rect 30609 15750 30621 15802
rect 30673 15750 30685 15802
rect 30737 15750 30749 15802
rect 30801 15750 34868 15802
rect 1104 15728 34868 15750
rect 1104 15258 35027 15280
rect 1104 15206 9390 15258
rect 9442 15206 9454 15258
rect 9506 15206 9518 15258
rect 9570 15206 9582 15258
rect 9634 15206 9646 15258
rect 9698 15206 17831 15258
rect 17883 15206 17895 15258
rect 17947 15206 17959 15258
rect 18011 15206 18023 15258
rect 18075 15206 18087 15258
rect 18139 15206 26272 15258
rect 26324 15206 26336 15258
rect 26388 15206 26400 15258
rect 26452 15206 26464 15258
rect 26516 15206 26528 15258
rect 26580 15206 34713 15258
rect 34765 15206 34777 15258
rect 34829 15206 34841 15258
rect 34893 15206 34905 15258
rect 34957 15206 34969 15258
rect 35021 15206 35027 15258
rect 1104 15184 35027 15206
rect 1104 14714 34868 14736
rect 1104 14662 5170 14714
rect 5222 14662 5234 14714
rect 5286 14662 5298 14714
rect 5350 14662 5362 14714
rect 5414 14662 5426 14714
rect 5478 14662 13611 14714
rect 13663 14662 13675 14714
rect 13727 14662 13739 14714
rect 13791 14662 13803 14714
rect 13855 14662 13867 14714
rect 13919 14662 22052 14714
rect 22104 14662 22116 14714
rect 22168 14662 22180 14714
rect 22232 14662 22244 14714
rect 22296 14662 22308 14714
rect 22360 14662 30493 14714
rect 30545 14662 30557 14714
rect 30609 14662 30621 14714
rect 30673 14662 30685 14714
rect 30737 14662 30749 14714
rect 30801 14662 34868 14714
rect 1104 14640 34868 14662
rect 1578 14560 1584 14612
rect 1636 14560 1642 14612
rect 934 14356 940 14408
rect 992 14396 998 14408
rect 1397 14399 1455 14405
rect 1397 14396 1409 14399
rect 992 14368 1409 14396
rect 992 14356 998 14368
rect 1397 14365 1409 14368
rect 1443 14365 1455 14399
rect 1397 14359 1455 14365
rect 1104 14170 35027 14192
rect 1104 14118 9390 14170
rect 9442 14118 9454 14170
rect 9506 14118 9518 14170
rect 9570 14118 9582 14170
rect 9634 14118 9646 14170
rect 9698 14118 17831 14170
rect 17883 14118 17895 14170
rect 17947 14118 17959 14170
rect 18011 14118 18023 14170
rect 18075 14118 18087 14170
rect 18139 14118 26272 14170
rect 26324 14118 26336 14170
rect 26388 14118 26400 14170
rect 26452 14118 26464 14170
rect 26516 14118 26528 14170
rect 26580 14118 34713 14170
rect 34765 14118 34777 14170
rect 34829 14118 34841 14170
rect 34893 14118 34905 14170
rect 34957 14118 34969 14170
rect 35021 14118 35027 14170
rect 1104 14096 35027 14118
rect 1104 13626 34868 13648
rect 1104 13574 5170 13626
rect 5222 13574 5234 13626
rect 5286 13574 5298 13626
rect 5350 13574 5362 13626
rect 5414 13574 5426 13626
rect 5478 13574 13611 13626
rect 13663 13574 13675 13626
rect 13727 13574 13739 13626
rect 13791 13574 13803 13626
rect 13855 13574 13867 13626
rect 13919 13574 22052 13626
rect 22104 13574 22116 13626
rect 22168 13574 22180 13626
rect 22232 13574 22244 13626
rect 22296 13574 22308 13626
rect 22360 13574 30493 13626
rect 30545 13574 30557 13626
rect 30609 13574 30621 13626
rect 30673 13574 30685 13626
rect 30737 13574 30749 13626
rect 30801 13574 34868 13626
rect 1104 13552 34868 13574
rect 34517 13311 34575 13317
rect 34517 13277 34529 13311
rect 34563 13308 34575 13311
rect 34563 13280 35204 13308
rect 34563 13277 34575 13280
rect 34517 13271 34575 13277
rect 35176 13184 35204 13280
rect 24026 13132 24032 13184
rect 24084 13172 24090 13184
rect 34333 13175 34391 13181
rect 34333 13172 34345 13175
rect 24084 13144 34345 13172
rect 24084 13132 24090 13144
rect 34333 13141 34345 13144
rect 34379 13141 34391 13175
rect 34333 13135 34391 13141
rect 35158 13132 35164 13184
rect 35216 13132 35222 13184
rect 1104 13082 35027 13104
rect 1104 13030 9390 13082
rect 9442 13030 9454 13082
rect 9506 13030 9518 13082
rect 9570 13030 9582 13082
rect 9634 13030 9646 13082
rect 9698 13030 17831 13082
rect 17883 13030 17895 13082
rect 17947 13030 17959 13082
rect 18011 13030 18023 13082
rect 18075 13030 18087 13082
rect 18139 13030 26272 13082
rect 26324 13030 26336 13082
rect 26388 13030 26400 13082
rect 26452 13030 26464 13082
rect 26516 13030 26528 13082
rect 26580 13030 34713 13082
rect 34765 13030 34777 13082
rect 34829 13030 34841 13082
rect 34893 13030 34905 13082
rect 34957 13030 34969 13082
rect 35021 13030 35027 13082
rect 1104 13008 35027 13030
rect 1104 12538 34868 12560
rect 1104 12486 5170 12538
rect 5222 12486 5234 12538
rect 5286 12486 5298 12538
rect 5350 12486 5362 12538
rect 5414 12486 5426 12538
rect 5478 12486 13611 12538
rect 13663 12486 13675 12538
rect 13727 12486 13739 12538
rect 13791 12486 13803 12538
rect 13855 12486 13867 12538
rect 13919 12486 22052 12538
rect 22104 12486 22116 12538
rect 22168 12486 22180 12538
rect 22232 12486 22244 12538
rect 22296 12486 22308 12538
rect 22360 12486 30493 12538
rect 30545 12486 30557 12538
rect 30609 12486 30621 12538
rect 30673 12486 30685 12538
rect 30737 12486 30749 12538
rect 30801 12486 34868 12538
rect 1104 12464 34868 12486
rect 1104 11994 35027 12016
rect 1104 11942 9390 11994
rect 9442 11942 9454 11994
rect 9506 11942 9518 11994
rect 9570 11942 9582 11994
rect 9634 11942 9646 11994
rect 9698 11942 17831 11994
rect 17883 11942 17895 11994
rect 17947 11942 17959 11994
rect 18011 11942 18023 11994
rect 18075 11942 18087 11994
rect 18139 11942 26272 11994
rect 26324 11942 26336 11994
rect 26388 11942 26400 11994
rect 26452 11942 26464 11994
rect 26516 11942 26528 11994
rect 26580 11942 34713 11994
rect 34765 11942 34777 11994
rect 34829 11942 34841 11994
rect 34893 11942 34905 11994
rect 34957 11942 34969 11994
rect 35021 11942 35027 11994
rect 1104 11920 35027 11942
rect 1104 11450 34868 11472
rect 1104 11398 5170 11450
rect 5222 11398 5234 11450
rect 5286 11398 5298 11450
rect 5350 11398 5362 11450
rect 5414 11398 5426 11450
rect 5478 11398 13611 11450
rect 13663 11398 13675 11450
rect 13727 11398 13739 11450
rect 13791 11398 13803 11450
rect 13855 11398 13867 11450
rect 13919 11398 22052 11450
rect 22104 11398 22116 11450
rect 22168 11398 22180 11450
rect 22232 11398 22244 11450
rect 22296 11398 22308 11450
rect 22360 11398 30493 11450
rect 30545 11398 30557 11450
rect 30609 11398 30621 11450
rect 30673 11398 30685 11450
rect 30737 11398 30749 11450
rect 30801 11398 34868 11450
rect 1104 11376 34868 11398
rect 1104 10906 35027 10928
rect 1104 10854 9390 10906
rect 9442 10854 9454 10906
rect 9506 10854 9518 10906
rect 9570 10854 9582 10906
rect 9634 10854 9646 10906
rect 9698 10854 17831 10906
rect 17883 10854 17895 10906
rect 17947 10854 17959 10906
rect 18011 10854 18023 10906
rect 18075 10854 18087 10906
rect 18139 10854 26272 10906
rect 26324 10854 26336 10906
rect 26388 10854 26400 10906
rect 26452 10854 26464 10906
rect 26516 10854 26528 10906
rect 26580 10854 34713 10906
rect 34765 10854 34777 10906
rect 34829 10854 34841 10906
rect 34893 10854 34905 10906
rect 34957 10854 34969 10906
rect 35021 10854 35027 10906
rect 1104 10832 35027 10854
rect 1104 10362 34868 10384
rect 1104 10310 5170 10362
rect 5222 10310 5234 10362
rect 5286 10310 5298 10362
rect 5350 10310 5362 10362
rect 5414 10310 5426 10362
rect 5478 10310 13611 10362
rect 13663 10310 13675 10362
rect 13727 10310 13739 10362
rect 13791 10310 13803 10362
rect 13855 10310 13867 10362
rect 13919 10310 22052 10362
rect 22104 10310 22116 10362
rect 22168 10310 22180 10362
rect 22232 10310 22244 10362
rect 22296 10310 22308 10362
rect 22360 10310 30493 10362
rect 30545 10310 30557 10362
rect 30609 10310 30621 10362
rect 30673 10310 30685 10362
rect 30737 10310 30749 10362
rect 30801 10310 34868 10362
rect 1104 10288 34868 10310
rect 1104 9818 35027 9840
rect 1104 9766 9390 9818
rect 9442 9766 9454 9818
rect 9506 9766 9518 9818
rect 9570 9766 9582 9818
rect 9634 9766 9646 9818
rect 9698 9766 17831 9818
rect 17883 9766 17895 9818
rect 17947 9766 17959 9818
rect 18011 9766 18023 9818
rect 18075 9766 18087 9818
rect 18139 9766 26272 9818
rect 26324 9766 26336 9818
rect 26388 9766 26400 9818
rect 26452 9766 26464 9818
rect 26516 9766 26528 9818
rect 26580 9766 34713 9818
rect 34765 9766 34777 9818
rect 34829 9766 34841 9818
rect 34893 9766 34905 9818
rect 34957 9766 34969 9818
rect 35021 9766 35027 9818
rect 1104 9744 35027 9766
rect 1104 9274 34868 9296
rect 1104 9222 5170 9274
rect 5222 9222 5234 9274
rect 5286 9222 5298 9274
rect 5350 9222 5362 9274
rect 5414 9222 5426 9274
rect 5478 9222 13611 9274
rect 13663 9222 13675 9274
rect 13727 9222 13739 9274
rect 13791 9222 13803 9274
rect 13855 9222 13867 9274
rect 13919 9222 22052 9274
rect 22104 9222 22116 9274
rect 22168 9222 22180 9274
rect 22232 9222 22244 9274
rect 22296 9222 22308 9274
rect 22360 9222 30493 9274
rect 30545 9222 30557 9274
rect 30609 9222 30621 9274
rect 30673 9222 30685 9274
rect 30737 9222 30749 9274
rect 30801 9222 34868 9274
rect 1104 9200 34868 9222
rect 1104 8730 35027 8752
rect 1104 8678 9390 8730
rect 9442 8678 9454 8730
rect 9506 8678 9518 8730
rect 9570 8678 9582 8730
rect 9634 8678 9646 8730
rect 9698 8678 17831 8730
rect 17883 8678 17895 8730
rect 17947 8678 17959 8730
rect 18011 8678 18023 8730
rect 18075 8678 18087 8730
rect 18139 8678 26272 8730
rect 26324 8678 26336 8730
rect 26388 8678 26400 8730
rect 26452 8678 26464 8730
rect 26516 8678 26528 8730
rect 26580 8678 34713 8730
rect 34765 8678 34777 8730
rect 34829 8678 34841 8730
rect 34893 8678 34905 8730
rect 34957 8678 34969 8730
rect 35021 8678 35027 8730
rect 1104 8656 35027 8678
rect 1104 8186 34868 8208
rect 1104 8134 5170 8186
rect 5222 8134 5234 8186
rect 5286 8134 5298 8186
rect 5350 8134 5362 8186
rect 5414 8134 5426 8186
rect 5478 8134 13611 8186
rect 13663 8134 13675 8186
rect 13727 8134 13739 8186
rect 13791 8134 13803 8186
rect 13855 8134 13867 8186
rect 13919 8134 22052 8186
rect 22104 8134 22116 8186
rect 22168 8134 22180 8186
rect 22232 8134 22244 8186
rect 22296 8134 22308 8186
rect 22360 8134 30493 8186
rect 30545 8134 30557 8186
rect 30609 8134 30621 8186
rect 30673 8134 30685 8186
rect 30737 8134 30749 8186
rect 30801 8134 34868 8186
rect 1104 8112 34868 8134
rect 1104 7642 35027 7664
rect 1104 7590 9390 7642
rect 9442 7590 9454 7642
rect 9506 7590 9518 7642
rect 9570 7590 9582 7642
rect 9634 7590 9646 7642
rect 9698 7590 17831 7642
rect 17883 7590 17895 7642
rect 17947 7590 17959 7642
rect 18011 7590 18023 7642
rect 18075 7590 18087 7642
rect 18139 7590 26272 7642
rect 26324 7590 26336 7642
rect 26388 7590 26400 7642
rect 26452 7590 26464 7642
rect 26516 7590 26528 7642
rect 26580 7590 34713 7642
rect 34765 7590 34777 7642
rect 34829 7590 34841 7642
rect 34893 7590 34905 7642
rect 34957 7590 34969 7642
rect 35021 7590 35027 7642
rect 1104 7568 35027 7590
rect 1394 7148 1400 7200
rect 1452 7148 1458 7200
rect 1104 7098 34868 7120
rect 1104 7046 5170 7098
rect 5222 7046 5234 7098
rect 5286 7046 5298 7098
rect 5350 7046 5362 7098
rect 5414 7046 5426 7098
rect 5478 7046 13611 7098
rect 13663 7046 13675 7098
rect 13727 7046 13739 7098
rect 13791 7046 13803 7098
rect 13855 7046 13867 7098
rect 13919 7046 22052 7098
rect 22104 7046 22116 7098
rect 22168 7046 22180 7098
rect 22232 7046 22244 7098
rect 22296 7046 22308 7098
rect 22360 7046 30493 7098
rect 30545 7046 30557 7098
rect 30609 7046 30621 7098
rect 30673 7046 30685 7098
rect 30737 7046 30749 7098
rect 30801 7046 34868 7098
rect 1104 7024 34868 7046
rect 1104 6554 35027 6576
rect 1104 6502 9390 6554
rect 9442 6502 9454 6554
rect 9506 6502 9518 6554
rect 9570 6502 9582 6554
rect 9634 6502 9646 6554
rect 9698 6502 17831 6554
rect 17883 6502 17895 6554
rect 17947 6502 17959 6554
rect 18011 6502 18023 6554
rect 18075 6502 18087 6554
rect 18139 6502 26272 6554
rect 26324 6502 26336 6554
rect 26388 6502 26400 6554
rect 26452 6502 26464 6554
rect 26516 6502 26528 6554
rect 26580 6502 34713 6554
rect 34765 6502 34777 6554
rect 34829 6502 34841 6554
rect 34893 6502 34905 6554
rect 34957 6502 34969 6554
rect 35021 6502 35027 6554
rect 1104 6480 35027 6502
rect 1104 6010 34868 6032
rect 1104 5958 5170 6010
rect 5222 5958 5234 6010
rect 5286 5958 5298 6010
rect 5350 5958 5362 6010
rect 5414 5958 5426 6010
rect 5478 5958 13611 6010
rect 13663 5958 13675 6010
rect 13727 5958 13739 6010
rect 13791 5958 13803 6010
rect 13855 5958 13867 6010
rect 13919 5958 22052 6010
rect 22104 5958 22116 6010
rect 22168 5958 22180 6010
rect 22232 5958 22244 6010
rect 22296 5958 22308 6010
rect 22360 5958 30493 6010
rect 30545 5958 30557 6010
rect 30609 5958 30621 6010
rect 30673 5958 30685 6010
rect 30737 5958 30749 6010
rect 30801 5958 34868 6010
rect 1104 5936 34868 5958
rect 34514 5584 34520 5636
rect 34572 5584 34578 5636
rect 1104 5466 35027 5488
rect 1104 5414 9390 5466
rect 9442 5414 9454 5466
rect 9506 5414 9518 5466
rect 9570 5414 9582 5466
rect 9634 5414 9646 5466
rect 9698 5414 17831 5466
rect 17883 5414 17895 5466
rect 17947 5414 17959 5466
rect 18011 5414 18023 5466
rect 18075 5414 18087 5466
rect 18139 5414 26272 5466
rect 26324 5414 26336 5466
rect 26388 5414 26400 5466
rect 26452 5414 26464 5466
rect 26516 5414 26528 5466
rect 26580 5414 34713 5466
rect 34765 5414 34777 5466
rect 34829 5414 34841 5466
rect 34893 5414 34905 5466
rect 34957 5414 34969 5466
rect 35021 5414 35027 5466
rect 1104 5392 35027 5414
rect 1104 4922 34868 4944
rect 1104 4870 5170 4922
rect 5222 4870 5234 4922
rect 5286 4870 5298 4922
rect 5350 4870 5362 4922
rect 5414 4870 5426 4922
rect 5478 4870 13611 4922
rect 13663 4870 13675 4922
rect 13727 4870 13739 4922
rect 13791 4870 13803 4922
rect 13855 4870 13867 4922
rect 13919 4870 22052 4922
rect 22104 4870 22116 4922
rect 22168 4870 22180 4922
rect 22232 4870 22244 4922
rect 22296 4870 22308 4922
rect 22360 4870 30493 4922
rect 30545 4870 30557 4922
rect 30609 4870 30621 4922
rect 30673 4870 30685 4922
rect 30737 4870 30749 4922
rect 30801 4870 34868 4922
rect 1104 4848 34868 4870
rect 1104 4378 35027 4400
rect 1104 4326 9390 4378
rect 9442 4326 9454 4378
rect 9506 4326 9518 4378
rect 9570 4326 9582 4378
rect 9634 4326 9646 4378
rect 9698 4326 17831 4378
rect 17883 4326 17895 4378
rect 17947 4326 17959 4378
rect 18011 4326 18023 4378
rect 18075 4326 18087 4378
rect 18139 4326 26272 4378
rect 26324 4326 26336 4378
rect 26388 4326 26400 4378
rect 26452 4326 26464 4378
rect 26516 4326 26528 4378
rect 26580 4326 34713 4378
rect 34765 4326 34777 4378
rect 34829 4326 34841 4378
rect 34893 4326 34905 4378
rect 34957 4326 34969 4378
rect 35021 4326 35027 4378
rect 1104 4304 35027 4326
rect 1104 3834 34868 3856
rect 1104 3782 5170 3834
rect 5222 3782 5234 3834
rect 5286 3782 5298 3834
rect 5350 3782 5362 3834
rect 5414 3782 5426 3834
rect 5478 3782 13611 3834
rect 13663 3782 13675 3834
rect 13727 3782 13739 3834
rect 13791 3782 13803 3834
rect 13855 3782 13867 3834
rect 13919 3782 22052 3834
rect 22104 3782 22116 3834
rect 22168 3782 22180 3834
rect 22232 3782 22244 3834
rect 22296 3782 22308 3834
rect 22360 3782 30493 3834
rect 30545 3782 30557 3834
rect 30609 3782 30621 3834
rect 30673 3782 30685 3834
rect 30737 3782 30749 3834
rect 30801 3782 34868 3834
rect 1104 3760 34868 3782
rect 1104 3290 35027 3312
rect 1104 3238 9390 3290
rect 9442 3238 9454 3290
rect 9506 3238 9518 3290
rect 9570 3238 9582 3290
rect 9634 3238 9646 3290
rect 9698 3238 17831 3290
rect 17883 3238 17895 3290
rect 17947 3238 17959 3290
rect 18011 3238 18023 3290
rect 18075 3238 18087 3290
rect 18139 3238 26272 3290
rect 26324 3238 26336 3290
rect 26388 3238 26400 3290
rect 26452 3238 26464 3290
rect 26516 3238 26528 3290
rect 26580 3238 34713 3290
rect 34765 3238 34777 3290
rect 34829 3238 34841 3290
rect 34893 3238 34905 3290
rect 34957 3238 34969 3290
rect 35021 3238 35027 3290
rect 1104 3216 35027 3238
rect 1104 2746 34868 2768
rect 1104 2694 5170 2746
rect 5222 2694 5234 2746
rect 5286 2694 5298 2746
rect 5350 2694 5362 2746
rect 5414 2694 5426 2746
rect 5478 2694 13611 2746
rect 13663 2694 13675 2746
rect 13727 2694 13739 2746
rect 13791 2694 13803 2746
rect 13855 2694 13867 2746
rect 13919 2694 22052 2746
rect 22104 2694 22116 2746
rect 22168 2694 22180 2746
rect 22232 2694 22244 2746
rect 22296 2694 22308 2746
rect 22360 2694 30493 2746
rect 30545 2694 30557 2746
rect 30609 2694 30621 2746
rect 30673 2694 30685 2746
rect 30737 2694 30749 2746
rect 30801 2694 34868 2746
rect 1104 2672 34868 2694
rect 20714 2456 20720 2508
rect 20772 2456 20778 2508
rect 13630 2388 13636 2440
rect 13688 2388 13694 2440
rect 20254 2388 20260 2440
rect 20312 2388 20318 2440
rect 14 2252 20 2304
rect 72 2292 78 2304
rect 1397 2295 1455 2301
rect 1397 2292 1409 2295
rect 72 2264 1409 2292
rect 72 2252 78 2264
rect 1397 2261 1409 2264
rect 1443 2261 1455 2295
rect 1397 2255 1455 2261
rect 6546 2252 6552 2304
rect 6604 2252 6610 2304
rect 27154 2252 27160 2304
rect 27212 2252 27218 2304
rect 34238 2252 34244 2304
rect 34296 2252 34302 2304
rect 1104 2202 35027 2224
rect 1104 2150 9390 2202
rect 9442 2150 9454 2202
rect 9506 2150 9518 2202
rect 9570 2150 9582 2202
rect 9634 2150 9646 2202
rect 9698 2150 17831 2202
rect 17883 2150 17895 2202
rect 17947 2150 17959 2202
rect 18011 2150 18023 2202
rect 18075 2150 18087 2202
rect 18139 2150 26272 2202
rect 26324 2150 26336 2202
rect 26388 2150 26400 2202
rect 26452 2150 26464 2202
rect 26516 2150 26528 2202
rect 26580 2150 34713 2202
rect 34765 2150 34777 2202
rect 34829 2150 34841 2202
rect 34893 2150 34905 2202
rect 34957 2150 34969 2202
rect 35021 2150 35027 2202
rect 1104 2128 35027 2150
<< via1 >>
rect 5170 39686 5222 39738
rect 5234 39686 5286 39738
rect 5298 39686 5350 39738
rect 5362 39686 5414 39738
rect 5426 39686 5478 39738
rect 13611 39686 13663 39738
rect 13675 39686 13727 39738
rect 13739 39686 13791 39738
rect 13803 39686 13855 39738
rect 13867 39686 13919 39738
rect 22052 39686 22104 39738
rect 22116 39686 22168 39738
rect 22180 39686 22232 39738
rect 22244 39686 22296 39738
rect 22308 39686 22360 39738
rect 30493 39686 30545 39738
rect 30557 39686 30609 39738
rect 30621 39686 30673 39738
rect 30685 39686 30737 39738
rect 30749 39686 30801 39738
rect 18328 39584 18380 39636
rect 3056 39423 3108 39432
rect 3056 39389 3065 39423
rect 3065 39389 3099 39423
rect 3099 39389 3108 39423
rect 3056 39380 3108 39389
rect 8392 39380 8444 39432
rect 14832 39380 14884 39432
rect 16396 39491 16448 39500
rect 16396 39457 16405 39491
rect 16405 39457 16439 39491
rect 16439 39457 16448 39491
rect 16396 39448 16448 39457
rect 4896 39244 4948 39296
rect 8484 39287 8536 39296
rect 8484 39253 8493 39287
rect 8493 39253 8527 39287
rect 8527 39253 8536 39287
rect 8484 39244 8536 39253
rect 13912 39244 13964 39296
rect 17500 39423 17552 39432
rect 17500 39389 17509 39423
rect 17509 39389 17543 39423
rect 17543 39389 17552 39423
rect 17500 39380 17552 39389
rect 17592 39423 17644 39432
rect 17592 39389 17601 39423
rect 17601 39389 17635 39423
rect 17635 39389 17644 39423
rect 17592 39380 17644 39389
rect 16120 39312 16172 39364
rect 18236 39423 18288 39432
rect 18236 39389 18245 39423
rect 18245 39389 18279 39423
rect 18279 39389 18288 39423
rect 18236 39380 18288 39389
rect 22836 39516 22888 39568
rect 21916 39448 21968 39500
rect 35440 39448 35492 39500
rect 19156 39312 19208 39364
rect 23112 39380 23164 39432
rect 22744 39312 22796 39364
rect 15292 39287 15344 39296
rect 15292 39253 15301 39287
rect 15301 39253 15335 39287
rect 15335 39253 15344 39287
rect 15292 39244 15344 39253
rect 15384 39244 15436 39296
rect 17040 39287 17092 39296
rect 17040 39253 17049 39287
rect 17049 39253 17083 39287
rect 17083 39253 17092 39287
rect 17040 39244 17092 39253
rect 17316 39287 17368 39296
rect 17316 39253 17325 39287
rect 17325 39253 17359 39287
rect 17359 39253 17368 39287
rect 17316 39244 17368 39253
rect 20536 39287 20588 39296
rect 20536 39253 20545 39287
rect 20545 39253 20579 39287
rect 20579 39253 20588 39287
rect 20536 39244 20588 39253
rect 21456 39287 21508 39296
rect 21456 39253 21465 39287
rect 21465 39253 21499 39287
rect 21499 39253 21508 39287
rect 21456 39244 21508 39253
rect 9390 39142 9442 39194
rect 9454 39142 9506 39194
rect 9518 39142 9570 39194
rect 9582 39142 9634 39194
rect 9646 39142 9698 39194
rect 17831 39142 17883 39194
rect 17895 39142 17947 39194
rect 17959 39142 18011 39194
rect 18023 39142 18075 39194
rect 18087 39142 18139 39194
rect 26272 39142 26324 39194
rect 26336 39142 26388 39194
rect 26400 39142 26452 39194
rect 26464 39142 26516 39194
rect 26528 39142 26580 39194
rect 34713 39142 34765 39194
rect 34777 39142 34829 39194
rect 34841 39142 34893 39194
rect 34905 39142 34957 39194
rect 34969 39142 35021 39194
rect 3056 39040 3108 39092
rect 13912 39040 13964 39092
rect 1308 38904 1360 38956
rect 16396 39040 16448 39092
rect 17040 39040 17092 39092
rect 20536 39040 20588 39092
rect 21456 39040 21508 39092
rect 21640 39040 21692 39092
rect 15384 38904 15436 38956
rect 14096 38879 14148 38888
rect 14096 38845 14105 38879
rect 14105 38845 14139 38879
rect 14139 38845 14148 38879
rect 14096 38836 14148 38845
rect 16120 38836 16172 38888
rect 19340 38836 19392 38888
rect 23204 38879 23256 38888
rect 23204 38845 23213 38879
rect 23213 38845 23247 38879
rect 23247 38845 23256 38879
rect 23204 38836 23256 38845
rect 15752 38743 15804 38752
rect 15752 38709 15761 38743
rect 15761 38709 15795 38743
rect 15795 38709 15804 38743
rect 15752 38700 15804 38709
rect 17040 38700 17092 38752
rect 18512 38743 18564 38752
rect 18512 38709 18521 38743
rect 18521 38709 18555 38743
rect 18555 38709 18564 38743
rect 18512 38700 18564 38709
rect 21824 38743 21876 38752
rect 21824 38709 21833 38743
rect 21833 38709 21867 38743
rect 21867 38709 21876 38743
rect 21824 38700 21876 38709
rect 23940 38743 23992 38752
rect 23940 38709 23949 38743
rect 23949 38709 23983 38743
rect 23983 38709 23992 38743
rect 23940 38700 23992 38709
rect 5170 38598 5222 38650
rect 5234 38598 5286 38650
rect 5298 38598 5350 38650
rect 5362 38598 5414 38650
rect 5426 38598 5478 38650
rect 13611 38598 13663 38650
rect 13675 38598 13727 38650
rect 13739 38598 13791 38650
rect 13803 38598 13855 38650
rect 13867 38598 13919 38650
rect 22052 38598 22104 38650
rect 22116 38598 22168 38650
rect 22180 38598 22232 38650
rect 22244 38598 22296 38650
rect 22308 38598 22360 38650
rect 30493 38598 30545 38650
rect 30557 38598 30609 38650
rect 30621 38598 30673 38650
rect 30685 38598 30737 38650
rect 30749 38598 30801 38650
rect 4896 38335 4948 38344
rect 4896 38301 4905 38335
rect 4905 38301 4939 38335
rect 4939 38301 4948 38335
rect 4896 38292 4948 38301
rect 7472 38292 7524 38344
rect 8392 38335 8444 38344
rect 8392 38301 8401 38335
rect 8401 38301 8435 38335
rect 8435 38301 8444 38335
rect 8392 38292 8444 38301
rect 8484 38335 8536 38344
rect 8484 38301 8493 38335
rect 8493 38301 8527 38335
rect 8527 38301 8536 38335
rect 8484 38292 8536 38301
rect 15292 38496 15344 38548
rect 18236 38496 18288 38548
rect 22744 38539 22796 38548
rect 22744 38505 22753 38539
rect 22753 38505 22787 38539
rect 22787 38505 22796 38539
rect 22744 38496 22796 38505
rect 22836 38496 22888 38548
rect 14096 38292 14148 38344
rect 15752 38292 15804 38344
rect 18512 38360 18564 38412
rect 21272 38403 21324 38412
rect 21272 38369 21281 38403
rect 21281 38369 21315 38403
rect 21315 38369 21324 38403
rect 21272 38360 21324 38369
rect 21824 38360 21876 38412
rect 23940 38360 23992 38412
rect 17040 38292 17092 38344
rect 17592 38335 17644 38344
rect 17592 38301 17601 38335
rect 17601 38301 17635 38335
rect 17635 38301 17644 38335
rect 17592 38292 17644 38301
rect 18236 38292 18288 38344
rect 19340 38292 19392 38344
rect 6920 38156 6972 38208
rect 8668 38199 8720 38208
rect 8668 38165 8677 38199
rect 8677 38165 8711 38199
rect 8711 38165 8720 38199
rect 8668 38156 8720 38165
rect 15568 38199 15620 38208
rect 15568 38165 15577 38199
rect 15577 38165 15611 38199
rect 15611 38165 15620 38199
rect 15568 38156 15620 38165
rect 20720 38224 20772 38276
rect 18420 38199 18472 38208
rect 18420 38165 18429 38199
rect 18429 38165 18463 38199
rect 18463 38165 18472 38199
rect 18420 38156 18472 38165
rect 22560 38156 22612 38208
rect 22652 38199 22704 38208
rect 22652 38165 22661 38199
rect 22661 38165 22695 38199
rect 22695 38165 22704 38199
rect 22652 38156 22704 38165
rect 9390 38054 9442 38106
rect 9454 38054 9506 38106
rect 9518 38054 9570 38106
rect 9582 38054 9634 38106
rect 9646 38054 9698 38106
rect 17831 38054 17883 38106
rect 17895 38054 17947 38106
rect 17959 38054 18011 38106
rect 18023 38054 18075 38106
rect 18087 38054 18139 38106
rect 26272 38054 26324 38106
rect 26336 38054 26388 38106
rect 26400 38054 26452 38106
rect 26464 38054 26516 38106
rect 26528 38054 26580 38106
rect 34713 38054 34765 38106
rect 34777 38054 34829 38106
rect 34841 38054 34893 38106
rect 34905 38054 34957 38106
rect 34969 38054 35021 38106
rect 8668 37952 8720 38004
rect 17684 37995 17736 38004
rect 17684 37961 17693 37995
rect 17693 37961 17727 37995
rect 17727 37961 17736 37995
rect 17684 37952 17736 37961
rect 20720 37995 20772 38004
rect 20720 37961 20729 37995
rect 20729 37961 20763 37995
rect 20763 37961 20772 37995
rect 20720 37952 20772 37961
rect 21272 37952 21324 38004
rect 21548 37952 21600 38004
rect 21916 37952 21968 38004
rect 6000 37748 6052 37800
rect 8392 37748 8444 37800
rect 10508 37816 10560 37868
rect 10692 37859 10744 37868
rect 10692 37825 10701 37859
rect 10701 37825 10735 37859
rect 10735 37825 10744 37859
rect 10692 37816 10744 37825
rect 10784 37816 10836 37868
rect 11152 37859 11204 37868
rect 11152 37825 11161 37859
rect 11161 37825 11195 37859
rect 11195 37825 11204 37859
rect 11152 37816 11204 37825
rect 11704 37859 11756 37868
rect 11704 37825 11713 37859
rect 11713 37825 11747 37859
rect 11747 37825 11756 37859
rect 11704 37816 11756 37825
rect 14004 37816 14056 37868
rect 14464 37859 14516 37868
rect 14464 37825 14473 37859
rect 14473 37825 14507 37859
rect 14507 37825 14516 37859
rect 14464 37816 14516 37825
rect 15384 37884 15436 37936
rect 18052 37884 18104 37936
rect 19156 37884 19208 37936
rect 19248 37884 19300 37936
rect 17592 37816 17644 37868
rect 18512 37816 18564 37868
rect 18604 37816 18656 37868
rect 11060 37791 11112 37800
rect 11060 37757 11069 37791
rect 11069 37757 11103 37791
rect 11103 37757 11112 37791
rect 11060 37748 11112 37757
rect 11980 37748 12032 37800
rect 14096 37748 14148 37800
rect 17408 37791 17460 37800
rect 17408 37757 17417 37791
rect 17417 37757 17451 37791
rect 17451 37757 17460 37791
rect 17408 37748 17460 37757
rect 17868 37791 17920 37800
rect 17868 37757 17877 37791
rect 17877 37757 17911 37791
rect 17911 37757 17920 37791
rect 17868 37748 17920 37757
rect 19340 37791 19392 37800
rect 19340 37757 19349 37791
rect 19349 37757 19383 37791
rect 19383 37757 19392 37791
rect 19340 37748 19392 37757
rect 20536 37816 20588 37868
rect 21548 37816 21600 37868
rect 21640 37859 21692 37868
rect 21640 37825 21649 37859
rect 21649 37825 21683 37859
rect 21683 37825 21692 37859
rect 21640 37816 21692 37825
rect 12992 37680 13044 37732
rect 16120 37723 16172 37732
rect 16120 37689 16129 37723
rect 16129 37689 16163 37723
rect 16163 37689 16172 37723
rect 16120 37680 16172 37689
rect 7288 37612 7340 37664
rect 9036 37655 9088 37664
rect 9036 37621 9045 37655
rect 9045 37621 9079 37655
rect 9079 37621 9088 37655
rect 9036 37612 9088 37621
rect 10140 37655 10192 37664
rect 10140 37621 10149 37655
rect 10149 37621 10183 37655
rect 10183 37621 10192 37655
rect 10140 37612 10192 37621
rect 10876 37655 10928 37664
rect 10876 37621 10885 37655
rect 10885 37621 10919 37655
rect 10919 37621 10928 37655
rect 10876 37612 10928 37621
rect 11520 37655 11572 37664
rect 11520 37621 11529 37655
rect 11529 37621 11563 37655
rect 11563 37621 11572 37655
rect 11520 37612 11572 37621
rect 12624 37612 12676 37664
rect 12900 37655 12952 37664
rect 12900 37621 12909 37655
rect 12909 37621 12943 37655
rect 12943 37621 12952 37655
rect 12900 37612 12952 37621
rect 17224 37655 17276 37664
rect 17224 37621 17233 37655
rect 17233 37621 17267 37655
rect 17267 37621 17276 37655
rect 17224 37612 17276 37621
rect 17500 37680 17552 37732
rect 17776 37680 17828 37732
rect 23388 37748 23440 37800
rect 18144 37612 18196 37664
rect 19432 37655 19484 37664
rect 19432 37621 19441 37655
rect 19441 37621 19475 37655
rect 19475 37621 19484 37655
rect 19432 37612 19484 37621
rect 21180 37655 21232 37664
rect 21180 37621 21189 37655
rect 21189 37621 21223 37655
rect 21223 37621 21232 37655
rect 21180 37612 21232 37621
rect 22376 37655 22428 37664
rect 22376 37621 22385 37655
rect 22385 37621 22419 37655
rect 22419 37621 22428 37655
rect 22376 37612 22428 37621
rect 5170 37510 5222 37562
rect 5234 37510 5286 37562
rect 5298 37510 5350 37562
rect 5362 37510 5414 37562
rect 5426 37510 5478 37562
rect 13611 37510 13663 37562
rect 13675 37510 13727 37562
rect 13739 37510 13791 37562
rect 13803 37510 13855 37562
rect 13867 37510 13919 37562
rect 22052 37510 22104 37562
rect 22116 37510 22168 37562
rect 22180 37510 22232 37562
rect 22244 37510 22296 37562
rect 22308 37510 22360 37562
rect 30493 37510 30545 37562
rect 30557 37510 30609 37562
rect 30621 37510 30673 37562
rect 30685 37510 30737 37562
rect 30749 37510 30801 37562
rect 11060 37408 11112 37460
rect 14004 37408 14056 37460
rect 14464 37408 14516 37460
rect 17316 37451 17368 37460
rect 17316 37417 17325 37451
rect 17325 37417 17359 37451
rect 17359 37417 17368 37451
rect 17316 37408 17368 37417
rect 17684 37408 17736 37460
rect 17868 37408 17920 37460
rect 19248 37408 19300 37460
rect 21180 37408 21232 37460
rect 22468 37408 22520 37460
rect 22652 37408 22704 37460
rect 15568 37340 15620 37392
rect 17776 37383 17828 37392
rect 7288 37315 7340 37324
rect 7288 37281 7297 37315
rect 7297 37281 7331 37315
rect 7331 37281 7340 37315
rect 7288 37272 7340 37281
rect 17776 37349 17785 37383
rect 17785 37349 17819 37383
rect 17819 37349 17828 37383
rect 17776 37340 17828 37349
rect 18052 37272 18104 37324
rect 8024 37136 8076 37188
rect 8852 37204 8904 37256
rect 14096 37204 14148 37256
rect 10140 37136 10192 37188
rect 11520 37136 11572 37188
rect 12900 37136 12952 37188
rect 13084 37136 13136 37188
rect 14372 37247 14424 37256
rect 14372 37213 14381 37247
rect 14381 37213 14415 37247
rect 14415 37213 14424 37247
rect 14372 37204 14424 37213
rect 17316 37204 17368 37256
rect 17592 37204 17644 37256
rect 18144 37247 18196 37256
rect 18144 37213 18153 37247
rect 18153 37213 18187 37247
rect 18187 37213 18196 37247
rect 18144 37204 18196 37213
rect 18236 37136 18288 37188
rect 9128 37068 9180 37120
rect 12440 37111 12492 37120
rect 12440 37077 12449 37111
rect 12449 37077 12483 37111
rect 12483 37077 12492 37111
rect 12440 37068 12492 37077
rect 13268 37068 13320 37120
rect 15384 37068 15436 37120
rect 16304 37068 16356 37120
rect 16948 37111 17000 37120
rect 16948 37077 16957 37111
rect 16957 37077 16991 37111
rect 16991 37077 17000 37111
rect 16948 37068 17000 37077
rect 17040 37068 17092 37120
rect 17684 37068 17736 37120
rect 18328 37068 18380 37120
rect 19340 37204 19392 37256
rect 20628 37247 20680 37256
rect 20628 37213 20637 37247
rect 20637 37213 20671 37247
rect 20671 37213 20680 37247
rect 20628 37204 20680 37213
rect 20720 37247 20772 37256
rect 20720 37213 20729 37247
rect 20729 37213 20763 37247
rect 20763 37213 20772 37247
rect 20720 37204 20772 37213
rect 19064 37136 19116 37188
rect 20536 37136 20588 37188
rect 21916 37204 21968 37256
rect 22560 37247 22612 37256
rect 22560 37213 22569 37247
rect 22569 37213 22603 37247
rect 22603 37213 22612 37247
rect 22560 37204 22612 37213
rect 21088 37111 21140 37120
rect 21088 37077 21097 37111
rect 21097 37077 21131 37111
rect 21131 37077 21140 37111
rect 21088 37068 21140 37077
rect 21640 37111 21692 37120
rect 21640 37077 21649 37111
rect 21649 37077 21683 37111
rect 21683 37077 21692 37111
rect 21640 37068 21692 37077
rect 23020 37111 23072 37120
rect 23020 37077 23029 37111
rect 23029 37077 23063 37111
rect 23063 37077 23072 37111
rect 23020 37068 23072 37077
rect 9390 36966 9442 37018
rect 9454 36966 9506 37018
rect 9518 36966 9570 37018
rect 9582 36966 9634 37018
rect 9646 36966 9698 37018
rect 17831 36966 17883 37018
rect 17895 36966 17947 37018
rect 17959 36966 18011 37018
rect 18023 36966 18075 37018
rect 18087 36966 18139 37018
rect 26272 36966 26324 37018
rect 26336 36966 26388 37018
rect 26400 36966 26452 37018
rect 26464 36966 26516 37018
rect 26528 36966 26580 37018
rect 34713 36966 34765 37018
rect 34777 36966 34829 37018
rect 34841 36966 34893 37018
rect 34905 36966 34957 37018
rect 34969 36966 35021 37018
rect 8024 36907 8076 36916
rect 8024 36873 8033 36907
rect 8033 36873 8067 36907
rect 8067 36873 8076 36907
rect 8024 36864 8076 36873
rect 12440 36864 12492 36916
rect 13268 36864 13320 36916
rect 14372 36864 14424 36916
rect 9036 36839 9088 36848
rect 9036 36805 9070 36839
rect 9070 36805 9088 36839
rect 9036 36796 9088 36805
rect 7472 36771 7524 36780
rect 7472 36737 7481 36771
rect 7481 36737 7515 36771
rect 7515 36737 7524 36771
rect 7472 36728 7524 36737
rect 8852 36728 8904 36780
rect 10048 36728 10100 36780
rect 12900 36771 12952 36780
rect 12900 36737 12909 36771
rect 12909 36737 12943 36771
rect 12943 36737 12952 36771
rect 12900 36728 12952 36737
rect 17040 36796 17092 36848
rect 17316 36864 17368 36916
rect 20536 36864 20588 36916
rect 21640 36864 21692 36916
rect 21916 36907 21968 36916
rect 21916 36873 21925 36907
rect 21925 36873 21959 36907
rect 21959 36873 21968 36907
rect 21916 36864 21968 36873
rect 23388 36907 23440 36916
rect 23388 36873 23397 36907
rect 23397 36873 23431 36907
rect 23431 36873 23440 36907
rect 23388 36864 23440 36873
rect 8576 36703 8628 36712
rect 8576 36669 8585 36703
rect 8585 36669 8619 36703
rect 8619 36669 8628 36703
rect 8576 36660 8628 36669
rect 10600 36703 10652 36712
rect 10600 36669 10609 36703
rect 10609 36669 10643 36703
rect 10643 36669 10652 36703
rect 10600 36660 10652 36669
rect 10876 36660 10928 36712
rect 12532 36703 12584 36712
rect 12532 36669 12541 36703
rect 12541 36669 12575 36703
rect 12575 36669 12584 36703
rect 12532 36660 12584 36669
rect 12716 36660 12768 36712
rect 13452 36660 13504 36712
rect 15936 36703 15988 36712
rect 15936 36669 15945 36703
rect 15945 36669 15979 36703
rect 15979 36669 15988 36703
rect 15936 36660 15988 36669
rect 7656 36567 7708 36576
rect 7656 36533 7665 36567
rect 7665 36533 7699 36567
rect 7699 36533 7708 36567
rect 7656 36524 7708 36533
rect 10232 36567 10284 36576
rect 10232 36533 10241 36567
rect 10241 36533 10275 36567
rect 10275 36533 10284 36567
rect 10232 36524 10284 36533
rect 11244 36524 11296 36576
rect 12440 36524 12492 36576
rect 13176 36567 13228 36576
rect 13176 36533 13185 36567
rect 13185 36533 13219 36567
rect 13219 36533 13228 36567
rect 13176 36524 13228 36533
rect 13360 36524 13412 36576
rect 14648 36567 14700 36576
rect 14648 36533 14657 36567
rect 14657 36533 14691 36567
rect 14691 36533 14700 36567
rect 14648 36524 14700 36533
rect 17684 36796 17736 36848
rect 19340 36796 19392 36848
rect 18604 36728 18656 36780
rect 19984 36771 20036 36780
rect 19984 36737 19993 36771
rect 19993 36737 20027 36771
rect 20027 36737 20036 36771
rect 19984 36728 20036 36737
rect 23020 36839 23072 36848
rect 23020 36805 23038 36839
rect 23038 36805 23072 36839
rect 23020 36796 23072 36805
rect 23204 36728 23256 36780
rect 24492 36771 24544 36780
rect 24492 36737 24510 36771
rect 24510 36737 24544 36771
rect 24492 36728 24544 36737
rect 19432 36660 19484 36712
rect 20536 36703 20588 36712
rect 20536 36669 20545 36703
rect 20545 36669 20579 36703
rect 20579 36669 20588 36703
rect 20536 36660 20588 36669
rect 20076 36567 20128 36576
rect 20076 36533 20085 36567
rect 20085 36533 20119 36567
rect 20119 36533 20128 36567
rect 20076 36524 20128 36533
rect 20720 36524 20772 36576
rect 5170 36422 5222 36474
rect 5234 36422 5286 36474
rect 5298 36422 5350 36474
rect 5362 36422 5414 36474
rect 5426 36422 5478 36474
rect 13611 36422 13663 36474
rect 13675 36422 13727 36474
rect 13739 36422 13791 36474
rect 13803 36422 13855 36474
rect 13867 36422 13919 36474
rect 22052 36422 22104 36474
rect 22116 36422 22168 36474
rect 22180 36422 22232 36474
rect 22244 36422 22296 36474
rect 22308 36422 22360 36474
rect 30493 36422 30545 36474
rect 30557 36422 30609 36474
rect 30621 36422 30673 36474
rect 30685 36422 30737 36474
rect 30749 36422 30801 36474
rect 8576 36320 8628 36372
rect 9128 36320 9180 36372
rect 10232 36320 10284 36372
rect 10600 36320 10652 36372
rect 11704 36320 11756 36372
rect 12532 36320 12584 36372
rect 12900 36320 12952 36372
rect 12992 36320 13044 36372
rect 13268 36320 13320 36372
rect 13360 36320 13412 36372
rect 940 36116 992 36168
rect 6920 36116 6972 36168
rect 10784 36227 10836 36236
rect 10784 36193 10793 36227
rect 10793 36193 10827 36227
rect 10827 36193 10836 36227
rect 10784 36184 10836 36193
rect 11152 36184 11204 36236
rect 12624 36184 12676 36236
rect 10692 36048 10744 36100
rect 10876 36116 10928 36168
rect 11980 36159 12032 36168
rect 11980 36125 11989 36159
rect 11989 36125 12023 36159
rect 12023 36125 12032 36159
rect 11980 36116 12032 36125
rect 15936 36320 15988 36372
rect 15476 36295 15528 36304
rect 15476 36261 15485 36295
rect 15485 36261 15519 36295
rect 15519 36261 15528 36295
rect 15476 36252 15528 36261
rect 16764 36184 16816 36236
rect 12716 36048 12768 36100
rect 14096 36159 14148 36168
rect 14096 36125 14105 36159
rect 14105 36125 14139 36159
rect 14139 36125 14148 36159
rect 14096 36116 14148 36125
rect 14648 36116 14700 36168
rect 9772 36023 9824 36032
rect 9772 35989 9781 36023
rect 9781 35989 9815 36023
rect 9815 35989 9824 36023
rect 9772 35980 9824 35989
rect 9956 36023 10008 36032
rect 9956 35989 9965 36023
rect 9965 35989 9999 36023
rect 9999 35989 10008 36023
rect 9956 35980 10008 35989
rect 12532 35980 12584 36032
rect 13084 35980 13136 36032
rect 13636 36023 13688 36032
rect 13636 35989 13645 36023
rect 13645 35989 13679 36023
rect 13679 35989 13688 36023
rect 13636 35980 13688 35989
rect 14556 35980 14608 36032
rect 16212 36023 16264 36032
rect 16212 35989 16221 36023
rect 16221 35989 16255 36023
rect 16255 35989 16264 36023
rect 16212 35980 16264 35989
rect 16948 36184 17000 36236
rect 19064 36363 19116 36372
rect 19064 36329 19073 36363
rect 19073 36329 19107 36363
rect 19107 36329 19116 36363
rect 19064 36320 19116 36329
rect 17316 36252 17368 36304
rect 20444 36252 20496 36304
rect 17224 36159 17276 36168
rect 17224 36125 17233 36159
rect 17233 36125 17267 36159
rect 17267 36125 17276 36159
rect 17224 36116 17276 36125
rect 17500 36116 17552 36168
rect 17868 36184 17920 36236
rect 18604 36184 18656 36236
rect 19156 36184 19208 36236
rect 20628 36184 20680 36236
rect 20812 36227 20864 36236
rect 20812 36193 20821 36227
rect 20821 36193 20855 36227
rect 20855 36193 20864 36227
rect 20812 36184 20864 36193
rect 18696 36159 18748 36168
rect 18696 36125 18705 36159
rect 18705 36125 18739 36159
rect 18739 36125 18748 36159
rect 18696 36116 18748 36125
rect 16488 35980 16540 36032
rect 16672 36023 16724 36032
rect 16672 35989 16681 36023
rect 16681 35989 16715 36023
rect 16715 35989 16724 36023
rect 16672 35980 16724 35989
rect 17868 36048 17920 36100
rect 19892 36159 19944 36168
rect 19892 36125 19901 36159
rect 19901 36125 19935 36159
rect 19935 36125 19944 36159
rect 19892 36116 19944 36125
rect 18420 35980 18472 36032
rect 20168 35980 20220 36032
rect 20720 36116 20772 36168
rect 23204 36116 23256 36168
rect 20904 35980 20956 36032
rect 21364 36048 21416 36100
rect 23848 36048 23900 36100
rect 21824 35980 21876 36032
rect 22192 36023 22244 36032
rect 22192 35989 22201 36023
rect 22201 35989 22235 36023
rect 22235 35989 22244 36023
rect 22192 35980 22244 35989
rect 22284 35980 22336 36032
rect 9390 35878 9442 35930
rect 9454 35878 9506 35930
rect 9518 35878 9570 35930
rect 9582 35878 9634 35930
rect 9646 35878 9698 35930
rect 17831 35878 17883 35930
rect 17895 35878 17947 35930
rect 17959 35878 18011 35930
rect 18023 35878 18075 35930
rect 18087 35878 18139 35930
rect 26272 35878 26324 35930
rect 26336 35878 26388 35930
rect 26400 35878 26452 35930
rect 26464 35878 26516 35930
rect 26528 35878 26580 35930
rect 34713 35878 34765 35930
rect 34777 35878 34829 35930
rect 34841 35878 34893 35930
rect 34905 35878 34957 35930
rect 34969 35878 35021 35930
rect 8760 35683 8812 35692
rect 8760 35649 8769 35683
rect 8769 35649 8803 35683
rect 8803 35649 8812 35683
rect 8760 35640 8812 35649
rect 8852 35640 8904 35692
rect 9772 35776 9824 35828
rect 11152 35776 11204 35828
rect 11796 35776 11848 35828
rect 11888 35683 11940 35692
rect 9312 35572 9364 35624
rect 11888 35649 11897 35683
rect 11897 35649 11931 35683
rect 11931 35649 11940 35683
rect 11888 35640 11940 35649
rect 12532 35776 12584 35828
rect 13176 35776 13228 35828
rect 13452 35776 13504 35828
rect 13636 35776 13688 35828
rect 16672 35776 16724 35828
rect 18696 35776 18748 35828
rect 20444 35776 20496 35828
rect 20536 35819 20588 35828
rect 20536 35785 20545 35819
rect 20545 35785 20579 35819
rect 20579 35785 20588 35819
rect 20536 35776 20588 35785
rect 21088 35776 21140 35828
rect 21364 35819 21416 35828
rect 21364 35785 21373 35819
rect 21373 35785 21407 35819
rect 21407 35785 21416 35819
rect 21364 35776 21416 35785
rect 21824 35819 21876 35828
rect 21824 35785 21833 35819
rect 21833 35785 21867 35819
rect 21867 35785 21876 35819
rect 21824 35776 21876 35785
rect 22468 35776 22520 35828
rect 23848 35819 23900 35828
rect 23848 35785 23857 35819
rect 23857 35785 23891 35819
rect 23891 35785 23900 35819
rect 23848 35776 23900 35785
rect 24492 35776 24544 35828
rect 12440 35572 12492 35624
rect 12992 35683 13044 35692
rect 12992 35649 13001 35683
rect 13001 35649 13035 35683
rect 13035 35649 13044 35683
rect 12992 35640 13044 35649
rect 14096 35640 14148 35692
rect 13360 35572 13412 35624
rect 16028 35640 16080 35692
rect 11612 35504 11664 35556
rect 13084 35504 13136 35556
rect 14556 35504 14608 35556
rect 16764 35751 16816 35760
rect 16764 35717 16773 35751
rect 16773 35717 16807 35751
rect 16807 35717 16816 35751
rect 16764 35708 16816 35717
rect 17316 35708 17368 35760
rect 18972 35708 19024 35760
rect 17684 35683 17736 35692
rect 17684 35649 17693 35683
rect 17693 35649 17727 35683
rect 17727 35649 17736 35683
rect 17684 35640 17736 35649
rect 20076 35708 20128 35760
rect 16304 35504 16356 35556
rect 22284 35640 22336 35692
rect 22468 35640 22520 35692
rect 21916 35572 21968 35624
rect 22192 35504 22244 35556
rect 22560 35504 22612 35556
rect 11704 35436 11756 35488
rect 12992 35436 13044 35488
rect 14740 35479 14792 35488
rect 14740 35445 14749 35479
rect 14749 35445 14783 35479
rect 14783 35445 14792 35479
rect 14740 35436 14792 35445
rect 16120 35436 16172 35488
rect 17224 35479 17276 35488
rect 17224 35445 17233 35479
rect 17233 35445 17267 35479
rect 17267 35445 17276 35479
rect 17224 35436 17276 35445
rect 21272 35479 21324 35488
rect 21272 35445 21281 35479
rect 21281 35445 21315 35479
rect 21315 35445 21324 35479
rect 21272 35436 21324 35445
rect 21824 35436 21876 35488
rect 22652 35436 22704 35488
rect 24124 35683 24176 35692
rect 24124 35649 24133 35683
rect 24133 35649 24167 35683
rect 24167 35649 24176 35683
rect 24124 35640 24176 35649
rect 5170 35334 5222 35386
rect 5234 35334 5286 35386
rect 5298 35334 5350 35386
rect 5362 35334 5414 35386
rect 5426 35334 5478 35386
rect 13611 35334 13663 35386
rect 13675 35334 13727 35386
rect 13739 35334 13791 35386
rect 13803 35334 13855 35386
rect 13867 35334 13919 35386
rect 22052 35334 22104 35386
rect 22116 35334 22168 35386
rect 22180 35334 22232 35386
rect 22244 35334 22296 35386
rect 22308 35334 22360 35386
rect 30493 35334 30545 35386
rect 30557 35334 30609 35386
rect 30621 35334 30673 35386
rect 30685 35334 30737 35386
rect 30749 35334 30801 35386
rect 8760 35232 8812 35284
rect 10784 35207 10836 35216
rect 10784 35173 10793 35207
rect 10793 35173 10827 35207
rect 10827 35173 10836 35207
rect 10784 35164 10836 35173
rect 9312 35096 9364 35148
rect 12900 35096 12952 35148
rect 9956 35028 10008 35080
rect 10048 34960 10100 35012
rect 11244 35071 11296 35080
rect 11244 35037 11253 35071
rect 11253 35037 11287 35071
rect 11287 35037 11296 35071
rect 11244 35028 11296 35037
rect 11336 35071 11388 35080
rect 11336 35037 11345 35071
rect 11345 35037 11379 35071
rect 11379 35037 11388 35071
rect 11336 35028 11388 35037
rect 11520 35028 11572 35080
rect 11612 35071 11664 35080
rect 11612 35037 11621 35071
rect 11621 35037 11655 35071
rect 11655 35037 11664 35071
rect 11612 35028 11664 35037
rect 11796 35028 11848 35080
rect 12624 34960 12676 35012
rect 14004 35028 14056 35080
rect 16120 35232 16172 35284
rect 17224 35232 17276 35284
rect 17408 35232 17460 35284
rect 19892 35232 19944 35284
rect 14556 35139 14608 35148
rect 14556 35105 14565 35139
rect 14565 35105 14599 35139
rect 14599 35105 14608 35139
rect 14556 35096 14608 35105
rect 16304 35028 16356 35080
rect 17224 35096 17276 35148
rect 15016 34960 15068 35012
rect 17684 35028 17736 35080
rect 18420 35071 18472 35080
rect 18420 35037 18429 35071
rect 18429 35037 18463 35071
rect 18463 35037 18472 35071
rect 18420 35028 18472 35037
rect 18880 35164 18932 35216
rect 12256 34892 12308 34944
rect 12716 34892 12768 34944
rect 15108 34892 15160 34944
rect 16856 34892 16908 34944
rect 19064 35028 19116 35080
rect 20904 35232 20956 35284
rect 21916 35232 21968 35284
rect 22560 35232 22612 35284
rect 24124 35232 24176 35284
rect 22376 35139 22428 35148
rect 22376 35105 22385 35139
rect 22385 35105 22419 35139
rect 22419 35105 22428 35139
rect 22376 35096 22428 35105
rect 20812 35028 20864 35080
rect 21824 35028 21876 35080
rect 21272 34960 21324 35012
rect 22468 35028 22520 35080
rect 22560 35071 22612 35080
rect 22560 35037 22569 35071
rect 22569 35037 22603 35071
rect 22603 35037 22612 35071
rect 22560 35028 22612 35037
rect 23572 35071 23624 35080
rect 23572 35037 23581 35071
rect 23581 35037 23615 35071
rect 23615 35037 23624 35071
rect 23572 35028 23624 35037
rect 22744 34935 22796 34944
rect 22744 34901 22753 34935
rect 22753 34901 22787 34935
rect 22787 34901 22796 34935
rect 22744 34892 22796 34901
rect 35164 34892 35216 34944
rect 9390 34790 9442 34842
rect 9454 34790 9506 34842
rect 9518 34790 9570 34842
rect 9582 34790 9634 34842
rect 9646 34790 9698 34842
rect 17831 34790 17883 34842
rect 17895 34790 17947 34842
rect 17959 34790 18011 34842
rect 18023 34790 18075 34842
rect 18087 34790 18139 34842
rect 26272 34790 26324 34842
rect 26336 34790 26388 34842
rect 26400 34790 26452 34842
rect 26464 34790 26516 34842
rect 26528 34790 26580 34842
rect 34713 34790 34765 34842
rect 34777 34790 34829 34842
rect 34841 34790 34893 34842
rect 34905 34790 34957 34842
rect 34969 34790 35021 34842
rect 10048 34688 10100 34740
rect 11244 34688 11296 34740
rect 11336 34731 11388 34740
rect 11336 34697 11345 34731
rect 11345 34697 11379 34731
rect 11379 34697 11388 34731
rect 11336 34688 11388 34697
rect 8576 34484 8628 34536
rect 9220 34595 9272 34604
rect 9220 34561 9229 34595
rect 9229 34561 9263 34595
rect 9263 34561 9272 34595
rect 9220 34552 9272 34561
rect 9956 34595 10008 34604
rect 9956 34561 9965 34595
rect 9965 34561 9999 34595
rect 9999 34561 10008 34595
rect 9956 34552 10008 34561
rect 10048 34552 10100 34604
rect 10784 34527 10836 34536
rect 10784 34493 10793 34527
rect 10793 34493 10827 34527
rect 10827 34493 10836 34527
rect 10784 34484 10836 34493
rect 12532 34688 12584 34740
rect 12992 34688 13044 34740
rect 13360 34731 13412 34740
rect 13360 34697 13369 34731
rect 13369 34697 13403 34731
rect 13403 34697 13412 34731
rect 13360 34688 13412 34697
rect 15016 34731 15068 34740
rect 15016 34697 15025 34731
rect 15025 34697 15059 34731
rect 15059 34697 15068 34731
rect 15016 34688 15068 34697
rect 16028 34731 16080 34740
rect 16028 34697 16037 34731
rect 16037 34697 16071 34731
rect 16071 34697 16080 34731
rect 16028 34688 16080 34697
rect 16120 34688 16172 34740
rect 16212 34688 16264 34740
rect 16304 34688 16356 34740
rect 16856 34688 16908 34740
rect 17224 34731 17276 34740
rect 17224 34697 17233 34731
rect 17233 34697 17267 34731
rect 17267 34697 17276 34731
rect 17224 34688 17276 34697
rect 18880 34688 18932 34740
rect 19064 34688 19116 34740
rect 19340 34688 19392 34740
rect 20628 34731 20680 34740
rect 20628 34697 20637 34731
rect 20637 34697 20671 34731
rect 20671 34697 20680 34731
rect 20628 34688 20680 34697
rect 24124 34688 24176 34740
rect 13084 34620 13136 34672
rect 11612 34595 11664 34604
rect 11612 34561 11621 34595
rect 11621 34561 11655 34595
rect 11655 34561 11664 34595
rect 11612 34552 11664 34561
rect 11704 34552 11756 34604
rect 12992 34552 13044 34604
rect 14740 34552 14792 34604
rect 15660 34552 15712 34604
rect 9680 34416 9732 34468
rect 11704 34416 11756 34468
rect 8944 34391 8996 34400
rect 8944 34357 8953 34391
rect 8953 34357 8987 34391
rect 8987 34357 8996 34391
rect 8944 34348 8996 34357
rect 10508 34348 10560 34400
rect 11796 34391 11848 34400
rect 11796 34357 11805 34391
rect 11805 34357 11839 34391
rect 11839 34357 11848 34391
rect 11796 34348 11848 34357
rect 14096 34416 14148 34468
rect 15844 34527 15896 34536
rect 15844 34493 15853 34527
rect 15853 34493 15887 34527
rect 15887 34493 15896 34527
rect 15844 34484 15896 34493
rect 16396 34552 16448 34604
rect 18420 34620 18472 34672
rect 19156 34620 19208 34672
rect 18972 34595 19024 34604
rect 18972 34561 18981 34595
rect 18981 34561 19015 34595
rect 19015 34561 19024 34595
rect 18972 34552 19024 34561
rect 19524 34595 19576 34604
rect 19524 34561 19558 34595
rect 19558 34561 19576 34595
rect 19524 34552 19576 34561
rect 20628 34552 20680 34604
rect 22468 34620 22520 34672
rect 24492 34595 24544 34604
rect 24492 34561 24510 34595
rect 24510 34561 24544 34595
rect 24492 34552 24544 34561
rect 22652 34484 22704 34536
rect 23020 34527 23072 34536
rect 23020 34493 23029 34527
rect 23029 34493 23063 34527
rect 23063 34493 23072 34527
rect 23020 34484 23072 34493
rect 24768 34527 24820 34536
rect 24768 34493 24777 34527
rect 24777 34493 24811 34527
rect 24811 34493 24820 34527
rect 24768 34484 24820 34493
rect 17316 34416 17368 34468
rect 12164 34348 12216 34400
rect 13360 34348 13412 34400
rect 14924 34348 14976 34400
rect 15108 34348 15160 34400
rect 15292 34391 15344 34400
rect 15292 34357 15301 34391
rect 15301 34357 15335 34391
rect 15335 34357 15344 34391
rect 15292 34348 15344 34357
rect 15384 34348 15436 34400
rect 20812 34348 20864 34400
rect 21364 34391 21416 34400
rect 21364 34357 21373 34391
rect 21373 34357 21407 34391
rect 21407 34357 21416 34391
rect 21364 34348 21416 34357
rect 24860 34391 24912 34400
rect 24860 34357 24869 34391
rect 24869 34357 24903 34391
rect 24903 34357 24912 34391
rect 24860 34348 24912 34357
rect 5170 34246 5222 34298
rect 5234 34246 5286 34298
rect 5298 34246 5350 34298
rect 5362 34246 5414 34298
rect 5426 34246 5478 34298
rect 13611 34246 13663 34298
rect 13675 34246 13727 34298
rect 13739 34246 13791 34298
rect 13803 34246 13855 34298
rect 13867 34246 13919 34298
rect 22052 34246 22104 34298
rect 22116 34246 22168 34298
rect 22180 34246 22232 34298
rect 22244 34246 22296 34298
rect 22308 34246 22360 34298
rect 30493 34246 30545 34298
rect 30557 34246 30609 34298
rect 30621 34246 30673 34298
rect 30685 34246 30737 34298
rect 30749 34246 30801 34298
rect 9220 34144 9272 34196
rect 14096 34187 14148 34196
rect 8392 34076 8444 34128
rect 14096 34153 14105 34187
rect 14105 34153 14139 34187
rect 14139 34153 14148 34187
rect 14096 34144 14148 34153
rect 14924 34144 14976 34196
rect 17684 34187 17736 34196
rect 17684 34153 17693 34187
rect 17693 34153 17727 34187
rect 17727 34153 17736 34187
rect 17684 34144 17736 34153
rect 18604 34144 18656 34196
rect 8760 34008 8812 34060
rect 13084 34076 13136 34128
rect 17500 34076 17552 34128
rect 20168 34144 20220 34196
rect 23204 34144 23256 34196
rect 8484 33983 8536 33992
rect 8484 33949 8493 33983
rect 8493 33949 8527 33983
rect 8527 33949 8536 33983
rect 8484 33940 8536 33949
rect 8944 33940 8996 33992
rect 8852 33872 8904 33924
rect 11980 33940 12032 33992
rect 13452 34051 13504 34060
rect 13452 34017 13461 34051
rect 13461 34017 13495 34051
rect 13495 34017 13504 34051
rect 13452 34008 13504 34017
rect 12532 33983 12584 33992
rect 12532 33949 12541 33983
rect 12541 33949 12575 33983
rect 12575 33949 12584 33983
rect 12532 33940 12584 33949
rect 14556 34008 14608 34060
rect 13820 33940 13872 33992
rect 14004 33940 14056 33992
rect 15292 33940 15344 33992
rect 18696 34008 18748 34060
rect 9772 33872 9824 33924
rect 10416 33915 10468 33924
rect 10416 33881 10425 33915
rect 10425 33881 10459 33915
rect 10459 33881 10468 33915
rect 10416 33872 10468 33881
rect 11704 33872 11756 33924
rect 8300 33847 8352 33856
rect 8300 33813 8309 33847
rect 8309 33813 8343 33847
rect 8343 33813 8352 33847
rect 8300 33804 8352 33813
rect 9220 33804 9272 33856
rect 10876 33804 10928 33856
rect 12164 33804 12216 33856
rect 12256 33847 12308 33856
rect 12256 33813 12265 33847
rect 12265 33813 12299 33847
rect 12299 33813 12308 33847
rect 12256 33804 12308 33813
rect 13728 33847 13780 33856
rect 13728 33813 13755 33847
rect 13755 33813 13780 33847
rect 13728 33804 13780 33813
rect 14188 33872 14240 33924
rect 14372 33872 14424 33924
rect 14004 33804 14056 33856
rect 15016 33804 15068 33856
rect 15936 33804 15988 33856
rect 18236 33940 18288 33992
rect 24860 34008 24912 34060
rect 19800 33983 19852 33992
rect 19800 33949 19809 33983
rect 19809 33949 19843 33983
rect 19843 33949 19852 33983
rect 19800 33940 19852 33949
rect 20812 33940 20864 33992
rect 18788 33915 18840 33924
rect 18788 33881 18797 33915
rect 18797 33881 18831 33915
rect 18831 33881 18840 33915
rect 18788 33872 18840 33881
rect 16948 33804 17000 33856
rect 18512 33804 18564 33856
rect 19156 33804 19208 33856
rect 19524 33804 19576 33856
rect 19708 33804 19760 33856
rect 20720 33804 20772 33856
rect 20996 33847 21048 33856
rect 20996 33813 21005 33847
rect 21005 33813 21039 33847
rect 21039 33813 21048 33847
rect 20996 33804 21048 33813
rect 24032 33940 24084 33992
rect 22284 33872 22336 33924
rect 22744 33915 22796 33924
rect 22744 33881 22778 33915
rect 22778 33881 22796 33915
rect 22744 33872 22796 33881
rect 23572 33872 23624 33924
rect 23848 33847 23900 33856
rect 23848 33813 23857 33847
rect 23857 33813 23891 33847
rect 23891 33813 23900 33847
rect 23848 33804 23900 33813
rect 23940 33847 23992 33856
rect 23940 33813 23949 33847
rect 23949 33813 23983 33847
rect 23983 33813 23992 33847
rect 23940 33804 23992 33813
rect 24308 33804 24360 33856
rect 9390 33702 9442 33754
rect 9454 33702 9506 33754
rect 9518 33702 9570 33754
rect 9582 33702 9634 33754
rect 9646 33702 9698 33754
rect 17831 33702 17883 33754
rect 17895 33702 17947 33754
rect 17959 33702 18011 33754
rect 18023 33702 18075 33754
rect 18087 33702 18139 33754
rect 26272 33702 26324 33754
rect 26336 33702 26388 33754
rect 26400 33702 26452 33754
rect 26464 33702 26516 33754
rect 26528 33702 26580 33754
rect 34713 33702 34765 33754
rect 34777 33702 34829 33754
rect 34841 33702 34893 33754
rect 34905 33702 34957 33754
rect 34969 33702 35021 33754
rect 8300 33600 8352 33652
rect 9312 33600 9364 33652
rect 10048 33600 10100 33652
rect 11244 33600 11296 33652
rect 13728 33600 13780 33652
rect 14280 33600 14332 33652
rect 15844 33600 15896 33652
rect 12164 33532 12216 33584
rect 12624 33507 12676 33516
rect 13820 33532 13872 33584
rect 12624 33473 12642 33507
rect 12642 33473 12676 33507
rect 12624 33464 12676 33473
rect 13544 33464 13596 33516
rect 14740 33507 14792 33516
rect 14740 33473 14749 33507
rect 14749 33473 14783 33507
rect 14783 33473 14792 33507
rect 14740 33464 14792 33473
rect 14924 33464 14976 33516
rect 7380 33439 7432 33448
rect 7380 33405 7389 33439
rect 7389 33405 7423 33439
rect 7423 33405 7432 33439
rect 7380 33396 7432 33405
rect 8760 33303 8812 33312
rect 8760 33269 8769 33303
rect 8769 33269 8803 33303
rect 8803 33269 8812 33303
rect 8760 33260 8812 33269
rect 11520 33303 11572 33312
rect 11520 33269 11529 33303
rect 11529 33269 11563 33303
rect 11563 33269 11572 33303
rect 11520 33260 11572 33269
rect 13360 33396 13412 33448
rect 14464 33439 14516 33448
rect 14464 33405 14473 33439
rect 14473 33405 14507 33439
rect 14507 33405 14516 33439
rect 14464 33396 14516 33405
rect 15476 33464 15528 33516
rect 18236 33600 18288 33652
rect 15752 33396 15804 33448
rect 16120 33507 16172 33516
rect 16120 33473 16129 33507
rect 16129 33473 16163 33507
rect 16163 33473 16172 33507
rect 16120 33464 16172 33473
rect 16580 33464 16632 33516
rect 16856 33507 16908 33516
rect 16856 33473 16865 33507
rect 16865 33473 16899 33507
rect 16899 33473 16908 33507
rect 16856 33464 16908 33473
rect 16948 33507 17000 33516
rect 16948 33473 16957 33507
rect 16957 33473 16991 33507
rect 16991 33473 17000 33507
rect 16948 33464 17000 33473
rect 17132 33507 17184 33516
rect 17132 33473 17141 33507
rect 17141 33473 17175 33507
rect 17175 33473 17184 33507
rect 17132 33464 17184 33473
rect 16212 33396 16264 33448
rect 18052 33507 18104 33516
rect 18052 33473 18061 33507
rect 18061 33473 18095 33507
rect 18095 33473 18104 33507
rect 18052 33464 18104 33473
rect 19708 33600 19760 33652
rect 19800 33600 19852 33652
rect 23020 33600 23072 33652
rect 23940 33600 23992 33652
rect 24492 33600 24544 33652
rect 24768 33600 24820 33652
rect 19156 33532 19208 33584
rect 15660 33371 15712 33380
rect 15660 33337 15669 33371
rect 15669 33337 15703 33371
rect 15703 33337 15712 33371
rect 15660 33328 15712 33337
rect 17316 33328 17368 33380
rect 18512 33328 18564 33380
rect 12716 33260 12768 33312
rect 13084 33303 13136 33312
rect 13084 33269 13093 33303
rect 13093 33269 13127 33303
rect 13127 33269 13136 33303
rect 13084 33260 13136 33269
rect 14372 33260 14424 33312
rect 14924 33260 14976 33312
rect 15568 33260 15620 33312
rect 16304 33260 16356 33312
rect 18696 33260 18748 33312
rect 20168 33507 20220 33516
rect 20168 33473 20177 33507
rect 20177 33473 20211 33507
rect 20211 33473 20220 33507
rect 21364 33532 21416 33584
rect 20168 33464 20220 33473
rect 20996 33464 21048 33516
rect 24032 33507 24084 33516
rect 24032 33473 24041 33507
rect 24041 33473 24075 33507
rect 24075 33473 24084 33507
rect 24032 33464 24084 33473
rect 24216 33507 24268 33516
rect 24216 33473 24225 33507
rect 24225 33473 24259 33507
rect 24259 33473 24268 33507
rect 24216 33464 24268 33473
rect 24308 33507 24360 33516
rect 24308 33473 24317 33507
rect 24317 33473 24351 33507
rect 24351 33473 24360 33507
rect 24308 33464 24360 33473
rect 19524 33328 19576 33380
rect 19616 33371 19668 33380
rect 19616 33337 19625 33371
rect 19625 33337 19659 33371
rect 19659 33337 19668 33371
rect 19616 33328 19668 33337
rect 19800 33260 19852 33312
rect 20168 33260 20220 33312
rect 20444 33303 20496 33312
rect 20444 33269 20453 33303
rect 20453 33269 20487 33303
rect 20487 33269 20496 33303
rect 20444 33260 20496 33269
rect 21088 33260 21140 33312
rect 22836 33260 22888 33312
rect 23296 33260 23348 33312
rect 5170 33158 5222 33210
rect 5234 33158 5286 33210
rect 5298 33158 5350 33210
rect 5362 33158 5414 33210
rect 5426 33158 5478 33210
rect 13611 33158 13663 33210
rect 13675 33158 13727 33210
rect 13739 33158 13791 33210
rect 13803 33158 13855 33210
rect 13867 33158 13919 33210
rect 22052 33158 22104 33210
rect 22116 33158 22168 33210
rect 22180 33158 22232 33210
rect 22244 33158 22296 33210
rect 22308 33158 22360 33210
rect 30493 33158 30545 33210
rect 30557 33158 30609 33210
rect 30621 33158 30673 33210
rect 30685 33158 30737 33210
rect 30749 33158 30801 33210
rect 8484 33056 8536 33108
rect 10048 33056 10100 33108
rect 10784 33056 10836 33108
rect 12532 33056 12584 33108
rect 14096 33056 14148 33108
rect 14740 33056 14792 33108
rect 16120 33099 16172 33108
rect 16120 33065 16129 33099
rect 16129 33065 16163 33099
rect 16163 33065 16172 33099
rect 16120 33056 16172 33065
rect 16856 33056 16908 33108
rect 7932 32988 7984 33040
rect 8760 32988 8812 33040
rect 8576 32852 8628 32904
rect 8300 32784 8352 32836
rect 7840 32716 7892 32768
rect 9036 32852 9088 32904
rect 9220 32895 9272 32904
rect 9220 32861 9254 32895
rect 9254 32861 9272 32895
rect 9220 32852 9272 32861
rect 12256 32920 12308 32972
rect 15476 32988 15528 33040
rect 14464 32920 14516 32972
rect 14740 32963 14792 32972
rect 14740 32929 14749 32963
rect 14749 32929 14783 32963
rect 14783 32929 14792 32963
rect 14740 32920 14792 32929
rect 15660 32920 15712 32972
rect 15752 32920 15804 32972
rect 9128 32784 9180 32836
rect 11520 32852 11572 32904
rect 13084 32852 13136 32904
rect 14280 32852 14332 32904
rect 14648 32895 14700 32904
rect 14648 32861 14657 32895
rect 14657 32861 14691 32895
rect 14691 32861 14700 32895
rect 14648 32852 14700 32861
rect 14832 32784 14884 32836
rect 9772 32716 9824 32768
rect 10324 32716 10376 32768
rect 11336 32716 11388 32768
rect 11520 32759 11572 32768
rect 11520 32725 11529 32759
rect 11529 32725 11563 32759
rect 11563 32725 11572 32759
rect 11520 32716 11572 32725
rect 12716 32716 12768 32768
rect 16212 32852 16264 32904
rect 17408 32988 17460 33040
rect 15476 32784 15528 32836
rect 16212 32716 16264 32768
rect 17132 32784 17184 32836
rect 17592 32784 17644 32836
rect 17776 32895 17828 32904
rect 17776 32861 17785 32895
rect 17785 32861 17819 32895
rect 17819 32861 17828 32895
rect 17776 32852 17828 32861
rect 18052 33056 18104 33108
rect 19616 33056 19668 33108
rect 20444 33056 20496 33108
rect 21088 33099 21140 33108
rect 21088 33065 21097 33099
rect 21097 33065 21131 33099
rect 21131 33065 21140 33099
rect 21088 33056 21140 33065
rect 22376 33056 22428 33108
rect 22560 33056 22612 33108
rect 24216 33056 24268 33108
rect 19800 32988 19852 33040
rect 20076 32988 20128 33040
rect 20720 32920 20772 32972
rect 18144 32852 18196 32904
rect 18604 32852 18656 32904
rect 19524 32895 19576 32904
rect 19524 32861 19533 32895
rect 19533 32861 19567 32895
rect 19567 32861 19576 32895
rect 19524 32852 19576 32861
rect 20076 32852 20128 32904
rect 20352 32895 20404 32904
rect 20352 32861 20361 32895
rect 20361 32861 20395 32895
rect 20395 32861 20404 32895
rect 20352 32852 20404 32861
rect 22836 32920 22888 32972
rect 21364 32895 21416 32904
rect 21364 32861 21373 32895
rect 21373 32861 21407 32895
rect 21407 32861 21416 32895
rect 21364 32852 21416 32861
rect 18788 32716 18840 32768
rect 19340 32716 19392 32768
rect 19800 32716 19852 32768
rect 22468 32895 22520 32904
rect 22468 32861 22477 32895
rect 22477 32861 22511 32895
rect 22511 32861 22520 32895
rect 22468 32852 22520 32861
rect 23296 32920 23348 32972
rect 22744 32784 22796 32836
rect 23848 32852 23900 32904
rect 25320 32895 25372 32904
rect 25320 32861 25329 32895
rect 25329 32861 25363 32895
rect 25363 32861 25372 32895
rect 25320 32852 25372 32861
rect 25504 32784 25556 32836
rect 20260 32716 20312 32768
rect 23480 32759 23532 32768
rect 23480 32725 23489 32759
rect 23489 32725 23523 32759
rect 23523 32725 23532 32759
rect 23480 32716 23532 32725
rect 24400 32759 24452 32768
rect 24400 32725 24409 32759
rect 24409 32725 24443 32759
rect 24443 32725 24452 32759
rect 24400 32716 24452 32725
rect 9390 32614 9442 32666
rect 9454 32614 9506 32666
rect 9518 32614 9570 32666
rect 9582 32614 9634 32666
rect 9646 32614 9698 32666
rect 17831 32614 17883 32666
rect 17895 32614 17947 32666
rect 17959 32614 18011 32666
rect 18023 32614 18075 32666
rect 18087 32614 18139 32666
rect 26272 32614 26324 32666
rect 26336 32614 26388 32666
rect 26400 32614 26452 32666
rect 26464 32614 26516 32666
rect 26528 32614 26580 32666
rect 34713 32614 34765 32666
rect 34777 32614 34829 32666
rect 34841 32614 34893 32666
rect 34905 32614 34957 32666
rect 34969 32614 35021 32666
rect 8484 32444 8536 32496
rect 7840 32419 7892 32428
rect 7840 32385 7849 32419
rect 7849 32385 7883 32419
rect 7883 32385 7892 32419
rect 7840 32376 7892 32385
rect 7932 32419 7984 32428
rect 7932 32385 7941 32419
rect 7941 32385 7975 32419
rect 7975 32385 7984 32419
rect 7932 32376 7984 32385
rect 8116 32376 8168 32428
rect 8392 32351 8444 32360
rect 8392 32317 8401 32351
rect 8401 32317 8435 32351
rect 8435 32317 8444 32351
rect 8392 32308 8444 32317
rect 8852 32308 8904 32360
rect 10232 32555 10284 32564
rect 10232 32521 10241 32555
rect 10241 32521 10275 32555
rect 10275 32521 10284 32555
rect 10232 32512 10284 32521
rect 10784 32512 10836 32564
rect 9128 32444 9180 32496
rect 9312 32419 9364 32428
rect 9312 32385 9321 32419
rect 9321 32385 9355 32419
rect 9355 32385 9364 32419
rect 9312 32376 9364 32385
rect 9864 32444 9916 32496
rect 9680 32419 9732 32428
rect 9680 32385 9689 32419
rect 9689 32385 9723 32419
rect 9723 32385 9732 32419
rect 9680 32376 9732 32385
rect 9956 32419 10008 32428
rect 9956 32385 9965 32419
rect 9965 32385 9999 32419
rect 9999 32385 10008 32419
rect 9956 32376 10008 32385
rect 10048 32419 10100 32428
rect 10048 32385 10057 32419
rect 10057 32385 10091 32419
rect 10091 32385 10100 32419
rect 10048 32376 10100 32385
rect 10600 32444 10652 32496
rect 10692 32444 10744 32496
rect 10508 32376 10560 32428
rect 11152 32444 11204 32496
rect 10876 32419 10928 32428
rect 10876 32385 10885 32419
rect 10885 32385 10919 32419
rect 10919 32385 10928 32419
rect 10876 32376 10928 32385
rect 11520 32512 11572 32564
rect 13360 32555 13412 32564
rect 13360 32521 13369 32555
rect 13369 32521 13403 32555
rect 13403 32521 13412 32555
rect 13360 32512 13412 32521
rect 14004 32512 14056 32564
rect 14648 32512 14700 32564
rect 14740 32512 14792 32564
rect 14832 32555 14884 32564
rect 14832 32521 14841 32555
rect 14841 32521 14875 32555
rect 14875 32521 14884 32555
rect 14832 32512 14884 32521
rect 13452 32444 13504 32496
rect 9220 32240 9272 32292
rect 8944 32215 8996 32224
rect 8944 32181 8953 32215
rect 8953 32181 8987 32215
rect 8987 32181 8996 32215
rect 8944 32172 8996 32181
rect 14096 32419 14148 32428
rect 14096 32385 14105 32419
rect 14105 32385 14139 32419
rect 14139 32385 14148 32419
rect 14096 32376 14148 32385
rect 14188 32376 14240 32428
rect 9864 32172 9916 32224
rect 10600 32172 10652 32224
rect 11428 32172 11480 32224
rect 12716 32172 12768 32224
rect 14280 32308 14332 32360
rect 14096 32240 14148 32292
rect 14832 32419 14884 32428
rect 14832 32385 14841 32419
rect 14841 32385 14875 32419
rect 14875 32385 14884 32419
rect 14832 32376 14884 32385
rect 15476 32512 15528 32564
rect 15660 32512 15712 32564
rect 16580 32512 16632 32564
rect 15016 32419 15068 32428
rect 15016 32385 15025 32419
rect 15025 32385 15059 32419
rect 15059 32385 15068 32419
rect 15016 32376 15068 32385
rect 15568 32419 15620 32428
rect 15568 32385 15577 32419
rect 15577 32385 15611 32419
rect 15611 32385 15620 32419
rect 15568 32376 15620 32385
rect 15108 32308 15160 32360
rect 15292 32308 15344 32360
rect 15752 32376 15804 32428
rect 16304 32376 16356 32428
rect 15844 32308 15896 32360
rect 14372 32215 14424 32224
rect 14372 32181 14381 32215
rect 14381 32181 14415 32215
rect 14415 32181 14424 32215
rect 14372 32172 14424 32181
rect 14556 32172 14608 32224
rect 17132 32376 17184 32428
rect 17224 32419 17276 32428
rect 17224 32385 17233 32419
rect 17233 32385 17267 32419
rect 17267 32385 17276 32419
rect 17224 32376 17276 32385
rect 17316 32419 17368 32428
rect 17316 32385 17325 32419
rect 17325 32385 17359 32419
rect 17359 32385 17368 32419
rect 17316 32376 17368 32385
rect 18788 32512 18840 32564
rect 20352 32512 20404 32564
rect 23664 32555 23716 32564
rect 23664 32521 23673 32555
rect 23673 32521 23707 32555
rect 23707 32521 23716 32555
rect 23664 32512 23716 32521
rect 23848 32555 23900 32564
rect 23848 32521 23857 32555
rect 23857 32521 23891 32555
rect 23891 32521 23900 32555
rect 23848 32512 23900 32521
rect 24032 32512 24084 32564
rect 24400 32512 24452 32564
rect 24492 32512 24544 32564
rect 25320 32512 25372 32564
rect 25504 32555 25556 32564
rect 25504 32521 25513 32555
rect 25513 32521 25547 32555
rect 25547 32521 25556 32555
rect 25504 32512 25556 32521
rect 18788 32376 18840 32428
rect 19432 32376 19484 32428
rect 19616 32376 19668 32428
rect 19800 32419 19852 32428
rect 19800 32385 19809 32419
rect 19809 32385 19843 32419
rect 19843 32385 19852 32419
rect 19800 32376 19852 32385
rect 20076 32376 20128 32428
rect 15660 32172 15712 32224
rect 17684 32308 17736 32360
rect 17776 32351 17828 32360
rect 17776 32317 17785 32351
rect 17785 32317 17819 32351
rect 17819 32317 17828 32351
rect 17776 32308 17828 32317
rect 18236 32351 18288 32360
rect 18236 32317 18245 32351
rect 18245 32317 18279 32351
rect 18279 32317 18288 32351
rect 18236 32308 18288 32317
rect 18972 32240 19024 32292
rect 19156 32283 19208 32292
rect 19156 32249 19165 32283
rect 19165 32249 19199 32283
rect 19199 32249 19208 32283
rect 19156 32240 19208 32249
rect 20076 32240 20128 32292
rect 22836 32419 22888 32428
rect 22836 32385 22845 32419
rect 22845 32385 22879 32419
rect 22879 32385 22888 32419
rect 22836 32376 22888 32385
rect 22928 32419 22980 32428
rect 22928 32385 22937 32419
rect 22937 32385 22971 32419
rect 22971 32385 22980 32419
rect 22928 32376 22980 32385
rect 23388 32444 23440 32496
rect 23204 32419 23256 32428
rect 23204 32385 23213 32419
rect 23213 32385 23247 32419
rect 23247 32385 23256 32419
rect 23204 32376 23256 32385
rect 21088 32351 21140 32360
rect 21088 32317 21097 32351
rect 21097 32317 21131 32351
rect 21131 32317 21140 32351
rect 21088 32308 21140 32317
rect 21456 32240 21508 32292
rect 23204 32240 23256 32292
rect 16856 32172 16908 32224
rect 17592 32215 17644 32224
rect 17592 32181 17601 32215
rect 17601 32181 17635 32215
rect 17635 32181 17644 32215
rect 17592 32172 17644 32181
rect 19432 32215 19484 32224
rect 19432 32181 19441 32215
rect 19441 32181 19475 32215
rect 19475 32181 19484 32215
rect 19432 32172 19484 32181
rect 22468 32215 22520 32224
rect 22468 32181 22477 32215
rect 22477 32181 22511 32215
rect 22511 32181 22520 32215
rect 22468 32172 22520 32181
rect 23020 32172 23072 32224
rect 23296 32172 23348 32224
rect 23940 32351 23992 32360
rect 23940 32317 23949 32351
rect 23949 32317 23983 32351
rect 23983 32317 23992 32351
rect 23940 32308 23992 32317
rect 25780 32172 25832 32224
rect 5170 32070 5222 32122
rect 5234 32070 5286 32122
rect 5298 32070 5350 32122
rect 5362 32070 5414 32122
rect 5426 32070 5478 32122
rect 13611 32070 13663 32122
rect 13675 32070 13727 32122
rect 13739 32070 13791 32122
rect 13803 32070 13855 32122
rect 13867 32070 13919 32122
rect 22052 32070 22104 32122
rect 22116 32070 22168 32122
rect 22180 32070 22232 32122
rect 22244 32070 22296 32122
rect 22308 32070 22360 32122
rect 30493 32070 30545 32122
rect 30557 32070 30609 32122
rect 30621 32070 30673 32122
rect 30685 32070 30737 32122
rect 30749 32070 30801 32122
rect 8852 31968 8904 32020
rect 9680 31968 9732 32020
rect 11060 31968 11112 32020
rect 11152 31968 11204 32020
rect 10324 31943 10376 31952
rect 10324 31909 10333 31943
rect 10333 31909 10367 31943
rect 10367 31909 10376 31943
rect 10324 31900 10376 31909
rect 14096 31968 14148 32020
rect 14832 31968 14884 32020
rect 15844 32011 15896 32020
rect 15844 31977 15853 32011
rect 15853 31977 15887 32011
rect 15887 31977 15896 32011
rect 15844 31968 15896 31977
rect 14648 31900 14700 31952
rect 7380 31875 7432 31884
rect 7380 31841 7389 31875
rect 7389 31841 7423 31875
rect 7423 31841 7432 31875
rect 7380 31832 7432 31841
rect 12256 31832 12308 31884
rect 13820 31875 13872 31884
rect 13820 31841 13829 31875
rect 13829 31841 13863 31875
rect 13863 31841 13872 31875
rect 13820 31832 13872 31841
rect 16212 31875 16264 31884
rect 16212 31841 16221 31875
rect 16221 31841 16255 31875
rect 16255 31841 16264 31875
rect 16212 31832 16264 31841
rect 9036 31764 9088 31816
rect 9220 31807 9272 31816
rect 9220 31773 9254 31807
rect 9254 31773 9272 31807
rect 9220 31764 9272 31773
rect 12716 31764 12768 31816
rect 13452 31764 13504 31816
rect 14096 31764 14148 31816
rect 14188 31764 14240 31816
rect 15936 31764 15988 31816
rect 8024 31696 8076 31748
rect 11336 31696 11388 31748
rect 12348 31671 12400 31680
rect 12348 31637 12357 31671
rect 12357 31637 12391 31671
rect 12391 31637 12400 31671
rect 12348 31628 12400 31637
rect 13268 31671 13320 31680
rect 13268 31637 13277 31671
rect 13277 31637 13311 31671
rect 13311 31637 13320 31671
rect 13268 31628 13320 31637
rect 14280 31628 14332 31680
rect 14740 31628 14792 31680
rect 15476 31628 15528 31680
rect 16672 31807 16724 31816
rect 16672 31773 16681 31807
rect 16681 31773 16715 31807
rect 16715 31773 16724 31807
rect 16672 31764 16724 31773
rect 18420 31968 18472 32020
rect 17132 31900 17184 31952
rect 17040 31807 17092 31816
rect 17040 31773 17049 31807
rect 17049 31773 17083 31807
rect 17083 31773 17092 31807
rect 17040 31764 17092 31773
rect 17684 31900 17736 31952
rect 17776 31900 17828 31952
rect 18236 31900 18288 31952
rect 18788 31968 18840 32020
rect 19708 31968 19760 32020
rect 20260 31968 20312 32020
rect 21180 31968 21232 32020
rect 22100 31968 22152 32020
rect 22928 32011 22980 32020
rect 22928 31977 22937 32011
rect 22937 31977 22971 32011
rect 22971 31977 22980 32011
rect 22928 31968 22980 31977
rect 23388 32011 23440 32020
rect 23388 31977 23397 32011
rect 23397 31977 23431 32011
rect 23431 31977 23440 32011
rect 23388 31968 23440 31977
rect 23664 31968 23716 32020
rect 24032 31968 24084 32020
rect 24308 31968 24360 32020
rect 24768 31968 24820 32020
rect 25780 32011 25832 32020
rect 25780 31977 25789 32011
rect 25789 31977 25823 32011
rect 25823 31977 25832 32011
rect 25780 31968 25832 31977
rect 18604 31900 18656 31952
rect 21456 31943 21508 31952
rect 21456 31909 21465 31943
rect 21465 31909 21499 31943
rect 21499 31909 21508 31943
rect 21456 31900 21508 31909
rect 19432 31832 19484 31884
rect 16948 31739 17000 31748
rect 16948 31705 16957 31739
rect 16957 31705 16991 31739
rect 16991 31705 17000 31739
rect 16948 31696 17000 31705
rect 17224 31696 17276 31748
rect 18696 31807 18748 31816
rect 18696 31773 18705 31807
rect 18705 31773 18739 31807
rect 18739 31773 18748 31807
rect 18696 31764 18748 31773
rect 18880 31807 18932 31816
rect 18880 31773 18889 31807
rect 18889 31773 18923 31807
rect 18923 31773 18932 31807
rect 18880 31764 18932 31773
rect 18972 31807 19024 31816
rect 18972 31773 18981 31807
rect 18981 31773 19015 31807
rect 19015 31773 19024 31807
rect 18972 31764 19024 31773
rect 19524 31807 19576 31816
rect 19524 31773 19533 31807
rect 19533 31773 19567 31807
rect 19567 31773 19576 31807
rect 19524 31764 19576 31773
rect 19708 31807 19760 31816
rect 19708 31773 19717 31807
rect 19717 31773 19751 31807
rect 19751 31773 19760 31807
rect 19708 31764 19760 31773
rect 18512 31696 18564 31748
rect 18788 31696 18840 31748
rect 20076 31807 20128 31816
rect 20076 31773 20085 31807
rect 20085 31773 20119 31807
rect 20119 31773 20128 31807
rect 20076 31764 20128 31773
rect 17500 31628 17552 31680
rect 17592 31671 17644 31680
rect 17592 31637 17601 31671
rect 17601 31637 17635 31671
rect 17635 31637 17644 31671
rect 17592 31628 17644 31637
rect 20996 31671 21048 31680
rect 20996 31637 21005 31671
rect 21005 31637 21039 31671
rect 21039 31637 21048 31671
rect 20996 31628 21048 31637
rect 21824 31696 21876 31748
rect 23204 31807 23256 31816
rect 23204 31773 23213 31807
rect 23213 31773 23247 31807
rect 23247 31773 23256 31807
rect 23204 31764 23256 31773
rect 23296 31764 23348 31816
rect 22560 31739 22612 31748
rect 22560 31705 22578 31739
rect 22578 31705 22612 31739
rect 22560 31696 22612 31705
rect 24124 31764 24176 31816
rect 24492 31764 24544 31816
rect 22652 31628 22704 31680
rect 23756 31628 23808 31680
rect 23848 31628 23900 31680
rect 9390 31526 9442 31578
rect 9454 31526 9506 31578
rect 9518 31526 9570 31578
rect 9582 31526 9634 31578
rect 9646 31526 9698 31578
rect 17831 31526 17883 31578
rect 17895 31526 17947 31578
rect 17959 31526 18011 31578
rect 18023 31526 18075 31578
rect 18087 31526 18139 31578
rect 26272 31526 26324 31578
rect 26336 31526 26388 31578
rect 26400 31526 26452 31578
rect 26464 31526 26516 31578
rect 26528 31526 26580 31578
rect 34713 31526 34765 31578
rect 34777 31526 34829 31578
rect 34841 31526 34893 31578
rect 34905 31526 34957 31578
rect 34969 31526 35021 31578
rect 8024 31467 8076 31476
rect 8024 31433 8033 31467
rect 8033 31433 8067 31467
rect 8067 31433 8076 31467
rect 8024 31424 8076 31433
rect 8484 31424 8536 31476
rect 8484 31331 8536 31340
rect 8484 31297 8493 31331
rect 8493 31297 8527 31331
rect 8527 31297 8536 31331
rect 8484 31288 8536 31297
rect 8944 31356 8996 31408
rect 8760 31331 8812 31340
rect 8760 31297 8769 31331
rect 8769 31297 8803 31331
rect 8803 31297 8812 31331
rect 8760 31288 8812 31297
rect 10232 31331 10284 31340
rect 10232 31297 10241 31331
rect 10241 31297 10275 31331
rect 10275 31297 10284 31331
rect 10232 31288 10284 31297
rect 11060 31288 11112 31340
rect 13268 31356 13320 31408
rect 13820 31424 13872 31476
rect 14556 31424 14608 31476
rect 14280 31356 14332 31408
rect 11612 31288 11664 31340
rect 11796 31331 11848 31340
rect 11796 31297 11805 31331
rect 11805 31297 11839 31331
rect 11839 31297 11848 31331
rect 11796 31288 11848 31297
rect 10508 31263 10560 31272
rect 10508 31229 10517 31263
rect 10517 31229 10551 31263
rect 10551 31229 10560 31263
rect 10508 31220 10560 31229
rect 12348 31331 12400 31340
rect 12348 31297 12357 31331
rect 12357 31297 12391 31331
rect 12391 31297 12400 31331
rect 12348 31288 12400 31297
rect 12440 31331 12492 31340
rect 12440 31297 12449 31331
rect 12449 31297 12483 31331
rect 12483 31297 12492 31331
rect 12440 31288 12492 31297
rect 13360 31288 13412 31340
rect 12716 31263 12768 31272
rect 12716 31229 12725 31263
rect 12725 31229 12759 31263
rect 12759 31229 12768 31263
rect 12716 31220 12768 31229
rect 14004 31288 14056 31340
rect 14372 31331 14424 31340
rect 14372 31297 14381 31331
rect 14381 31297 14415 31331
rect 14415 31297 14424 31331
rect 14372 31288 14424 31297
rect 14464 31288 14516 31340
rect 14648 31331 14700 31340
rect 14648 31297 14657 31331
rect 14657 31297 14691 31331
rect 14691 31297 14700 31331
rect 14648 31288 14700 31297
rect 10048 31127 10100 31136
rect 10048 31093 10057 31127
rect 10057 31093 10091 31127
rect 10091 31093 10100 31127
rect 10048 31084 10100 31093
rect 11152 31127 11204 31136
rect 11152 31093 11161 31127
rect 11161 31093 11195 31127
rect 11195 31093 11204 31127
rect 11152 31084 11204 31093
rect 12532 31084 12584 31136
rect 13452 31084 13504 31136
rect 14188 31084 14240 31136
rect 14648 31152 14700 31204
rect 15016 31288 15068 31340
rect 17224 31424 17276 31476
rect 17592 31424 17644 31476
rect 19616 31424 19668 31476
rect 21088 31424 21140 31476
rect 23664 31424 23716 31476
rect 23848 31467 23900 31476
rect 23848 31433 23857 31467
rect 23857 31433 23891 31467
rect 23891 31433 23900 31467
rect 23848 31424 23900 31433
rect 23940 31467 23992 31476
rect 23940 31433 23949 31467
rect 23949 31433 23983 31467
rect 23983 31433 23992 31467
rect 23940 31424 23992 31433
rect 24124 31424 24176 31476
rect 24308 31467 24360 31476
rect 24308 31433 24317 31467
rect 24317 31433 24351 31467
rect 24351 31433 24360 31467
rect 24308 31424 24360 31433
rect 24492 31424 24544 31476
rect 16948 31356 17000 31408
rect 15568 31152 15620 31204
rect 16764 31220 16816 31272
rect 17868 31331 17920 31340
rect 17868 31297 17877 31331
rect 17877 31297 17911 31331
rect 17911 31297 17920 31331
rect 17868 31288 17920 31297
rect 18512 31356 18564 31408
rect 20996 31399 21048 31408
rect 20996 31365 21014 31399
rect 21014 31365 21048 31399
rect 20996 31356 21048 31365
rect 22100 31399 22152 31408
rect 22100 31365 22134 31399
rect 22134 31365 22152 31399
rect 22100 31356 22152 31365
rect 18236 31288 18288 31340
rect 21824 31331 21876 31340
rect 21824 31297 21833 31331
rect 21833 31297 21867 31331
rect 21867 31297 21876 31331
rect 21824 31288 21876 31297
rect 23664 31331 23716 31340
rect 23664 31297 23673 31331
rect 23673 31297 23707 31331
rect 23707 31297 23716 31331
rect 23664 31288 23716 31297
rect 24308 31288 24360 31340
rect 24676 31288 24728 31340
rect 19800 31220 19852 31272
rect 23756 31220 23808 31272
rect 24768 31220 24820 31272
rect 15016 31084 15068 31136
rect 15660 31127 15712 31136
rect 15660 31093 15669 31127
rect 15669 31093 15703 31127
rect 15703 31093 15712 31127
rect 15660 31084 15712 31093
rect 16028 31127 16080 31136
rect 16028 31093 16037 31127
rect 16037 31093 16071 31127
rect 16071 31093 16080 31127
rect 16028 31084 16080 31093
rect 18972 31084 19024 31136
rect 20352 31084 20404 31136
rect 25504 31127 25556 31136
rect 25504 31093 25513 31127
rect 25513 31093 25547 31127
rect 25547 31093 25556 31127
rect 25504 31084 25556 31093
rect 5170 30982 5222 31034
rect 5234 30982 5286 31034
rect 5298 30982 5350 31034
rect 5362 30982 5414 31034
rect 5426 30982 5478 31034
rect 13611 30982 13663 31034
rect 13675 30982 13727 31034
rect 13739 30982 13791 31034
rect 13803 30982 13855 31034
rect 13867 30982 13919 31034
rect 22052 30982 22104 31034
rect 22116 30982 22168 31034
rect 22180 30982 22232 31034
rect 22244 30982 22296 31034
rect 22308 30982 22360 31034
rect 30493 30982 30545 31034
rect 30557 30982 30609 31034
rect 30621 30982 30673 31034
rect 30685 30982 30737 31034
rect 30749 30982 30801 31034
rect 8116 30880 8168 30932
rect 10508 30880 10560 30932
rect 15752 30880 15804 30932
rect 15016 30812 15068 30864
rect 16764 30880 16816 30932
rect 16948 30880 17000 30932
rect 17500 30880 17552 30932
rect 17684 30923 17736 30932
rect 17684 30889 17693 30923
rect 17693 30889 17727 30923
rect 17727 30889 17736 30923
rect 17684 30880 17736 30889
rect 8944 30719 8996 30728
rect 8944 30685 8953 30719
rect 8953 30685 8987 30719
rect 8987 30685 8996 30719
rect 12716 30744 12768 30796
rect 19800 30744 19852 30796
rect 8944 30676 8996 30685
rect 12532 30676 12584 30728
rect 13360 30676 13412 30728
rect 13452 30676 13504 30728
rect 6920 30608 6972 30660
rect 9864 30608 9916 30660
rect 10416 30651 10468 30660
rect 10416 30617 10425 30651
rect 10425 30617 10459 30651
rect 10459 30617 10468 30651
rect 10416 30608 10468 30617
rect 14188 30608 14240 30660
rect 14464 30676 14516 30728
rect 14740 30719 14792 30728
rect 14740 30685 14749 30719
rect 14749 30685 14783 30719
rect 14783 30685 14792 30719
rect 14740 30676 14792 30685
rect 15108 30719 15160 30728
rect 15108 30685 15117 30719
rect 15117 30685 15151 30719
rect 15151 30685 15160 30719
rect 15108 30676 15160 30685
rect 15384 30676 15436 30728
rect 18236 30676 18288 30728
rect 18972 30676 19024 30728
rect 19340 30719 19392 30728
rect 19340 30685 19349 30719
rect 19349 30685 19383 30719
rect 19383 30685 19392 30719
rect 19340 30676 19392 30685
rect 19616 30719 19668 30728
rect 19616 30685 19625 30719
rect 19625 30685 19659 30719
rect 19659 30685 19668 30719
rect 19616 30676 19668 30685
rect 19892 30676 19944 30728
rect 21548 30812 21600 30864
rect 21824 30812 21876 30864
rect 22008 30812 22060 30864
rect 22652 30923 22704 30932
rect 22652 30889 22661 30923
rect 22661 30889 22695 30923
rect 22695 30889 22704 30923
rect 22652 30880 22704 30889
rect 23112 30880 23164 30932
rect 23664 30880 23716 30932
rect 25504 30880 25556 30932
rect 23480 30744 23532 30796
rect 14556 30651 14608 30660
rect 14556 30617 14565 30651
rect 14565 30617 14599 30651
rect 14599 30617 14608 30651
rect 14556 30608 14608 30617
rect 12072 30540 12124 30592
rect 14096 30583 14148 30592
rect 14096 30549 14105 30583
rect 14105 30549 14139 30583
rect 14139 30549 14148 30583
rect 14096 30540 14148 30549
rect 14280 30540 14332 30592
rect 15292 30540 15344 30592
rect 19524 30651 19576 30660
rect 19524 30617 19533 30651
rect 19533 30617 19567 30651
rect 19567 30617 19576 30651
rect 19524 30608 19576 30617
rect 17500 30583 17552 30592
rect 17500 30549 17509 30583
rect 17509 30549 17543 30583
rect 17543 30549 17552 30583
rect 17500 30540 17552 30549
rect 20260 30719 20312 30728
rect 20260 30685 20269 30719
rect 20269 30685 20303 30719
rect 20303 30685 20312 30719
rect 20260 30676 20312 30685
rect 20444 30676 20496 30728
rect 21088 30676 21140 30728
rect 22836 30719 22888 30728
rect 22836 30685 22845 30719
rect 22845 30685 22879 30719
rect 22879 30685 22888 30719
rect 22836 30676 22888 30685
rect 23204 30676 23256 30728
rect 20536 30540 20588 30592
rect 23940 30583 23992 30592
rect 23940 30549 23949 30583
rect 23949 30549 23983 30583
rect 23983 30549 23992 30583
rect 23940 30540 23992 30549
rect 9390 30438 9442 30490
rect 9454 30438 9506 30490
rect 9518 30438 9570 30490
rect 9582 30438 9634 30490
rect 9646 30438 9698 30490
rect 17831 30438 17883 30490
rect 17895 30438 17947 30490
rect 17959 30438 18011 30490
rect 18023 30438 18075 30490
rect 18087 30438 18139 30490
rect 26272 30438 26324 30490
rect 26336 30438 26388 30490
rect 26400 30438 26452 30490
rect 26464 30438 26516 30490
rect 26528 30438 26580 30490
rect 34713 30438 34765 30490
rect 34777 30438 34829 30490
rect 34841 30438 34893 30490
rect 34905 30438 34957 30490
rect 34969 30438 35021 30490
rect 10232 30336 10284 30388
rect 14648 30336 14700 30388
rect 15108 30336 15160 30388
rect 16948 30336 17000 30388
rect 17684 30336 17736 30388
rect 10048 30268 10100 30320
rect 14096 30268 14148 30320
rect 6552 30243 6604 30252
rect 6552 30209 6561 30243
rect 6561 30209 6595 30243
rect 6595 30209 6604 30243
rect 6552 30200 6604 30209
rect 8116 30243 8168 30252
rect 8116 30209 8125 30243
rect 8125 30209 8159 30243
rect 8159 30209 8168 30243
rect 8116 30200 8168 30209
rect 8944 30200 8996 30252
rect 6920 30132 6972 30184
rect 9404 30200 9456 30252
rect 11520 30243 11572 30252
rect 11520 30209 11529 30243
rect 11529 30209 11563 30243
rect 11563 30209 11572 30243
rect 11520 30200 11572 30209
rect 12716 30200 12768 30252
rect 7932 30039 7984 30048
rect 7932 30005 7941 30039
rect 7941 30005 7975 30039
rect 7975 30005 7984 30039
rect 7932 29996 7984 30005
rect 14004 30175 14056 30184
rect 14004 30141 14013 30175
rect 14013 30141 14047 30175
rect 14047 30141 14056 30175
rect 14004 30132 14056 30141
rect 11152 30064 11204 30116
rect 14556 30132 14608 30184
rect 10968 30039 11020 30048
rect 10968 30005 10977 30039
rect 10977 30005 11011 30039
rect 11011 30005 11020 30039
rect 10968 29996 11020 30005
rect 11704 30039 11756 30048
rect 11704 30005 11713 30039
rect 11713 30005 11747 30039
rect 11747 30005 11756 30039
rect 11704 29996 11756 30005
rect 13268 30039 13320 30048
rect 13268 30005 13277 30039
rect 13277 30005 13311 30039
rect 13311 30005 13320 30039
rect 13268 29996 13320 30005
rect 14004 29996 14056 30048
rect 15936 30268 15988 30320
rect 15476 30243 15528 30252
rect 15476 30209 15485 30243
rect 15485 30209 15519 30243
rect 15519 30209 15528 30243
rect 15476 30200 15528 30209
rect 15568 30243 15620 30252
rect 15568 30209 15577 30243
rect 15577 30209 15611 30243
rect 15611 30209 15620 30243
rect 15568 30200 15620 30209
rect 16764 30243 16816 30252
rect 16764 30209 16773 30243
rect 16773 30209 16807 30243
rect 16807 30209 16816 30243
rect 16764 30200 16816 30209
rect 16948 30243 17000 30252
rect 16948 30209 16957 30243
rect 16957 30209 16991 30243
rect 16991 30209 17000 30243
rect 16948 30200 17000 30209
rect 17040 30243 17092 30252
rect 17040 30209 17049 30243
rect 17049 30209 17083 30243
rect 17083 30209 17092 30243
rect 17040 30200 17092 30209
rect 17224 30243 17276 30252
rect 17224 30209 17233 30243
rect 17233 30209 17267 30243
rect 17267 30209 17276 30243
rect 17224 30200 17276 30209
rect 17500 30200 17552 30252
rect 16856 30132 16908 30184
rect 16028 30064 16080 30116
rect 16580 30064 16632 30116
rect 18696 30243 18748 30252
rect 18696 30209 18705 30243
rect 18705 30209 18739 30243
rect 18739 30209 18748 30243
rect 18696 30200 18748 30209
rect 18880 30243 18932 30252
rect 18880 30209 18889 30243
rect 18889 30209 18923 30243
rect 18923 30209 18932 30243
rect 18880 30200 18932 30209
rect 19156 30243 19208 30252
rect 19156 30209 19165 30243
rect 19165 30209 19199 30243
rect 19199 30209 19208 30243
rect 19156 30200 19208 30209
rect 20260 30336 20312 30388
rect 20444 30336 20496 30388
rect 24676 30379 24728 30388
rect 24676 30345 24685 30379
rect 24685 30345 24719 30379
rect 24719 30345 24728 30379
rect 24676 30336 24728 30345
rect 19892 30268 19944 30320
rect 21732 30268 21784 30320
rect 23204 30268 23256 30320
rect 19432 30200 19484 30252
rect 14740 30039 14792 30048
rect 14740 30005 14749 30039
rect 14749 30005 14783 30039
rect 14783 30005 14792 30039
rect 14740 29996 14792 30005
rect 15752 30039 15804 30048
rect 15752 30005 15761 30039
rect 15761 30005 15795 30039
rect 15795 30005 15804 30039
rect 15752 29996 15804 30005
rect 17132 29996 17184 30048
rect 19892 30132 19944 30184
rect 20168 30200 20220 30252
rect 20352 30200 20404 30252
rect 20996 30200 21048 30252
rect 21640 30200 21692 30252
rect 22008 30200 22060 30252
rect 23848 30200 23900 30252
rect 18788 30064 18840 30116
rect 18972 30064 19024 30116
rect 19524 30064 19576 30116
rect 18880 30039 18932 30048
rect 18880 30005 18889 30039
rect 18889 30005 18923 30039
rect 18923 30005 18932 30039
rect 18880 29996 18932 30005
rect 19340 29996 19392 30048
rect 20720 30132 20772 30184
rect 21272 30064 21324 30116
rect 20260 30039 20312 30048
rect 20260 30005 20269 30039
rect 20269 30005 20303 30039
rect 20303 30005 20312 30039
rect 20260 29996 20312 30005
rect 20536 29996 20588 30048
rect 21824 29996 21876 30048
rect 22652 29996 22704 30048
rect 23572 29996 23624 30048
rect 5170 29894 5222 29946
rect 5234 29894 5286 29946
rect 5298 29894 5350 29946
rect 5362 29894 5414 29946
rect 5426 29894 5478 29946
rect 13611 29894 13663 29946
rect 13675 29894 13727 29946
rect 13739 29894 13791 29946
rect 13803 29894 13855 29946
rect 13867 29894 13919 29946
rect 22052 29894 22104 29946
rect 22116 29894 22168 29946
rect 22180 29894 22232 29946
rect 22244 29894 22296 29946
rect 22308 29894 22360 29946
rect 30493 29894 30545 29946
rect 30557 29894 30609 29946
rect 30621 29894 30673 29946
rect 30685 29894 30737 29946
rect 30749 29894 30801 29946
rect 6552 29792 6604 29844
rect 9864 29792 9916 29844
rect 10232 29724 10284 29776
rect 10968 29724 11020 29776
rect 6000 29656 6052 29708
rect 8852 29656 8904 29708
rect 9404 29656 9456 29708
rect 11980 29792 12032 29844
rect 12716 29792 12768 29844
rect 15384 29792 15436 29844
rect 15568 29792 15620 29844
rect 16672 29792 16724 29844
rect 6092 29631 6144 29640
rect 6092 29597 6101 29631
rect 6101 29597 6135 29631
rect 6135 29597 6144 29631
rect 6092 29588 6144 29597
rect 7380 29631 7432 29640
rect 7380 29597 7389 29631
rect 7389 29597 7423 29631
rect 7423 29597 7432 29631
rect 7380 29588 7432 29597
rect 7932 29588 7984 29640
rect 9312 29588 9364 29640
rect 8484 29452 8536 29504
rect 8944 29495 8996 29504
rect 8944 29461 8953 29495
rect 8953 29461 8987 29495
rect 8987 29461 8996 29495
rect 8944 29452 8996 29461
rect 12072 29588 12124 29640
rect 12164 29631 12216 29640
rect 12164 29597 12173 29631
rect 12173 29597 12207 29631
rect 12207 29597 12216 29631
rect 12164 29588 12216 29597
rect 10692 29452 10744 29504
rect 10784 29495 10836 29504
rect 10784 29461 10793 29495
rect 10793 29461 10827 29495
rect 10827 29461 10836 29495
rect 13360 29588 13412 29640
rect 14740 29588 14792 29640
rect 12440 29520 12492 29572
rect 15476 29656 15528 29708
rect 18420 29835 18472 29844
rect 18420 29801 18429 29835
rect 18429 29801 18463 29835
rect 18463 29801 18472 29835
rect 18420 29792 18472 29801
rect 19156 29792 19208 29844
rect 19340 29792 19392 29844
rect 18512 29724 18564 29776
rect 19064 29724 19116 29776
rect 19892 29792 19944 29844
rect 21640 29792 21692 29844
rect 23848 29835 23900 29844
rect 23848 29801 23857 29835
rect 23857 29801 23891 29835
rect 23891 29801 23900 29835
rect 23848 29792 23900 29801
rect 19984 29724 20036 29776
rect 20352 29724 20404 29776
rect 21732 29767 21784 29776
rect 21732 29733 21741 29767
rect 21741 29733 21775 29767
rect 21775 29733 21784 29767
rect 21732 29724 21784 29733
rect 15292 29588 15344 29640
rect 15660 29588 15712 29640
rect 15844 29631 15896 29640
rect 15844 29597 15853 29631
rect 15853 29597 15887 29631
rect 15887 29597 15896 29631
rect 15844 29588 15896 29597
rect 10784 29452 10836 29461
rect 12348 29452 12400 29504
rect 14464 29452 14516 29504
rect 17868 29520 17920 29572
rect 18420 29588 18472 29640
rect 18604 29588 18656 29640
rect 18972 29588 19024 29640
rect 19064 29631 19116 29640
rect 19064 29597 19073 29631
rect 19073 29597 19107 29631
rect 19107 29597 19116 29631
rect 19064 29588 19116 29597
rect 19340 29588 19392 29640
rect 20444 29631 20496 29640
rect 20444 29597 20453 29631
rect 20453 29597 20487 29631
rect 20487 29597 20496 29631
rect 20444 29588 20496 29597
rect 20628 29631 20680 29640
rect 20628 29597 20637 29631
rect 20637 29597 20671 29631
rect 20671 29597 20680 29631
rect 20628 29588 20680 29597
rect 20720 29588 20772 29640
rect 20812 29588 20864 29640
rect 18052 29563 18104 29572
rect 18052 29529 18061 29563
rect 18061 29529 18095 29563
rect 18095 29529 18104 29563
rect 18052 29520 18104 29529
rect 18144 29520 18196 29572
rect 18328 29452 18380 29504
rect 18604 29495 18656 29504
rect 18604 29461 18613 29495
rect 18613 29461 18647 29495
rect 18647 29461 18656 29495
rect 18604 29452 18656 29461
rect 18696 29452 18748 29504
rect 19156 29452 19208 29504
rect 19708 29520 19760 29572
rect 21272 29588 21324 29640
rect 21824 29588 21876 29640
rect 21916 29631 21968 29640
rect 21916 29597 21925 29631
rect 21925 29597 21959 29631
rect 21959 29597 21968 29631
rect 21916 29588 21968 29597
rect 23572 29631 23624 29640
rect 23572 29597 23581 29631
rect 23581 29597 23615 29631
rect 23615 29597 23624 29631
rect 23572 29588 23624 29597
rect 23940 29588 23992 29640
rect 24032 29631 24084 29640
rect 24032 29597 24041 29631
rect 24041 29597 24075 29631
rect 24075 29597 24084 29631
rect 24032 29588 24084 29597
rect 29000 29588 29052 29640
rect 19892 29495 19944 29504
rect 19892 29461 19901 29495
rect 19901 29461 19935 29495
rect 19935 29461 19944 29495
rect 19892 29452 19944 29461
rect 21180 29452 21232 29504
rect 22744 29452 22796 29504
rect 23296 29495 23348 29504
rect 23296 29461 23305 29495
rect 23305 29461 23339 29495
rect 23339 29461 23348 29495
rect 23296 29452 23348 29461
rect 9390 29350 9442 29402
rect 9454 29350 9506 29402
rect 9518 29350 9570 29402
rect 9582 29350 9634 29402
rect 9646 29350 9698 29402
rect 17831 29350 17883 29402
rect 17895 29350 17947 29402
rect 17959 29350 18011 29402
rect 18023 29350 18075 29402
rect 18087 29350 18139 29402
rect 26272 29350 26324 29402
rect 26336 29350 26388 29402
rect 26400 29350 26452 29402
rect 26464 29350 26516 29402
rect 26528 29350 26580 29402
rect 34713 29350 34765 29402
rect 34777 29350 34829 29402
rect 34841 29350 34893 29402
rect 34905 29350 34957 29402
rect 34969 29350 35021 29402
rect 6092 29248 6144 29300
rect 8116 29248 8168 29300
rect 8944 29248 8996 29300
rect 9312 29248 9364 29300
rect 9772 29248 9824 29300
rect 11520 29248 11572 29300
rect 11796 29248 11848 29300
rect 1400 29155 1452 29164
rect 1400 29121 1409 29155
rect 1409 29121 1443 29155
rect 1443 29121 1452 29155
rect 1400 29112 1452 29121
rect 1584 29112 1636 29164
rect 6644 29112 6696 29164
rect 7380 29112 7432 29164
rect 8116 29112 8168 29164
rect 8852 29180 8904 29232
rect 9220 29180 9272 29232
rect 12256 29223 12308 29232
rect 12256 29189 12265 29223
rect 12265 29189 12299 29223
rect 12299 29189 12308 29223
rect 12256 29180 12308 29189
rect 9496 29155 9548 29164
rect 9496 29121 9505 29155
rect 9505 29121 9539 29155
rect 9539 29121 9548 29155
rect 9496 29112 9548 29121
rect 10048 29155 10100 29164
rect 10048 29121 10057 29155
rect 10057 29121 10091 29155
rect 10091 29121 10100 29155
rect 10048 29112 10100 29121
rect 10324 29112 10376 29164
rect 10784 29112 10836 29164
rect 13360 29248 13412 29300
rect 14004 29248 14056 29300
rect 14188 29291 14240 29300
rect 14188 29257 14197 29291
rect 14197 29257 14231 29291
rect 14231 29257 14240 29291
rect 14188 29248 14240 29257
rect 14464 29291 14516 29300
rect 14464 29257 14473 29291
rect 14473 29257 14507 29291
rect 14507 29257 14516 29291
rect 14464 29248 14516 29257
rect 13268 29180 13320 29232
rect 14740 29180 14792 29232
rect 13176 29155 13228 29164
rect 13176 29121 13185 29155
rect 13185 29121 13219 29155
rect 13219 29121 13228 29155
rect 13176 29112 13228 29121
rect 8484 29044 8536 29096
rect 10876 29044 10928 29096
rect 6000 28976 6052 29028
rect 9312 28976 9364 29028
rect 9956 28976 10008 29028
rect 11244 29044 11296 29096
rect 12348 28976 12400 29028
rect 14372 29155 14424 29164
rect 14372 29121 14381 29155
rect 14381 29121 14415 29155
rect 14415 29121 14424 29155
rect 14372 29112 14424 29121
rect 14096 28976 14148 29028
rect 14740 28976 14792 29028
rect 16764 29248 16816 29300
rect 16948 29248 17000 29300
rect 16580 29180 16632 29232
rect 18420 29248 18472 29300
rect 18604 29248 18656 29300
rect 18880 29248 18932 29300
rect 18972 29248 19024 29300
rect 19156 29291 19208 29300
rect 19156 29257 19165 29291
rect 19165 29257 19199 29291
rect 19199 29257 19208 29291
rect 19156 29248 19208 29257
rect 16028 29155 16080 29164
rect 16028 29121 16037 29155
rect 16037 29121 16071 29155
rect 16071 29121 16080 29155
rect 16028 29112 16080 29121
rect 16212 29112 16264 29164
rect 6184 28951 6236 28960
rect 6184 28917 6193 28951
rect 6193 28917 6227 28951
rect 6227 28917 6236 28951
rect 6184 28908 6236 28917
rect 8300 28908 8352 28960
rect 10232 28908 10284 28960
rect 10508 28951 10560 28960
rect 10508 28917 10517 28951
rect 10517 28917 10551 28951
rect 10551 28917 10560 28951
rect 10508 28908 10560 28917
rect 10600 28908 10652 28960
rect 11796 28908 11848 28960
rect 12716 28951 12768 28960
rect 12716 28917 12725 28951
rect 12725 28917 12759 28951
rect 12759 28917 12768 28951
rect 12716 28908 12768 28917
rect 12900 28951 12952 28960
rect 12900 28917 12909 28951
rect 12909 28917 12943 28951
rect 12943 28917 12952 28951
rect 12900 28908 12952 28917
rect 15660 28976 15712 29028
rect 15752 29019 15804 29028
rect 15752 28985 15761 29019
rect 15761 28985 15795 29019
rect 15795 28985 15804 29019
rect 15752 28976 15804 28985
rect 16672 29044 16724 29096
rect 16856 29155 16908 29164
rect 16856 29121 16865 29155
rect 16865 29121 16899 29155
rect 16899 29121 16908 29155
rect 16856 29112 16908 29121
rect 17684 29155 17736 29164
rect 17684 29121 17693 29155
rect 17693 29121 17727 29155
rect 17727 29121 17736 29155
rect 17684 29112 17736 29121
rect 17592 29044 17644 29096
rect 18052 29180 18104 29232
rect 18512 29180 18564 29232
rect 19248 29112 19300 29164
rect 19340 29155 19392 29164
rect 19340 29121 19349 29155
rect 19349 29121 19383 29155
rect 19383 29121 19392 29155
rect 19340 29112 19392 29121
rect 20996 29291 21048 29300
rect 20996 29257 21005 29291
rect 21005 29257 21039 29291
rect 21039 29257 21048 29291
rect 20996 29248 21048 29257
rect 23296 29248 23348 29300
rect 24032 29248 24084 29300
rect 19524 29112 19576 29164
rect 21272 29180 21324 29232
rect 19708 29112 19760 29164
rect 19892 29155 19944 29164
rect 19892 29121 19926 29155
rect 19926 29121 19944 29155
rect 19892 29112 19944 29121
rect 21180 29112 21232 29164
rect 23756 29155 23808 29164
rect 23756 29121 23765 29155
rect 23765 29121 23799 29155
rect 23799 29121 23808 29155
rect 23756 29112 23808 29121
rect 23940 29155 23992 29164
rect 23940 29121 23949 29155
rect 23949 29121 23983 29155
rect 23983 29121 23992 29155
rect 23940 29112 23992 29121
rect 16212 28908 16264 28960
rect 16764 28908 16816 28960
rect 17500 28908 17552 28960
rect 18604 28951 18656 28960
rect 18604 28917 18613 28951
rect 18613 28917 18647 28951
rect 18647 28917 18656 28951
rect 18604 28908 18656 28917
rect 19156 28976 19208 29028
rect 20352 28908 20404 28960
rect 23296 28951 23348 28960
rect 23296 28917 23305 28951
rect 23305 28917 23339 28951
rect 23339 28917 23348 28951
rect 23296 28908 23348 28917
rect 24216 28951 24268 28960
rect 24216 28917 24225 28951
rect 24225 28917 24259 28951
rect 24259 28917 24268 28951
rect 24216 28908 24268 28917
rect 5170 28806 5222 28858
rect 5234 28806 5286 28858
rect 5298 28806 5350 28858
rect 5362 28806 5414 28858
rect 5426 28806 5478 28858
rect 13611 28806 13663 28858
rect 13675 28806 13727 28858
rect 13739 28806 13791 28858
rect 13803 28806 13855 28858
rect 13867 28806 13919 28858
rect 22052 28806 22104 28858
rect 22116 28806 22168 28858
rect 22180 28806 22232 28858
rect 22244 28806 22296 28858
rect 22308 28806 22360 28858
rect 30493 28806 30545 28858
rect 30557 28806 30609 28858
rect 30621 28806 30673 28858
rect 30685 28806 30737 28858
rect 30749 28806 30801 28858
rect 6644 28704 6696 28756
rect 9312 28704 9364 28756
rect 10508 28704 10560 28756
rect 10692 28704 10744 28756
rect 11612 28704 11664 28756
rect 8300 28568 8352 28620
rect 8944 28568 8996 28620
rect 9496 28568 9548 28620
rect 9864 28568 9916 28620
rect 12164 28704 12216 28756
rect 13176 28747 13228 28756
rect 13176 28713 13185 28747
rect 13185 28713 13219 28747
rect 13219 28713 13228 28747
rect 13176 28704 13228 28713
rect 14372 28704 14424 28756
rect 16856 28704 16908 28756
rect 17592 28747 17644 28756
rect 17592 28713 17601 28747
rect 17601 28713 17635 28747
rect 17635 28713 17644 28747
rect 17592 28704 17644 28713
rect 17684 28704 17736 28756
rect 19708 28704 19760 28756
rect 20444 28704 20496 28756
rect 20536 28747 20588 28756
rect 20536 28713 20545 28747
rect 20545 28713 20579 28747
rect 20579 28713 20588 28747
rect 20536 28704 20588 28713
rect 22744 28747 22796 28756
rect 22744 28713 22753 28747
rect 22753 28713 22787 28747
rect 22787 28713 22796 28747
rect 22744 28704 22796 28713
rect 6184 28500 6236 28552
rect 8116 28500 8168 28552
rect 8208 28543 8260 28552
rect 8208 28509 8217 28543
rect 8217 28509 8251 28543
rect 8251 28509 8260 28543
rect 8208 28500 8260 28509
rect 8484 28543 8536 28552
rect 8484 28509 8493 28543
rect 8493 28509 8527 28543
rect 8527 28509 8536 28543
rect 8484 28500 8536 28509
rect 9220 28432 9272 28484
rect 9956 28500 10008 28552
rect 10232 28543 10284 28552
rect 10232 28509 10241 28543
rect 10241 28509 10275 28543
rect 10275 28509 10284 28543
rect 10232 28500 10284 28509
rect 10324 28500 10376 28552
rect 10784 28500 10836 28552
rect 10876 28500 10928 28552
rect 11704 28500 11756 28552
rect 12900 28568 12952 28620
rect 13360 28611 13412 28620
rect 13360 28577 13369 28611
rect 13369 28577 13403 28611
rect 13403 28577 13412 28611
rect 13360 28568 13412 28577
rect 16672 28679 16724 28688
rect 16672 28645 16681 28679
rect 16681 28645 16715 28679
rect 16715 28645 16724 28679
rect 16672 28636 16724 28645
rect 20628 28636 20680 28688
rect 23296 28704 23348 28756
rect 11520 28432 11572 28484
rect 12808 28500 12860 28552
rect 13544 28543 13596 28552
rect 13544 28509 13553 28543
rect 13553 28509 13587 28543
rect 13587 28509 13596 28543
rect 13544 28500 13596 28509
rect 17316 28568 17368 28620
rect 18052 28568 18104 28620
rect 18236 28611 18288 28620
rect 18236 28577 18245 28611
rect 18245 28577 18279 28611
rect 18279 28577 18288 28611
rect 18236 28568 18288 28577
rect 18604 28568 18656 28620
rect 20076 28611 20128 28620
rect 20076 28577 20085 28611
rect 20085 28577 20119 28611
rect 20119 28577 20128 28611
rect 20076 28568 20128 28577
rect 20168 28568 20220 28620
rect 13912 28432 13964 28484
rect 15200 28432 15252 28484
rect 15384 28475 15436 28484
rect 15384 28441 15402 28475
rect 15402 28441 15436 28475
rect 15384 28432 15436 28441
rect 7196 28364 7248 28416
rect 7472 28364 7524 28416
rect 9036 28407 9088 28416
rect 9036 28373 9045 28407
rect 9045 28373 9079 28407
rect 9079 28373 9088 28407
rect 9036 28364 9088 28373
rect 9956 28407 10008 28416
rect 9956 28373 9965 28407
rect 9965 28373 9999 28407
rect 9999 28373 10008 28407
rect 9956 28364 10008 28373
rect 10600 28364 10652 28416
rect 11704 28364 11756 28416
rect 14280 28364 14332 28416
rect 16028 28543 16080 28552
rect 16028 28509 16037 28543
rect 16037 28509 16071 28543
rect 16071 28509 16080 28543
rect 16028 28500 16080 28509
rect 16672 28500 16724 28552
rect 16764 28543 16816 28552
rect 16764 28509 16773 28543
rect 16773 28509 16807 28543
rect 16807 28509 16816 28543
rect 16764 28500 16816 28509
rect 20260 28500 20312 28552
rect 20996 28568 21048 28620
rect 22744 28568 22796 28620
rect 17500 28432 17552 28484
rect 22652 28500 22704 28552
rect 24216 28500 24268 28552
rect 17316 28364 17368 28416
rect 17408 28407 17460 28416
rect 17408 28373 17417 28407
rect 17417 28373 17451 28407
rect 17451 28373 17460 28407
rect 17408 28364 17460 28373
rect 18420 28407 18472 28416
rect 18420 28373 18429 28407
rect 18429 28373 18463 28407
rect 18463 28373 18472 28407
rect 18420 28364 18472 28373
rect 22284 28407 22336 28416
rect 22284 28373 22293 28407
rect 22293 28373 22327 28407
rect 22327 28373 22336 28407
rect 22284 28364 22336 28373
rect 22560 28364 22612 28416
rect 9390 28262 9442 28314
rect 9454 28262 9506 28314
rect 9518 28262 9570 28314
rect 9582 28262 9634 28314
rect 9646 28262 9698 28314
rect 17831 28262 17883 28314
rect 17895 28262 17947 28314
rect 17959 28262 18011 28314
rect 18023 28262 18075 28314
rect 18087 28262 18139 28314
rect 26272 28262 26324 28314
rect 26336 28262 26388 28314
rect 26400 28262 26452 28314
rect 26464 28262 26516 28314
rect 26528 28262 26580 28314
rect 34713 28262 34765 28314
rect 34777 28262 34829 28314
rect 34841 28262 34893 28314
rect 34905 28262 34957 28314
rect 34969 28262 35021 28314
rect 7196 28160 7248 28212
rect 8208 28160 8260 28212
rect 9956 28160 10008 28212
rect 10600 28160 10652 28212
rect 11520 28203 11572 28212
rect 11520 28169 11529 28203
rect 11529 28169 11563 28203
rect 11563 28169 11572 28203
rect 11520 28160 11572 28169
rect 11888 28160 11940 28212
rect 7472 28024 7524 28076
rect 9220 28024 9272 28076
rect 12348 28092 12400 28144
rect 11796 28067 11848 28076
rect 11796 28033 11805 28067
rect 11805 28033 11839 28067
rect 11839 28033 11848 28067
rect 11796 28024 11848 28033
rect 12716 28067 12768 28076
rect 12716 28033 12725 28067
rect 12725 28033 12759 28067
rect 12759 28033 12768 28067
rect 12716 28024 12768 28033
rect 13360 28160 13412 28212
rect 13544 28160 13596 28212
rect 15384 28160 15436 28212
rect 16212 28160 16264 28212
rect 18236 28160 18288 28212
rect 19524 28160 19576 28212
rect 20076 28160 20128 28212
rect 13176 28024 13228 28076
rect 7380 27956 7432 28008
rect 9864 27999 9916 28008
rect 9864 27965 9873 27999
rect 9873 27965 9907 27999
rect 9907 27965 9916 27999
rect 9864 27956 9916 27965
rect 12900 27956 12952 28008
rect 13268 27956 13320 28008
rect 13912 28067 13964 28076
rect 13912 28033 13921 28067
rect 13921 28033 13955 28067
rect 13955 28033 13964 28067
rect 13912 28024 13964 28033
rect 14188 28067 14240 28076
rect 14188 28033 14222 28067
rect 14222 28033 14240 28067
rect 14188 28024 14240 28033
rect 15936 28024 15988 28076
rect 8944 27931 8996 27940
rect 8944 27897 8953 27931
rect 8953 27897 8987 27931
rect 8987 27897 8996 27931
rect 8944 27888 8996 27897
rect 12256 27888 12308 27940
rect 16488 27999 16540 28008
rect 16488 27965 16497 27999
rect 16497 27965 16531 27999
rect 16531 27965 16540 27999
rect 16488 27956 16540 27965
rect 16672 27999 16724 28008
rect 16672 27965 16681 27999
rect 16681 27965 16715 27999
rect 16715 27965 16724 27999
rect 17408 28024 17460 28076
rect 17776 28024 17828 28076
rect 21364 28092 21416 28144
rect 21548 28092 21600 28144
rect 22560 28092 22612 28144
rect 18420 28024 18472 28076
rect 20352 28067 20404 28076
rect 20352 28033 20361 28067
rect 20361 28033 20395 28067
rect 20395 28033 20404 28067
rect 20352 28024 20404 28033
rect 21916 28024 21968 28076
rect 16672 27956 16724 27965
rect 7196 27863 7248 27872
rect 7196 27829 7205 27863
rect 7205 27829 7239 27863
rect 7239 27829 7248 27863
rect 7196 27820 7248 27829
rect 13452 27820 13504 27872
rect 15292 27863 15344 27872
rect 15292 27829 15301 27863
rect 15301 27829 15335 27863
rect 15335 27829 15344 27863
rect 15292 27820 15344 27829
rect 19800 27863 19852 27872
rect 19800 27829 19809 27863
rect 19809 27829 19843 27863
rect 19843 27829 19852 27863
rect 19800 27820 19852 27829
rect 21088 27863 21140 27872
rect 21088 27829 21097 27863
rect 21097 27829 21131 27863
rect 21131 27829 21140 27863
rect 21088 27820 21140 27829
rect 21456 27820 21508 27872
rect 22284 27820 22336 27872
rect 23848 27820 23900 27872
rect 5170 27718 5222 27770
rect 5234 27718 5286 27770
rect 5298 27718 5350 27770
rect 5362 27718 5414 27770
rect 5426 27718 5478 27770
rect 13611 27718 13663 27770
rect 13675 27718 13727 27770
rect 13739 27718 13791 27770
rect 13803 27718 13855 27770
rect 13867 27718 13919 27770
rect 22052 27718 22104 27770
rect 22116 27718 22168 27770
rect 22180 27718 22232 27770
rect 22244 27718 22296 27770
rect 22308 27718 22360 27770
rect 30493 27718 30545 27770
rect 30557 27718 30609 27770
rect 30621 27718 30673 27770
rect 30685 27718 30737 27770
rect 30749 27718 30801 27770
rect 9220 27616 9272 27668
rect 10876 27616 10928 27668
rect 14188 27659 14240 27668
rect 14188 27625 14197 27659
rect 14197 27625 14231 27659
rect 14231 27625 14240 27659
rect 14188 27616 14240 27625
rect 15936 27659 15988 27668
rect 15936 27625 15945 27659
rect 15945 27625 15979 27659
rect 15979 27625 15988 27659
rect 15936 27616 15988 27625
rect 16028 27659 16080 27668
rect 16028 27625 16037 27659
rect 16037 27625 16071 27659
rect 16071 27625 16080 27659
rect 16028 27616 16080 27625
rect 21272 27616 21324 27668
rect 23020 27616 23072 27668
rect 19248 27591 19300 27600
rect 19248 27557 19257 27591
rect 19257 27557 19291 27591
rect 19291 27557 19300 27591
rect 19248 27548 19300 27557
rect 19800 27548 19852 27600
rect 20720 27548 20772 27600
rect 12440 27480 12492 27532
rect 13084 27480 13136 27532
rect 7196 27412 7248 27464
rect 7380 27455 7432 27464
rect 7380 27421 7389 27455
rect 7389 27421 7423 27455
rect 7423 27421 7432 27455
rect 7380 27412 7432 27421
rect 9864 27412 9916 27464
rect 12256 27412 12308 27464
rect 12532 27412 12584 27464
rect 12900 27455 12952 27464
rect 12900 27421 12909 27455
rect 12909 27421 12943 27455
rect 12943 27421 12952 27455
rect 12900 27412 12952 27421
rect 9772 27344 9824 27396
rect 14096 27412 14148 27464
rect 15292 27412 15344 27464
rect 12624 27276 12676 27328
rect 13544 27319 13596 27328
rect 13544 27285 13553 27319
rect 13553 27285 13587 27319
rect 13587 27285 13596 27319
rect 13544 27276 13596 27285
rect 13912 27276 13964 27328
rect 15752 27412 15804 27464
rect 17132 27455 17184 27464
rect 17132 27421 17150 27455
rect 17150 27421 17184 27455
rect 17132 27412 17184 27421
rect 17776 27412 17828 27464
rect 15660 27276 15712 27328
rect 19064 27319 19116 27328
rect 19064 27285 19073 27319
rect 19073 27285 19107 27319
rect 19107 27285 19116 27319
rect 21180 27412 21232 27464
rect 21732 27523 21784 27532
rect 21732 27489 21741 27523
rect 21741 27489 21775 27523
rect 21775 27489 21784 27523
rect 21732 27480 21784 27489
rect 21640 27455 21692 27464
rect 21640 27421 21649 27455
rect 21649 27421 21683 27455
rect 21683 27421 21692 27455
rect 21640 27412 21692 27421
rect 22744 27412 22796 27464
rect 22652 27344 22704 27396
rect 23296 27455 23348 27464
rect 23296 27421 23305 27455
rect 23305 27421 23339 27455
rect 23339 27421 23348 27455
rect 23296 27412 23348 27421
rect 34520 27455 34572 27464
rect 34520 27421 34529 27455
rect 34529 27421 34563 27455
rect 34563 27421 34572 27455
rect 34520 27412 34572 27421
rect 19064 27276 19116 27285
rect 20904 27319 20956 27328
rect 20904 27285 20913 27319
rect 20913 27285 20947 27319
rect 20947 27285 20956 27319
rect 20904 27276 20956 27285
rect 20996 27276 21048 27328
rect 21180 27276 21232 27328
rect 21916 27276 21968 27328
rect 22928 27319 22980 27328
rect 22928 27285 22937 27319
rect 22937 27285 22971 27319
rect 22971 27285 22980 27319
rect 22928 27276 22980 27285
rect 23940 27319 23992 27328
rect 23940 27285 23949 27319
rect 23949 27285 23983 27319
rect 23983 27285 23992 27319
rect 23940 27276 23992 27285
rect 24584 27276 24636 27328
rect 24860 27319 24912 27328
rect 24860 27285 24869 27319
rect 24869 27285 24903 27319
rect 24903 27285 24912 27319
rect 24860 27276 24912 27285
rect 9390 27174 9442 27226
rect 9454 27174 9506 27226
rect 9518 27174 9570 27226
rect 9582 27174 9634 27226
rect 9646 27174 9698 27226
rect 17831 27174 17883 27226
rect 17895 27174 17947 27226
rect 17959 27174 18011 27226
rect 18023 27174 18075 27226
rect 18087 27174 18139 27226
rect 26272 27174 26324 27226
rect 26336 27174 26388 27226
rect 26400 27174 26452 27226
rect 26464 27174 26516 27226
rect 26528 27174 26580 27226
rect 34713 27174 34765 27226
rect 34777 27174 34829 27226
rect 34841 27174 34893 27226
rect 34905 27174 34957 27226
rect 34969 27174 35021 27226
rect 8852 27072 8904 27124
rect 10048 27072 10100 27124
rect 11980 27072 12032 27124
rect 12440 27072 12492 27124
rect 12532 27115 12584 27124
rect 12532 27081 12541 27115
rect 12541 27081 12575 27115
rect 12575 27081 12584 27115
rect 12532 27072 12584 27081
rect 13544 27072 13596 27124
rect 13912 27072 13964 27124
rect 9036 26979 9088 26988
rect 9036 26945 9045 26979
rect 9045 26945 9079 26979
rect 9079 26945 9088 26979
rect 9036 26936 9088 26945
rect 11704 27004 11756 27056
rect 12808 27004 12860 27056
rect 11152 26936 11204 26988
rect 12164 26979 12216 26988
rect 12164 26945 12173 26979
rect 12173 26945 12207 26979
rect 12207 26945 12216 26979
rect 12164 26936 12216 26945
rect 12072 26800 12124 26852
rect 13360 26936 13412 26988
rect 14004 26936 14056 26988
rect 16488 27072 16540 27124
rect 19800 27072 19852 27124
rect 20904 27072 20956 27124
rect 21456 27115 21508 27124
rect 21456 27081 21465 27115
rect 21465 27081 21499 27115
rect 21499 27081 21508 27115
rect 21456 27072 21508 27081
rect 21640 27072 21692 27124
rect 22652 27072 22704 27124
rect 22928 27072 22980 27124
rect 23296 27072 23348 27124
rect 23940 27072 23992 27124
rect 15476 27004 15528 27056
rect 15016 26800 15068 26852
rect 15660 26936 15712 26988
rect 17408 27004 17460 27056
rect 18788 26979 18840 26988
rect 15936 26868 15988 26920
rect 18788 26945 18797 26979
rect 18797 26945 18831 26979
rect 18831 26945 18840 26979
rect 18788 26936 18840 26945
rect 21364 27004 21416 27056
rect 21272 26979 21324 26988
rect 21272 26945 21281 26979
rect 21281 26945 21315 26979
rect 21315 26945 21324 26979
rect 21272 26936 21324 26945
rect 21548 26936 21600 26988
rect 23204 27004 23256 27056
rect 17132 26911 17184 26920
rect 17132 26877 17141 26911
rect 17141 26877 17175 26911
rect 17175 26877 17184 26911
rect 17132 26868 17184 26877
rect 18420 26911 18472 26920
rect 18420 26877 18429 26911
rect 18429 26877 18463 26911
rect 18463 26877 18472 26911
rect 18420 26868 18472 26877
rect 19616 26868 19668 26920
rect 17592 26800 17644 26852
rect 22284 26800 22336 26852
rect 11612 26775 11664 26784
rect 11612 26741 11621 26775
rect 11621 26741 11655 26775
rect 11655 26741 11664 26775
rect 11612 26732 11664 26741
rect 12624 26732 12676 26784
rect 12808 26732 12860 26784
rect 12992 26732 13044 26784
rect 15108 26732 15160 26784
rect 15384 26775 15436 26784
rect 15384 26741 15393 26775
rect 15393 26741 15427 26775
rect 15427 26741 15436 26775
rect 15384 26732 15436 26741
rect 15568 26775 15620 26784
rect 15568 26741 15577 26775
rect 15577 26741 15611 26775
rect 15611 26741 15620 26775
rect 15568 26732 15620 26741
rect 15752 26732 15804 26784
rect 15844 26775 15896 26784
rect 15844 26741 15853 26775
rect 15853 26741 15887 26775
rect 15887 26741 15896 26775
rect 15844 26732 15896 26741
rect 17040 26775 17092 26784
rect 17040 26741 17049 26775
rect 17049 26741 17083 26775
rect 17083 26741 17092 26775
rect 17040 26732 17092 26741
rect 17776 26775 17828 26784
rect 17776 26741 17785 26775
rect 17785 26741 17819 26775
rect 17819 26741 17828 26775
rect 17776 26732 17828 26741
rect 19708 26775 19760 26784
rect 19708 26741 19717 26775
rect 19717 26741 19751 26775
rect 19751 26741 19760 26775
rect 19708 26732 19760 26741
rect 21640 26775 21692 26784
rect 21640 26741 21649 26775
rect 21649 26741 21683 26775
rect 21683 26741 21692 26775
rect 21640 26732 21692 26741
rect 21824 26732 21876 26784
rect 22468 26732 22520 26784
rect 22744 26979 22796 26988
rect 22744 26945 22753 26979
rect 22753 26945 22787 26979
rect 22787 26945 22796 26979
rect 22744 26936 22796 26945
rect 24860 26936 24912 26988
rect 23020 26868 23072 26920
rect 24584 26775 24636 26784
rect 24584 26741 24593 26775
rect 24593 26741 24627 26775
rect 24627 26741 24636 26775
rect 24584 26732 24636 26741
rect 5170 26630 5222 26682
rect 5234 26630 5286 26682
rect 5298 26630 5350 26682
rect 5362 26630 5414 26682
rect 5426 26630 5478 26682
rect 13611 26630 13663 26682
rect 13675 26630 13727 26682
rect 13739 26630 13791 26682
rect 13803 26630 13855 26682
rect 13867 26630 13919 26682
rect 22052 26630 22104 26682
rect 22116 26630 22168 26682
rect 22180 26630 22232 26682
rect 22244 26630 22296 26682
rect 22308 26630 22360 26682
rect 30493 26630 30545 26682
rect 30557 26630 30609 26682
rect 30621 26630 30673 26682
rect 30685 26630 30737 26682
rect 30749 26630 30801 26682
rect 11612 26528 11664 26580
rect 12900 26528 12952 26580
rect 12072 26392 12124 26444
rect 12164 26392 12216 26444
rect 8300 26324 8352 26376
rect 9864 26324 9916 26376
rect 11336 26324 11388 26376
rect 10692 26256 10744 26308
rect 11980 26367 12032 26376
rect 11980 26333 11989 26367
rect 11989 26333 12023 26367
rect 12023 26333 12032 26367
rect 11980 26324 12032 26333
rect 12624 26392 12676 26444
rect 17132 26571 17184 26580
rect 17132 26537 17141 26571
rect 17141 26537 17175 26571
rect 17175 26537 17184 26571
rect 17132 26528 17184 26537
rect 19708 26528 19760 26580
rect 21088 26528 21140 26580
rect 21640 26528 21692 26580
rect 22376 26528 22428 26580
rect 12348 26324 12400 26376
rect 12992 26367 13044 26376
rect 12992 26333 13001 26367
rect 13001 26333 13035 26367
rect 13035 26333 13044 26367
rect 12992 26324 13044 26333
rect 15016 26460 15068 26512
rect 19616 26460 19668 26512
rect 11244 26231 11296 26240
rect 11244 26197 11253 26231
rect 11253 26197 11287 26231
rect 11287 26197 11296 26231
rect 11244 26188 11296 26197
rect 11612 26188 11664 26240
rect 11796 26188 11848 26240
rect 13452 26367 13504 26376
rect 13452 26333 13461 26367
rect 13461 26333 13495 26367
rect 13495 26333 13504 26367
rect 13452 26324 13504 26333
rect 14280 26367 14332 26376
rect 14280 26333 14289 26367
rect 14289 26333 14323 26367
rect 14323 26333 14332 26367
rect 14280 26324 14332 26333
rect 14648 26324 14700 26376
rect 16672 26392 16724 26444
rect 17684 26435 17736 26444
rect 17684 26401 17693 26435
rect 17693 26401 17727 26435
rect 17727 26401 17736 26435
rect 17684 26392 17736 26401
rect 15844 26367 15896 26376
rect 15844 26333 15862 26367
rect 15862 26333 15896 26367
rect 15844 26324 15896 26333
rect 16396 26367 16448 26376
rect 16396 26333 16405 26367
rect 16405 26333 16439 26367
rect 16439 26333 16448 26367
rect 16396 26324 16448 26333
rect 17040 26324 17092 26376
rect 14832 26256 14884 26308
rect 15200 26188 15252 26240
rect 16488 26256 16540 26308
rect 17776 26324 17828 26376
rect 18420 26324 18472 26376
rect 19432 26324 19484 26376
rect 15476 26188 15528 26240
rect 16948 26188 17000 26240
rect 17132 26188 17184 26240
rect 19708 26256 19760 26308
rect 20720 26299 20772 26308
rect 20720 26265 20729 26299
rect 20729 26265 20763 26299
rect 20763 26265 20772 26299
rect 20720 26256 20772 26265
rect 21456 26435 21508 26444
rect 21456 26401 21465 26435
rect 21465 26401 21499 26435
rect 21499 26401 21508 26435
rect 21456 26392 21508 26401
rect 22100 26392 22152 26444
rect 23204 26460 23256 26512
rect 21548 26324 21600 26376
rect 21732 26324 21784 26376
rect 18604 26188 18656 26240
rect 19800 26231 19852 26240
rect 19800 26197 19809 26231
rect 19809 26197 19843 26231
rect 19843 26197 19852 26231
rect 19800 26188 19852 26197
rect 20352 26231 20404 26240
rect 20352 26197 20361 26231
rect 20361 26197 20395 26231
rect 20395 26197 20404 26231
rect 20352 26188 20404 26197
rect 20996 26256 21048 26308
rect 21824 26256 21876 26308
rect 20904 26188 20956 26240
rect 21364 26188 21416 26240
rect 21916 26231 21968 26240
rect 21916 26197 21925 26231
rect 21925 26197 21959 26231
rect 21959 26197 21968 26231
rect 22652 26367 22704 26376
rect 22652 26333 22661 26367
rect 22661 26333 22695 26367
rect 22695 26333 22704 26367
rect 22652 26324 22704 26333
rect 23204 26367 23256 26376
rect 23204 26333 23213 26367
rect 23213 26333 23247 26367
rect 23247 26333 23256 26367
rect 23204 26324 23256 26333
rect 21916 26188 21968 26197
rect 23112 26188 23164 26240
rect 9390 26086 9442 26138
rect 9454 26086 9506 26138
rect 9518 26086 9570 26138
rect 9582 26086 9634 26138
rect 9646 26086 9698 26138
rect 17831 26086 17883 26138
rect 17895 26086 17947 26138
rect 17959 26086 18011 26138
rect 18023 26086 18075 26138
rect 18087 26086 18139 26138
rect 26272 26086 26324 26138
rect 26336 26086 26388 26138
rect 26400 26086 26452 26138
rect 26464 26086 26516 26138
rect 26528 26086 26580 26138
rect 34713 26086 34765 26138
rect 34777 26086 34829 26138
rect 34841 26086 34893 26138
rect 34905 26086 34957 26138
rect 34969 26086 35021 26138
rect 8300 26027 8352 26036
rect 8300 25993 8309 26027
rect 8309 25993 8343 26027
rect 8343 25993 8352 26027
rect 8300 25984 8352 25993
rect 10692 25959 10744 25968
rect 10692 25925 10701 25959
rect 10701 25925 10735 25959
rect 10735 25925 10744 25959
rect 10692 25916 10744 25925
rect 12348 25916 12400 25968
rect 13268 25916 13320 25968
rect 10416 25848 10468 25900
rect 11244 25891 11296 25900
rect 11244 25857 11253 25891
rect 11253 25857 11287 25891
rect 11287 25857 11296 25891
rect 11244 25848 11296 25857
rect 11612 25848 11664 25900
rect 12440 25891 12492 25900
rect 12440 25857 12449 25891
rect 12449 25857 12483 25891
rect 12483 25857 12492 25891
rect 12440 25848 12492 25857
rect 12624 25848 12676 25900
rect 12716 25891 12768 25900
rect 12716 25857 12725 25891
rect 12725 25857 12759 25891
rect 12759 25857 12768 25891
rect 12716 25848 12768 25857
rect 12992 25848 13044 25900
rect 13176 25848 13228 25900
rect 13544 25891 13596 25900
rect 13544 25857 13553 25891
rect 13553 25857 13587 25891
rect 13587 25857 13596 25891
rect 13544 25848 13596 25857
rect 14188 25848 14240 25900
rect 14832 25916 14884 25968
rect 15200 25916 15252 25968
rect 15568 25916 15620 25968
rect 15660 25959 15712 25968
rect 15660 25925 15669 25959
rect 15669 25925 15703 25959
rect 15703 25925 15712 25959
rect 15660 25916 15712 25925
rect 15108 25891 15160 25900
rect 15108 25857 15117 25891
rect 15117 25857 15151 25891
rect 15151 25857 15160 25891
rect 15108 25848 15160 25857
rect 15384 25848 15436 25900
rect 15752 25891 15804 25900
rect 15752 25857 15761 25891
rect 15761 25857 15795 25891
rect 15795 25857 15804 25891
rect 15752 25848 15804 25857
rect 16672 25891 16724 25900
rect 16672 25857 16681 25891
rect 16681 25857 16715 25891
rect 16715 25857 16724 25891
rect 16672 25848 16724 25857
rect 16948 25891 17000 25900
rect 16948 25857 16982 25891
rect 16982 25857 17000 25891
rect 16948 25848 17000 25857
rect 21272 25984 21324 26036
rect 21364 25984 21416 26036
rect 21916 25984 21968 26036
rect 19984 25959 20036 25968
rect 19984 25925 19993 25959
rect 19993 25925 20027 25959
rect 20027 25925 20036 25959
rect 19984 25916 20036 25925
rect 18328 25848 18380 25900
rect 19340 25848 19392 25900
rect 19800 25848 19852 25900
rect 20352 25848 20404 25900
rect 21456 25916 21508 25968
rect 21824 25916 21876 25968
rect 21088 25891 21140 25900
rect 21088 25857 21097 25891
rect 21097 25857 21131 25891
rect 21131 25857 21140 25891
rect 21088 25848 21140 25857
rect 21640 25897 21692 25900
rect 21640 25863 21649 25897
rect 21649 25863 21683 25897
rect 21683 25863 21692 25897
rect 21640 25848 21692 25863
rect 10600 25712 10652 25764
rect 11336 25644 11388 25696
rect 11980 25644 12032 25696
rect 12072 25644 12124 25696
rect 16120 25780 16172 25832
rect 16396 25780 16448 25832
rect 21364 25823 21416 25832
rect 21364 25789 21373 25823
rect 21373 25789 21407 25823
rect 21407 25789 21416 25823
rect 21364 25780 21416 25789
rect 18420 25712 18472 25764
rect 19524 25712 19576 25764
rect 22284 25891 22336 25900
rect 22284 25857 22293 25891
rect 22293 25857 22327 25891
rect 22327 25857 22336 25891
rect 22284 25848 22336 25857
rect 22652 25916 22704 25968
rect 23112 25891 23164 25900
rect 23112 25857 23121 25891
rect 23121 25857 23155 25891
rect 23155 25857 23164 25891
rect 23112 25848 23164 25857
rect 23756 25823 23808 25832
rect 23756 25789 23765 25823
rect 23765 25789 23799 25823
rect 23799 25789 23808 25823
rect 23756 25780 23808 25789
rect 23848 25780 23900 25832
rect 13176 25644 13228 25696
rect 14556 25687 14608 25696
rect 14556 25653 14565 25687
rect 14565 25653 14599 25687
rect 14599 25653 14608 25687
rect 14556 25644 14608 25653
rect 14832 25644 14884 25696
rect 15200 25644 15252 25696
rect 15936 25644 15988 25696
rect 16488 25687 16540 25696
rect 16488 25653 16497 25687
rect 16497 25653 16531 25687
rect 16531 25653 16540 25687
rect 16488 25644 16540 25653
rect 20076 25687 20128 25696
rect 20076 25653 20085 25687
rect 20085 25653 20119 25687
rect 20119 25653 20128 25687
rect 20076 25644 20128 25653
rect 22100 25644 22152 25696
rect 22376 25644 22428 25696
rect 22560 25687 22612 25696
rect 22560 25653 22569 25687
rect 22569 25653 22603 25687
rect 22603 25653 22612 25687
rect 22560 25644 22612 25653
rect 22652 25687 22704 25696
rect 22652 25653 22661 25687
rect 22661 25653 22695 25687
rect 22695 25653 22704 25687
rect 22652 25644 22704 25653
rect 23112 25644 23164 25696
rect 5170 25542 5222 25594
rect 5234 25542 5286 25594
rect 5298 25542 5350 25594
rect 5362 25542 5414 25594
rect 5426 25542 5478 25594
rect 13611 25542 13663 25594
rect 13675 25542 13727 25594
rect 13739 25542 13791 25594
rect 13803 25542 13855 25594
rect 13867 25542 13919 25594
rect 22052 25542 22104 25594
rect 22116 25542 22168 25594
rect 22180 25542 22232 25594
rect 22244 25542 22296 25594
rect 22308 25542 22360 25594
rect 30493 25542 30545 25594
rect 30557 25542 30609 25594
rect 30621 25542 30673 25594
rect 30685 25542 30737 25594
rect 30749 25542 30801 25594
rect 12072 25440 12124 25492
rect 12716 25440 12768 25492
rect 13360 25483 13412 25492
rect 13360 25449 13369 25483
rect 13369 25449 13403 25483
rect 13403 25449 13412 25483
rect 13360 25440 13412 25449
rect 13452 25440 13504 25492
rect 13728 25483 13780 25492
rect 13728 25449 13737 25483
rect 13737 25449 13771 25483
rect 13771 25449 13780 25483
rect 14832 25483 14884 25492
rect 13728 25440 13780 25449
rect 14832 25449 14841 25483
rect 14841 25449 14875 25483
rect 14875 25449 14884 25483
rect 14832 25440 14884 25449
rect 15200 25440 15252 25492
rect 10232 25372 10284 25424
rect 10140 25304 10192 25356
rect 11244 25304 11296 25356
rect 14556 25372 14608 25424
rect 15292 25372 15344 25424
rect 11888 25304 11940 25356
rect 11980 25304 12032 25356
rect 10600 25236 10652 25288
rect 11336 25236 11388 25288
rect 11428 25279 11480 25288
rect 11428 25245 11437 25279
rect 11437 25245 11471 25279
rect 11471 25245 11480 25279
rect 11428 25236 11480 25245
rect 12164 25279 12216 25288
rect 12164 25245 12173 25279
rect 12173 25245 12207 25279
rect 12207 25245 12216 25279
rect 12164 25236 12216 25245
rect 12256 25279 12308 25288
rect 12256 25245 12265 25279
rect 12265 25245 12299 25279
rect 12299 25245 12308 25279
rect 12256 25236 12308 25245
rect 12624 25236 12676 25288
rect 12900 25304 12952 25356
rect 10968 25168 11020 25220
rect 11980 25211 12032 25220
rect 11980 25177 11989 25211
rect 11989 25177 12023 25211
rect 12023 25177 12032 25211
rect 11980 25168 12032 25177
rect 13176 25236 13228 25288
rect 11520 25100 11572 25152
rect 13360 25100 13412 25152
rect 14188 25168 14240 25220
rect 14464 25211 14516 25220
rect 14464 25177 14473 25211
rect 14473 25177 14507 25211
rect 14507 25177 14516 25211
rect 14464 25168 14516 25177
rect 14924 25279 14976 25288
rect 14924 25245 14933 25279
rect 14933 25245 14967 25279
rect 14967 25245 14976 25279
rect 14924 25236 14976 25245
rect 15108 25236 15160 25288
rect 16580 25440 16632 25492
rect 17408 25440 17460 25492
rect 19708 25440 19760 25492
rect 20076 25440 20128 25492
rect 20904 25440 20956 25492
rect 22376 25440 22428 25492
rect 18788 25304 18840 25356
rect 19524 25304 19576 25356
rect 15660 25279 15712 25288
rect 15660 25245 15669 25279
rect 15669 25245 15703 25279
rect 15703 25245 15712 25279
rect 15660 25236 15712 25245
rect 16488 25279 16540 25288
rect 16488 25245 16522 25279
rect 16522 25245 16540 25279
rect 16488 25236 16540 25245
rect 14372 25100 14424 25152
rect 16120 25168 16172 25220
rect 19432 25279 19484 25288
rect 19432 25245 19436 25279
rect 19436 25245 19470 25279
rect 19470 25245 19484 25279
rect 19432 25236 19484 25245
rect 19616 25279 19668 25288
rect 19616 25245 19625 25279
rect 19625 25245 19659 25279
rect 19659 25245 19668 25279
rect 19616 25236 19668 25245
rect 21272 25372 21324 25424
rect 20168 25236 20220 25288
rect 21732 25304 21784 25356
rect 21916 25347 21968 25356
rect 21916 25313 21925 25347
rect 21925 25313 21959 25347
rect 21959 25313 21968 25347
rect 21916 25304 21968 25313
rect 22836 25347 22888 25356
rect 22836 25313 22845 25347
rect 22845 25313 22879 25347
rect 22879 25313 22888 25347
rect 22836 25304 22888 25313
rect 18604 25143 18656 25152
rect 18604 25109 18613 25143
rect 18613 25109 18647 25143
rect 18647 25109 18656 25143
rect 18604 25100 18656 25109
rect 19524 25211 19576 25220
rect 19524 25177 19533 25211
rect 19533 25177 19567 25211
rect 19567 25177 19576 25211
rect 19524 25168 19576 25177
rect 20444 25168 20496 25220
rect 21180 25236 21232 25288
rect 21640 25236 21692 25288
rect 23112 25279 23164 25288
rect 21824 25168 21876 25220
rect 22560 25168 22612 25220
rect 23112 25245 23146 25279
rect 23146 25245 23164 25279
rect 23112 25236 23164 25245
rect 24216 25236 24268 25288
rect 23020 25168 23072 25220
rect 20168 25100 20220 25152
rect 20720 25100 20772 25152
rect 20812 25100 20864 25152
rect 23848 25100 23900 25152
rect 24216 25143 24268 25152
rect 24216 25109 24225 25143
rect 24225 25109 24259 25143
rect 24259 25109 24268 25143
rect 24216 25100 24268 25109
rect 24860 25143 24912 25152
rect 24860 25109 24869 25143
rect 24869 25109 24903 25143
rect 24903 25109 24912 25143
rect 24860 25100 24912 25109
rect 9390 24998 9442 25050
rect 9454 24998 9506 25050
rect 9518 24998 9570 25050
rect 9582 24998 9634 25050
rect 9646 24998 9698 25050
rect 17831 24998 17883 25050
rect 17895 24998 17947 25050
rect 17959 24998 18011 25050
rect 18023 24998 18075 25050
rect 18087 24998 18139 25050
rect 26272 24998 26324 25050
rect 26336 24998 26388 25050
rect 26400 24998 26452 25050
rect 26464 24998 26516 25050
rect 26528 24998 26580 25050
rect 34713 24998 34765 25050
rect 34777 24998 34829 25050
rect 34841 24998 34893 25050
rect 34905 24998 34957 25050
rect 34969 24998 35021 25050
rect 10600 24896 10652 24948
rect 11060 24896 11112 24948
rect 11980 24896 12032 24948
rect 12164 24939 12216 24948
rect 12164 24905 12173 24939
rect 12173 24905 12207 24939
rect 12207 24905 12216 24939
rect 12164 24896 12216 24905
rect 12256 24896 12308 24948
rect 14924 24896 14976 24948
rect 17408 24939 17460 24948
rect 17408 24905 17417 24939
rect 17417 24905 17451 24939
rect 17451 24905 17460 24939
rect 17408 24896 17460 24905
rect 19524 24896 19576 24948
rect 10140 24760 10192 24812
rect 10232 24803 10284 24812
rect 10232 24769 10241 24803
rect 10241 24769 10275 24803
rect 10275 24769 10284 24803
rect 10232 24760 10284 24769
rect 10508 24760 10560 24812
rect 10600 24803 10652 24812
rect 10600 24769 10609 24803
rect 10609 24769 10643 24803
rect 10643 24769 10652 24803
rect 10600 24760 10652 24769
rect 10968 24803 11020 24812
rect 10968 24769 10977 24803
rect 10977 24769 11011 24803
rect 11011 24769 11020 24803
rect 10968 24760 11020 24769
rect 11060 24760 11112 24812
rect 11152 24760 11204 24812
rect 10048 24599 10100 24608
rect 10048 24565 10057 24599
rect 10057 24565 10091 24599
rect 10091 24565 10100 24599
rect 10048 24556 10100 24565
rect 11244 24692 11296 24744
rect 12992 24803 13044 24812
rect 12992 24769 13001 24803
rect 13001 24769 13035 24803
rect 13035 24769 13044 24803
rect 12992 24760 13044 24769
rect 13360 24760 13412 24812
rect 13728 24803 13780 24812
rect 13728 24769 13737 24803
rect 13737 24769 13771 24803
rect 13771 24769 13780 24803
rect 13728 24760 13780 24769
rect 14004 24760 14056 24812
rect 12532 24735 12584 24744
rect 12532 24701 12541 24735
rect 12541 24701 12575 24735
rect 12575 24701 12584 24735
rect 12532 24692 12584 24701
rect 13176 24692 13228 24744
rect 14188 24760 14240 24812
rect 14464 24828 14516 24880
rect 15108 24871 15160 24880
rect 14556 24803 14608 24812
rect 14556 24769 14565 24803
rect 14565 24769 14599 24803
rect 14599 24769 14608 24803
rect 14556 24760 14608 24769
rect 15108 24837 15117 24871
rect 15117 24837 15151 24871
rect 15151 24837 15160 24871
rect 15108 24828 15160 24837
rect 14832 24803 14884 24812
rect 14832 24769 14841 24803
rect 14841 24769 14875 24803
rect 14875 24769 14884 24803
rect 14832 24760 14884 24769
rect 15384 24692 15436 24744
rect 11336 24556 11388 24608
rect 11704 24599 11756 24608
rect 11704 24565 11713 24599
rect 11713 24565 11747 24599
rect 11747 24565 11756 24599
rect 11704 24556 11756 24565
rect 14096 24624 14148 24676
rect 14280 24624 14332 24676
rect 16120 24760 16172 24812
rect 17316 24760 17368 24812
rect 17592 24803 17644 24812
rect 17592 24769 17601 24803
rect 17601 24769 17635 24803
rect 17635 24769 17644 24803
rect 17592 24760 17644 24769
rect 19432 24871 19484 24880
rect 19432 24837 19441 24871
rect 19441 24837 19475 24871
rect 19475 24837 19484 24871
rect 19432 24828 19484 24837
rect 15660 24692 15712 24744
rect 15844 24735 15896 24744
rect 15844 24701 15853 24735
rect 15853 24701 15887 24735
rect 15887 24701 15896 24735
rect 15844 24692 15896 24701
rect 15936 24692 15988 24744
rect 18144 24803 18196 24812
rect 18144 24769 18153 24803
rect 18153 24769 18187 24803
rect 18187 24769 18196 24803
rect 18144 24760 18196 24769
rect 18236 24760 18288 24812
rect 20720 24896 20772 24948
rect 21548 24896 21600 24948
rect 22652 24896 22704 24948
rect 17040 24624 17092 24676
rect 19984 24803 20036 24812
rect 19984 24769 19993 24803
rect 19993 24769 20027 24803
rect 20027 24769 20036 24803
rect 19984 24760 20036 24769
rect 20260 24803 20312 24812
rect 20260 24769 20294 24803
rect 20294 24769 20312 24803
rect 20260 24760 20312 24769
rect 22468 24760 22520 24812
rect 21456 24692 21508 24744
rect 23020 24803 23072 24812
rect 23020 24769 23029 24803
rect 23029 24769 23063 24803
rect 23063 24769 23072 24803
rect 23020 24760 23072 24769
rect 24860 24760 24912 24812
rect 11888 24556 11940 24608
rect 15660 24599 15712 24608
rect 15660 24565 15669 24599
rect 15669 24565 15703 24599
rect 15703 24565 15712 24599
rect 15660 24556 15712 24565
rect 15752 24599 15804 24608
rect 15752 24565 15761 24599
rect 15761 24565 15795 24599
rect 15795 24565 15804 24599
rect 15752 24556 15804 24565
rect 18328 24556 18380 24608
rect 19524 24556 19576 24608
rect 19800 24599 19852 24608
rect 19800 24565 19809 24599
rect 19809 24565 19843 24599
rect 19843 24565 19852 24599
rect 19800 24556 19852 24565
rect 23756 24692 23808 24744
rect 22652 24624 22704 24676
rect 24216 24556 24268 24608
rect 5170 24454 5222 24506
rect 5234 24454 5286 24506
rect 5298 24454 5350 24506
rect 5362 24454 5414 24506
rect 5426 24454 5478 24506
rect 13611 24454 13663 24506
rect 13675 24454 13727 24506
rect 13739 24454 13791 24506
rect 13803 24454 13855 24506
rect 13867 24454 13919 24506
rect 22052 24454 22104 24506
rect 22116 24454 22168 24506
rect 22180 24454 22232 24506
rect 22244 24454 22296 24506
rect 22308 24454 22360 24506
rect 30493 24454 30545 24506
rect 30557 24454 30609 24506
rect 30621 24454 30673 24506
rect 30685 24454 30737 24506
rect 30749 24454 30801 24506
rect 10048 24352 10100 24404
rect 8944 24191 8996 24200
rect 8944 24157 8953 24191
rect 8953 24157 8987 24191
rect 8987 24157 8996 24191
rect 8944 24148 8996 24157
rect 10508 24284 10560 24336
rect 10692 24327 10744 24336
rect 10692 24293 10701 24327
rect 10701 24293 10735 24327
rect 10735 24293 10744 24327
rect 12532 24352 12584 24404
rect 13176 24352 13228 24404
rect 14004 24352 14056 24404
rect 14096 24352 14148 24404
rect 14832 24352 14884 24404
rect 15384 24352 15436 24404
rect 18144 24352 18196 24404
rect 20260 24352 20312 24404
rect 20996 24352 21048 24404
rect 22652 24352 22704 24404
rect 10692 24284 10744 24293
rect 14004 24216 14056 24268
rect 12716 24191 12768 24200
rect 12716 24157 12725 24191
rect 12725 24157 12759 24191
rect 12759 24157 12768 24191
rect 12716 24148 12768 24157
rect 12992 24148 13044 24200
rect 13452 24191 13504 24200
rect 13452 24157 13461 24191
rect 13461 24157 13495 24191
rect 13495 24157 13504 24191
rect 13452 24148 13504 24157
rect 14556 24284 14608 24336
rect 14372 24216 14424 24268
rect 9312 24080 9364 24132
rect 13728 24080 13780 24132
rect 14280 24191 14332 24200
rect 14280 24157 14289 24191
rect 14289 24157 14323 24191
rect 14323 24157 14332 24191
rect 14280 24148 14332 24157
rect 18604 24284 18656 24336
rect 19156 24284 19208 24336
rect 15292 24148 15344 24200
rect 17684 24148 17736 24200
rect 18696 24259 18748 24268
rect 18696 24225 18705 24259
rect 18705 24225 18739 24259
rect 18739 24225 18748 24259
rect 21732 24284 21784 24336
rect 22560 24284 22612 24336
rect 18696 24216 18748 24225
rect 19432 24216 19484 24268
rect 19616 24216 19668 24268
rect 21548 24259 21600 24268
rect 21548 24225 21557 24259
rect 21557 24225 21591 24259
rect 21591 24225 21600 24259
rect 21548 24216 21600 24225
rect 14464 24123 14516 24132
rect 14464 24089 14473 24123
rect 14473 24089 14507 24123
rect 14507 24089 14516 24123
rect 14464 24080 14516 24089
rect 17500 24080 17552 24132
rect 11244 24055 11296 24064
rect 11244 24021 11253 24055
rect 11253 24021 11287 24055
rect 11287 24021 11296 24055
rect 11244 24012 11296 24021
rect 12164 24055 12216 24064
rect 12164 24021 12173 24055
rect 12173 24021 12207 24055
rect 12207 24021 12216 24055
rect 12164 24012 12216 24021
rect 12900 24055 12952 24064
rect 12900 24021 12909 24055
rect 12909 24021 12943 24055
rect 12943 24021 12952 24055
rect 12900 24012 12952 24021
rect 13360 24012 13412 24064
rect 15476 24012 15528 24064
rect 15936 24055 15988 24064
rect 15936 24021 15945 24055
rect 15945 24021 15979 24055
rect 15979 24021 15988 24055
rect 15936 24012 15988 24021
rect 18236 24055 18288 24064
rect 18236 24021 18245 24055
rect 18245 24021 18279 24055
rect 18279 24021 18288 24055
rect 18236 24012 18288 24021
rect 21272 24191 21324 24200
rect 21272 24157 21281 24191
rect 21281 24157 21315 24191
rect 21315 24157 21324 24191
rect 21272 24148 21324 24157
rect 21824 24148 21876 24200
rect 23204 24191 23256 24200
rect 23204 24157 23213 24191
rect 23213 24157 23247 24191
rect 23247 24157 23256 24191
rect 23204 24148 23256 24157
rect 19432 24012 19484 24064
rect 22284 24012 22336 24064
rect 22928 24055 22980 24064
rect 22928 24021 22937 24055
rect 22937 24021 22971 24055
rect 22971 24021 22980 24055
rect 22928 24012 22980 24021
rect 23848 24055 23900 24064
rect 23848 24021 23857 24055
rect 23857 24021 23891 24055
rect 23891 24021 23900 24055
rect 23848 24012 23900 24021
rect 24492 24012 24544 24064
rect 24584 24012 24636 24064
rect 9390 23910 9442 23962
rect 9454 23910 9506 23962
rect 9518 23910 9570 23962
rect 9582 23910 9634 23962
rect 9646 23910 9698 23962
rect 17831 23910 17883 23962
rect 17895 23910 17947 23962
rect 17959 23910 18011 23962
rect 18023 23910 18075 23962
rect 18087 23910 18139 23962
rect 26272 23910 26324 23962
rect 26336 23910 26388 23962
rect 26400 23910 26452 23962
rect 26464 23910 26516 23962
rect 26528 23910 26580 23962
rect 34713 23910 34765 23962
rect 34777 23910 34829 23962
rect 34841 23910 34893 23962
rect 34905 23910 34957 23962
rect 34969 23910 35021 23962
rect 9312 23808 9364 23860
rect 11152 23808 11204 23860
rect 11244 23808 11296 23860
rect 11520 23808 11572 23860
rect 11704 23808 11756 23860
rect 12716 23808 12768 23860
rect 13452 23808 13504 23860
rect 13728 23808 13780 23860
rect 14280 23851 14332 23860
rect 14280 23817 14289 23851
rect 14289 23817 14323 23851
rect 14323 23817 14332 23851
rect 14280 23808 14332 23817
rect 14464 23808 14516 23860
rect 14648 23808 14700 23860
rect 14832 23808 14884 23860
rect 15660 23851 15712 23860
rect 15660 23817 15669 23851
rect 15669 23817 15703 23851
rect 15703 23817 15712 23851
rect 15660 23808 15712 23817
rect 15752 23808 15804 23860
rect 15844 23808 15896 23860
rect 10140 23647 10192 23656
rect 10140 23613 10149 23647
rect 10149 23613 10183 23647
rect 10183 23613 10192 23647
rect 10140 23604 10192 23613
rect 11520 23715 11572 23724
rect 11520 23681 11529 23715
rect 11529 23681 11563 23715
rect 11563 23681 11572 23715
rect 11520 23672 11572 23681
rect 11244 23647 11296 23656
rect 11244 23613 11253 23647
rect 11253 23613 11287 23647
rect 11287 23613 11296 23647
rect 11244 23604 11296 23613
rect 11888 23647 11940 23656
rect 11888 23613 11897 23647
rect 11897 23613 11931 23647
rect 11931 23613 11940 23647
rect 11888 23604 11940 23613
rect 12992 23672 13044 23724
rect 13176 23715 13228 23724
rect 13176 23681 13185 23715
rect 13185 23681 13219 23715
rect 13219 23681 13228 23715
rect 13176 23672 13228 23681
rect 13728 23672 13780 23724
rect 14188 23715 14240 23724
rect 14188 23681 14197 23715
rect 14197 23681 14231 23715
rect 14231 23681 14240 23715
rect 14188 23672 14240 23681
rect 14372 23672 14424 23724
rect 15292 23783 15344 23792
rect 15292 23749 15301 23783
rect 15301 23749 15335 23783
rect 15335 23749 15344 23783
rect 15292 23740 15344 23749
rect 14740 23715 14792 23724
rect 14740 23681 14749 23715
rect 14749 23681 14783 23715
rect 14783 23681 14792 23715
rect 14740 23672 14792 23681
rect 14924 23715 14976 23724
rect 14924 23681 14933 23715
rect 14933 23681 14967 23715
rect 14967 23681 14976 23715
rect 14924 23672 14976 23681
rect 15108 23672 15160 23724
rect 15568 23672 15620 23724
rect 16120 23808 16172 23860
rect 17500 23808 17552 23860
rect 18328 23808 18380 23860
rect 19616 23851 19668 23860
rect 19616 23817 19625 23851
rect 19625 23817 19659 23851
rect 19659 23817 19668 23851
rect 19616 23808 19668 23817
rect 19800 23808 19852 23860
rect 22376 23808 22428 23860
rect 22468 23808 22520 23860
rect 22928 23808 22980 23860
rect 23204 23808 23256 23860
rect 23848 23808 23900 23860
rect 17316 23672 17368 23724
rect 19616 23672 19668 23724
rect 20168 23672 20220 23724
rect 15384 23536 15436 23588
rect 11060 23468 11112 23520
rect 11888 23468 11940 23520
rect 13176 23468 13228 23520
rect 14464 23468 14516 23520
rect 14648 23468 14700 23520
rect 21640 23604 21692 23656
rect 22652 23715 22704 23724
rect 22652 23681 22661 23715
rect 22661 23681 22695 23715
rect 22695 23681 22704 23715
rect 22652 23672 22704 23681
rect 23664 23672 23716 23724
rect 24584 23672 24636 23724
rect 22468 23604 22520 23656
rect 22836 23604 22888 23656
rect 17684 23468 17736 23520
rect 18236 23468 18288 23520
rect 19708 23511 19760 23520
rect 19708 23477 19717 23511
rect 19717 23477 19751 23511
rect 19751 23477 19760 23511
rect 19708 23468 19760 23477
rect 19892 23468 19944 23520
rect 22560 23468 22612 23520
rect 24492 23511 24544 23520
rect 24492 23477 24501 23511
rect 24501 23477 24535 23511
rect 24535 23477 24544 23511
rect 24492 23468 24544 23477
rect 5170 23366 5222 23418
rect 5234 23366 5286 23418
rect 5298 23366 5350 23418
rect 5362 23366 5414 23418
rect 5426 23366 5478 23418
rect 13611 23366 13663 23418
rect 13675 23366 13727 23418
rect 13739 23366 13791 23418
rect 13803 23366 13855 23418
rect 13867 23366 13919 23418
rect 22052 23366 22104 23418
rect 22116 23366 22168 23418
rect 22180 23366 22232 23418
rect 22244 23366 22296 23418
rect 22308 23366 22360 23418
rect 30493 23366 30545 23418
rect 30557 23366 30609 23418
rect 30621 23366 30673 23418
rect 30685 23366 30737 23418
rect 30749 23366 30801 23418
rect 10600 23307 10652 23316
rect 10600 23273 10609 23307
rect 10609 23273 10643 23307
rect 10643 23273 10652 23307
rect 10600 23264 10652 23273
rect 11244 23264 11296 23316
rect 14188 23264 14240 23316
rect 14464 23307 14516 23316
rect 14464 23273 14473 23307
rect 14473 23273 14507 23307
rect 14507 23273 14516 23307
rect 14464 23264 14516 23273
rect 17316 23307 17368 23316
rect 17316 23273 17325 23307
rect 17325 23273 17359 23307
rect 17359 23273 17368 23307
rect 17316 23264 17368 23273
rect 19432 23307 19484 23316
rect 19432 23273 19441 23307
rect 19441 23273 19475 23307
rect 19475 23273 19484 23307
rect 19432 23264 19484 23273
rect 19524 23264 19576 23316
rect 22192 23264 22244 23316
rect 22468 23307 22520 23316
rect 22468 23273 22477 23307
rect 22477 23273 22511 23307
rect 22511 23273 22520 23307
rect 22468 23264 22520 23273
rect 22560 23264 22612 23316
rect 14096 23196 14148 23248
rect 15016 23196 15068 23248
rect 18144 23196 18196 23248
rect 21640 23196 21692 23248
rect 14740 23128 14792 23180
rect 18236 23171 18288 23180
rect 18236 23137 18245 23171
rect 18245 23137 18279 23171
rect 18279 23137 18288 23171
rect 18236 23128 18288 23137
rect 19616 23128 19668 23180
rect 21916 23171 21968 23180
rect 21916 23137 21925 23171
rect 21925 23137 21959 23171
rect 21959 23137 21968 23171
rect 21916 23128 21968 23137
rect 10692 23103 10744 23112
rect 10692 23069 10701 23103
rect 10701 23069 10735 23103
rect 10735 23069 10744 23103
rect 10692 23060 10744 23069
rect 12164 23103 12216 23112
rect 12164 23069 12182 23103
rect 12182 23069 12216 23103
rect 12164 23060 12216 23069
rect 12532 23103 12584 23112
rect 12532 23069 12541 23103
rect 12541 23069 12575 23103
rect 12575 23069 12584 23103
rect 12532 23060 12584 23069
rect 13544 23060 13596 23112
rect 14648 23103 14700 23112
rect 14648 23069 14657 23103
rect 14657 23069 14691 23103
rect 14691 23069 14700 23103
rect 14648 23060 14700 23069
rect 15292 23060 15344 23112
rect 16120 23060 16172 23112
rect 17040 23060 17092 23112
rect 12900 22992 12952 23044
rect 17408 23060 17460 23112
rect 19064 23103 19116 23112
rect 19064 23069 19073 23103
rect 19073 23069 19107 23103
rect 19107 23069 19116 23103
rect 19064 23060 19116 23069
rect 19156 23060 19208 23112
rect 20536 23103 20588 23112
rect 20536 23069 20545 23103
rect 20545 23069 20579 23103
rect 20579 23069 20588 23103
rect 20536 23060 20588 23069
rect 21364 23103 21416 23112
rect 21364 23069 21373 23103
rect 21373 23069 21407 23103
rect 21407 23069 21416 23103
rect 21364 23060 21416 23069
rect 21548 23060 21600 23112
rect 21824 23103 21876 23112
rect 21824 23069 21833 23103
rect 21833 23069 21867 23103
rect 21867 23069 21876 23103
rect 21824 23060 21876 23069
rect 22008 23103 22060 23112
rect 22008 23069 22017 23103
rect 22017 23069 22051 23103
rect 22051 23069 22060 23103
rect 22008 23060 22060 23069
rect 15568 22967 15620 22976
rect 15568 22933 15577 22967
rect 15577 22933 15611 22967
rect 15611 22933 15620 22967
rect 15568 22924 15620 22933
rect 18236 22924 18288 22976
rect 19892 22924 19944 22976
rect 21640 22967 21692 22976
rect 21640 22933 21649 22967
rect 21649 22933 21683 22967
rect 21683 22933 21692 22967
rect 21640 22924 21692 22933
rect 21916 22992 21968 23044
rect 23020 23128 23072 23180
rect 22468 23060 22520 23112
rect 22928 23103 22980 23112
rect 22928 23069 22937 23103
rect 22937 23069 22971 23103
rect 22971 23069 22980 23103
rect 22928 23060 22980 23069
rect 23848 23035 23900 23044
rect 23848 23001 23857 23035
rect 23857 23001 23891 23035
rect 23891 23001 23900 23035
rect 23848 22992 23900 23001
rect 22284 22924 22336 22976
rect 22560 22924 22612 22976
rect 23296 22924 23348 22976
rect 24400 23128 24452 23180
rect 24124 22924 24176 22976
rect 24216 22924 24268 22976
rect 24308 22924 24360 22976
rect 9390 22822 9442 22874
rect 9454 22822 9506 22874
rect 9518 22822 9570 22874
rect 9582 22822 9634 22874
rect 9646 22822 9698 22874
rect 17831 22822 17883 22874
rect 17895 22822 17947 22874
rect 17959 22822 18011 22874
rect 18023 22822 18075 22874
rect 18087 22822 18139 22874
rect 26272 22822 26324 22874
rect 26336 22822 26388 22874
rect 26400 22822 26452 22874
rect 26464 22822 26516 22874
rect 26528 22822 26580 22874
rect 34713 22822 34765 22874
rect 34777 22822 34829 22874
rect 34841 22822 34893 22874
rect 34905 22822 34957 22874
rect 34969 22822 35021 22874
rect 11244 22720 11296 22772
rect 9036 22652 9088 22704
rect 9864 22627 9916 22636
rect 9864 22593 9873 22627
rect 9873 22593 9907 22627
rect 9907 22593 9916 22627
rect 9864 22584 9916 22593
rect 12808 22584 12860 22636
rect 13084 22584 13136 22636
rect 14188 22720 14240 22772
rect 14556 22720 14608 22772
rect 13452 22652 13504 22704
rect 14096 22627 14148 22636
rect 14096 22593 14105 22627
rect 14105 22593 14139 22627
rect 14139 22593 14148 22627
rect 14096 22584 14148 22593
rect 15476 22720 15528 22772
rect 15568 22720 15620 22772
rect 16120 22763 16172 22772
rect 16120 22729 16129 22763
rect 16129 22729 16163 22763
rect 16163 22729 16172 22763
rect 16120 22720 16172 22729
rect 19708 22720 19760 22772
rect 22008 22720 22060 22772
rect 22192 22720 22244 22772
rect 14832 22584 14884 22636
rect 16488 22627 16540 22636
rect 16488 22593 16497 22627
rect 16497 22593 16531 22627
rect 16531 22593 16540 22627
rect 16488 22584 16540 22593
rect 16672 22584 16724 22636
rect 17408 22584 17460 22636
rect 18236 22584 18288 22636
rect 10784 22559 10836 22568
rect 10784 22525 10793 22559
rect 10793 22525 10827 22559
rect 10827 22525 10836 22559
rect 10784 22516 10836 22525
rect 11520 22516 11572 22568
rect 13544 22516 13596 22568
rect 13176 22448 13228 22500
rect 9864 22423 9916 22432
rect 9864 22389 9873 22423
rect 9873 22389 9907 22423
rect 9907 22389 9916 22423
rect 9864 22380 9916 22389
rect 10232 22423 10284 22432
rect 10232 22389 10241 22423
rect 10241 22389 10275 22423
rect 10275 22389 10284 22423
rect 10232 22380 10284 22389
rect 11152 22423 11204 22432
rect 11152 22389 11161 22423
rect 11161 22389 11195 22423
rect 11195 22389 11204 22423
rect 11152 22380 11204 22389
rect 12440 22380 12492 22432
rect 13268 22423 13320 22432
rect 13268 22389 13277 22423
rect 13277 22389 13311 22423
rect 13311 22389 13320 22423
rect 13268 22380 13320 22389
rect 13360 22380 13412 22432
rect 14648 22448 14700 22500
rect 17132 22559 17184 22568
rect 17132 22525 17141 22559
rect 17141 22525 17175 22559
rect 17175 22525 17184 22559
rect 17132 22516 17184 22525
rect 19616 22627 19668 22636
rect 19616 22593 19625 22627
rect 19625 22593 19659 22627
rect 19659 22593 19668 22627
rect 19616 22584 19668 22593
rect 19892 22584 19944 22636
rect 20260 22584 20312 22636
rect 20168 22516 20220 22568
rect 14280 22423 14332 22432
rect 14280 22389 14289 22423
rect 14289 22389 14323 22423
rect 14323 22389 14332 22423
rect 14280 22380 14332 22389
rect 15108 22380 15160 22432
rect 16120 22380 16172 22432
rect 16396 22423 16448 22432
rect 16396 22389 16405 22423
rect 16405 22389 16439 22423
rect 16439 22389 16448 22423
rect 16396 22380 16448 22389
rect 17500 22380 17552 22432
rect 17960 22423 18012 22432
rect 17960 22389 17969 22423
rect 17969 22389 18003 22423
rect 18003 22389 18012 22423
rect 17960 22380 18012 22389
rect 19432 22448 19484 22500
rect 19616 22380 19668 22432
rect 20352 22380 20404 22432
rect 21364 22584 21416 22636
rect 21548 22584 21600 22636
rect 21732 22584 21784 22636
rect 22560 22720 22612 22772
rect 22928 22720 22980 22772
rect 22468 22652 22520 22704
rect 23296 22652 23348 22704
rect 24400 22763 24452 22772
rect 24400 22729 24409 22763
rect 24409 22729 24443 22763
rect 24443 22729 24452 22763
rect 24400 22720 24452 22729
rect 22100 22448 22152 22500
rect 22376 22559 22428 22568
rect 22376 22525 22385 22559
rect 22385 22525 22419 22559
rect 22419 22525 22428 22559
rect 22376 22516 22428 22525
rect 23572 22584 23624 22636
rect 24124 22584 24176 22636
rect 22836 22559 22888 22568
rect 22836 22525 22845 22559
rect 22845 22525 22879 22559
rect 22879 22525 22888 22559
rect 22836 22516 22888 22525
rect 24216 22423 24268 22432
rect 24216 22389 24225 22423
rect 24225 22389 24259 22423
rect 24259 22389 24268 22423
rect 24216 22380 24268 22389
rect 5170 22278 5222 22330
rect 5234 22278 5286 22330
rect 5298 22278 5350 22330
rect 5362 22278 5414 22330
rect 5426 22278 5478 22330
rect 13611 22278 13663 22330
rect 13675 22278 13727 22330
rect 13739 22278 13791 22330
rect 13803 22278 13855 22330
rect 13867 22278 13919 22330
rect 22052 22278 22104 22330
rect 22116 22278 22168 22330
rect 22180 22278 22232 22330
rect 22244 22278 22296 22330
rect 22308 22278 22360 22330
rect 30493 22278 30545 22330
rect 30557 22278 30609 22330
rect 30621 22278 30673 22330
rect 30685 22278 30737 22330
rect 30749 22278 30801 22330
rect 13084 22176 13136 22228
rect 16120 22176 16172 22228
rect 8944 22083 8996 22092
rect 8944 22049 8953 22083
rect 8953 22049 8987 22083
rect 8987 22049 8996 22083
rect 8944 22040 8996 22049
rect 10784 22108 10836 22160
rect 12440 22108 12492 22160
rect 14372 22108 14424 22160
rect 11980 22040 12032 22092
rect 940 21904 992 21956
rect 9312 21904 9364 21956
rect 10968 22015 11020 22024
rect 10968 21981 10977 22015
rect 10977 21981 11011 22015
rect 11011 21981 11020 22015
rect 10968 21972 11020 21981
rect 11152 21972 11204 22024
rect 11244 22015 11296 22024
rect 11244 21981 11253 22015
rect 11253 21981 11287 22015
rect 11287 21981 11296 22015
rect 11244 21972 11296 21981
rect 11520 22015 11572 22024
rect 11520 21981 11529 22015
rect 11529 21981 11563 22015
rect 11563 21981 11572 22015
rect 11520 21972 11572 21981
rect 12072 22015 12124 22024
rect 12072 21981 12081 22015
rect 12081 21981 12115 22015
rect 12115 21981 12124 22015
rect 12072 21972 12124 21981
rect 12624 22015 12676 22024
rect 12624 21981 12633 22015
rect 12633 21981 12667 22015
rect 12667 21981 12676 22015
rect 12624 21972 12676 21981
rect 13268 22040 13320 22092
rect 13820 21972 13872 22024
rect 14188 21972 14240 22024
rect 15292 22108 15344 22160
rect 14648 22015 14700 22024
rect 14648 21981 14656 22015
rect 14656 21981 14690 22015
rect 14690 21981 14700 22015
rect 14648 21972 14700 21981
rect 14740 22015 14792 22024
rect 14740 21981 14749 22015
rect 14749 21981 14783 22015
rect 14783 21981 14792 22015
rect 14740 21972 14792 21981
rect 15108 22015 15160 22024
rect 15108 21981 15117 22015
rect 15117 21981 15151 22015
rect 15151 21981 15160 22015
rect 15108 21972 15160 21981
rect 15200 22015 15252 22024
rect 15200 21981 15209 22015
rect 15209 21981 15243 22015
rect 15243 21981 15252 22015
rect 15200 21972 15252 21981
rect 15844 21972 15896 22024
rect 11888 21879 11940 21888
rect 11888 21845 11897 21879
rect 11897 21845 11931 21879
rect 11931 21845 11940 21879
rect 11888 21836 11940 21845
rect 12348 21836 12400 21888
rect 12716 21836 12768 21888
rect 12992 21879 13044 21888
rect 12992 21845 13001 21879
rect 13001 21845 13035 21879
rect 13035 21845 13044 21879
rect 12992 21836 13044 21845
rect 13728 21879 13780 21888
rect 13728 21845 13737 21879
rect 13737 21845 13771 21879
rect 13771 21845 13780 21879
rect 13728 21836 13780 21845
rect 14004 21836 14056 21888
rect 14096 21879 14148 21888
rect 14096 21845 14105 21879
rect 14105 21845 14139 21879
rect 14139 21845 14148 21879
rect 14096 21836 14148 21845
rect 14832 21836 14884 21888
rect 15384 21879 15436 21888
rect 15384 21845 15393 21879
rect 15393 21845 15427 21879
rect 15427 21845 15436 21879
rect 15384 21836 15436 21845
rect 17408 21972 17460 22024
rect 17684 22015 17736 22024
rect 17684 21981 17693 22015
rect 17693 21981 17727 22015
rect 17727 21981 17736 22015
rect 17684 21972 17736 21981
rect 17960 22015 18012 22024
rect 17960 21981 17994 22015
rect 17994 21981 18012 22015
rect 17960 21972 18012 21981
rect 18420 21972 18472 22024
rect 20812 22219 20864 22228
rect 20812 22185 20821 22219
rect 20821 22185 20855 22219
rect 20855 22185 20864 22219
rect 20812 22176 20864 22185
rect 21364 22176 21416 22228
rect 21916 22176 21968 22228
rect 20076 22040 20128 22092
rect 21548 22108 21600 22160
rect 23664 22176 23716 22228
rect 21916 22040 21968 22092
rect 24308 22040 24360 22092
rect 19432 21972 19484 22024
rect 20168 21972 20220 22024
rect 20260 22015 20312 22024
rect 20260 21981 20268 22015
rect 20268 21981 20302 22015
rect 20302 21981 20312 22015
rect 20260 21972 20312 21981
rect 20352 22015 20404 22024
rect 20352 21981 20361 22015
rect 20361 21981 20395 22015
rect 20395 21981 20404 22015
rect 20352 21972 20404 21981
rect 16764 21879 16816 21888
rect 16764 21845 16773 21879
rect 16773 21845 16807 21879
rect 16807 21845 16816 21879
rect 16764 21836 16816 21845
rect 17316 21836 17368 21888
rect 18788 21836 18840 21888
rect 19248 21879 19300 21888
rect 19248 21845 19257 21879
rect 19257 21845 19291 21879
rect 19291 21845 19300 21879
rect 19248 21836 19300 21845
rect 19616 21947 19668 21956
rect 19616 21913 19625 21947
rect 19625 21913 19659 21947
rect 19659 21913 19668 21947
rect 19616 21904 19668 21913
rect 19432 21879 19484 21888
rect 19432 21845 19454 21879
rect 19454 21845 19484 21879
rect 19432 21836 19484 21845
rect 19892 21836 19944 21888
rect 20904 21972 20956 22024
rect 20996 22015 21048 22024
rect 20996 21981 21005 22015
rect 21005 21981 21039 22015
rect 21039 21981 21048 22015
rect 20996 21972 21048 21981
rect 22468 21972 22520 22024
rect 23572 22015 23624 22024
rect 23572 21981 23581 22015
rect 23581 21981 23615 22015
rect 23615 21981 23624 22015
rect 23572 21972 23624 21981
rect 21272 21879 21324 21888
rect 21272 21845 21281 21879
rect 21281 21845 21315 21879
rect 21315 21845 21324 21879
rect 21272 21836 21324 21845
rect 9390 21734 9442 21786
rect 9454 21734 9506 21786
rect 9518 21734 9570 21786
rect 9582 21734 9634 21786
rect 9646 21734 9698 21786
rect 17831 21734 17883 21786
rect 17895 21734 17947 21786
rect 17959 21734 18011 21786
rect 18023 21734 18075 21786
rect 18087 21734 18139 21786
rect 26272 21734 26324 21786
rect 26336 21734 26388 21786
rect 26400 21734 26452 21786
rect 26464 21734 26516 21786
rect 26528 21734 26580 21786
rect 34713 21734 34765 21786
rect 34777 21734 34829 21786
rect 34841 21734 34893 21786
rect 34905 21734 34957 21786
rect 34969 21734 35021 21786
rect 9312 21632 9364 21684
rect 10968 21632 11020 21684
rect 11152 21632 11204 21684
rect 10232 21564 10284 21616
rect 9864 21496 9916 21548
rect 10692 21496 10744 21548
rect 10784 21539 10836 21548
rect 10784 21505 10793 21539
rect 10793 21505 10827 21539
rect 10827 21505 10836 21539
rect 10784 21496 10836 21505
rect 10968 21539 11020 21548
rect 10968 21505 10977 21539
rect 10977 21505 11011 21539
rect 11011 21505 11020 21539
rect 10968 21496 11020 21505
rect 11888 21632 11940 21684
rect 12624 21632 12676 21684
rect 12992 21632 13044 21684
rect 11888 21539 11940 21548
rect 11888 21505 11897 21539
rect 11897 21505 11931 21539
rect 11931 21505 11940 21539
rect 11888 21496 11940 21505
rect 12072 21539 12124 21548
rect 12072 21505 12080 21539
rect 12080 21505 12114 21539
rect 12114 21505 12124 21539
rect 12072 21496 12124 21505
rect 12440 21496 12492 21548
rect 12624 21539 12676 21548
rect 12624 21505 12633 21539
rect 12633 21505 12667 21539
rect 12667 21505 12676 21539
rect 12624 21496 12676 21505
rect 13728 21632 13780 21684
rect 14096 21564 14148 21616
rect 15108 21675 15160 21684
rect 15108 21641 15117 21675
rect 15117 21641 15151 21675
rect 15151 21641 15160 21675
rect 15108 21632 15160 21641
rect 15476 21632 15528 21684
rect 16488 21632 16540 21684
rect 16764 21632 16816 21684
rect 17316 21632 17368 21684
rect 17408 21632 17460 21684
rect 18420 21675 18472 21684
rect 18420 21641 18429 21675
rect 18429 21641 18463 21675
rect 18463 21641 18472 21675
rect 18420 21632 18472 21641
rect 13268 21539 13320 21548
rect 13268 21505 13277 21539
rect 13277 21505 13311 21539
rect 13311 21505 13320 21539
rect 13268 21496 13320 21505
rect 13544 21539 13596 21548
rect 13544 21505 13559 21539
rect 13559 21505 13593 21539
rect 13593 21505 13596 21539
rect 13544 21496 13596 21505
rect 13452 21471 13504 21480
rect 13452 21437 13461 21471
rect 13461 21437 13495 21471
rect 13495 21437 13504 21471
rect 13452 21428 13504 21437
rect 14188 21428 14240 21480
rect 14924 21539 14976 21548
rect 14924 21505 14933 21539
rect 14933 21505 14967 21539
rect 14967 21505 14976 21539
rect 14924 21496 14976 21505
rect 15016 21496 15068 21548
rect 15200 21539 15252 21548
rect 15200 21505 15209 21539
rect 15209 21505 15243 21539
rect 15243 21505 15252 21539
rect 15200 21496 15252 21505
rect 16672 21496 16724 21548
rect 17500 21496 17552 21548
rect 19432 21632 19484 21684
rect 20168 21632 20220 21684
rect 20812 21632 20864 21684
rect 21824 21632 21876 21684
rect 22468 21632 22520 21684
rect 15660 21428 15712 21480
rect 9036 21335 9088 21344
rect 9036 21301 9045 21335
rect 9045 21301 9079 21335
rect 9079 21301 9088 21335
rect 9036 21292 9088 21301
rect 9220 21292 9272 21344
rect 9956 21292 10008 21344
rect 14464 21360 14516 21412
rect 16948 21471 17000 21480
rect 16948 21437 16957 21471
rect 16957 21437 16991 21471
rect 16991 21437 17000 21471
rect 16948 21428 17000 21437
rect 21088 21564 21140 21616
rect 21548 21564 21600 21616
rect 19892 21539 19944 21548
rect 19892 21505 19901 21539
rect 19901 21505 19935 21539
rect 19935 21505 19944 21539
rect 19892 21496 19944 21505
rect 20076 21539 20128 21548
rect 20076 21505 20085 21539
rect 20085 21505 20119 21539
rect 20119 21505 20128 21539
rect 20076 21496 20128 21505
rect 18420 21360 18472 21412
rect 20352 21428 20404 21480
rect 21272 21496 21324 21548
rect 21824 21539 21876 21548
rect 21824 21505 21833 21539
rect 21833 21505 21867 21539
rect 21867 21505 21876 21539
rect 21824 21496 21876 21505
rect 20720 21428 20772 21480
rect 22652 21539 22704 21548
rect 22652 21505 22661 21539
rect 22661 21505 22695 21539
rect 22695 21505 22704 21539
rect 22652 21496 22704 21505
rect 23480 21471 23532 21480
rect 23480 21437 23489 21471
rect 23489 21437 23523 21471
rect 23523 21437 23532 21471
rect 23480 21428 23532 21437
rect 13084 21335 13136 21344
rect 13084 21301 13093 21335
rect 13093 21301 13127 21335
rect 13127 21301 13136 21335
rect 13084 21292 13136 21301
rect 13176 21292 13228 21344
rect 14740 21335 14792 21344
rect 14740 21301 14749 21335
rect 14749 21301 14783 21335
rect 14783 21301 14792 21335
rect 14740 21292 14792 21301
rect 15108 21292 15160 21344
rect 15752 21292 15804 21344
rect 16488 21335 16540 21344
rect 16488 21301 16497 21335
rect 16497 21301 16531 21335
rect 16531 21301 16540 21335
rect 16488 21292 16540 21301
rect 20628 21335 20680 21344
rect 20628 21301 20637 21335
rect 20637 21301 20671 21335
rect 20671 21301 20680 21335
rect 20628 21292 20680 21301
rect 20812 21335 20864 21344
rect 20812 21301 20821 21335
rect 20821 21301 20855 21335
rect 20855 21301 20864 21335
rect 20812 21292 20864 21301
rect 20904 21292 20956 21344
rect 21732 21292 21784 21344
rect 22376 21292 22428 21344
rect 22560 21292 22612 21344
rect 5170 21190 5222 21242
rect 5234 21190 5286 21242
rect 5298 21190 5350 21242
rect 5362 21190 5414 21242
rect 5426 21190 5478 21242
rect 13611 21190 13663 21242
rect 13675 21190 13727 21242
rect 13739 21190 13791 21242
rect 13803 21190 13855 21242
rect 13867 21190 13919 21242
rect 22052 21190 22104 21242
rect 22116 21190 22168 21242
rect 22180 21190 22232 21242
rect 22244 21190 22296 21242
rect 22308 21190 22360 21242
rect 30493 21190 30545 21242
rect 30557 21190 30609 21242
rect 30621 21190 30673 21242
rect 30685 21190 30737 21242
rect 30749 21190 30801 21242
rect 9772 21088 9824 21140
rect 13084 21088 13136 21140
rect 13176 21088 13228 21140
rect 13452 21088 13504 21140
rect 14188 21088 14240 21140
rect 10968 20952 11020 21004
rect 8484 20927 8536 20936
rect 8484 20893 8493 20927
rect 8493 20893 8527 20927
rect 8527 20893 8536 20927
rect 8484 20884 8536 20893
rect 9312 20748 9364 20800
rect 10416 20927 10468 20936
rect 10416 20893 10425 20927
rect 10425 20893 10459 20927
rect 10459 20893 10468 20927
rect 10416 20884 10468 20893
rect 14096 21020 14148 21072
rect 14464 21063 14516 21072
rect 14464 21029 14473 21063
rect 14473 21029 14507 21063
rect 14507 21029 14516 21063
rect 14464 21020 14516 21029
rect 14740 21088 14792 21140
rect 14832 21088 14884 21140
rect 15200 21020 15252 21072
rect 12808 20927 12860 20936
rect 12808 20893 12817 20927
rect 12817 20893 12851 20927
rect 12851 20893 12860 20927
rect 12808 20884 12860 20893
rect 12532 20816 12584 20868
rect 13820 20884 13872 20936
rect 14280 20952 14332 21004
rect 15476 21088 15528 21140
rect 15660 21131 15712 21140
rect 15660 21097 15669 21131
rect 15669 21097 15703 21131
rect 15703 21097 15712 21131
rect 15660 21088 15712 21097
rect 15752 21088 15804 21140
rect 15384 21020 15436 21072
rect 15844 21020 15896 21072
rect 17500 21020 17552 21072
rect 18696 21063 18748 21072
rect 18696 21029 18705 21063
rect 18705 21029 18739 21063
rect 18739 21029 18748 21063
rect 18696 21020 18748 21029
rect 11060 20748 11112 20800
rect 11704 20791 11756 20800
rect 11704 20757 11713 20791
rect 11713 20757 11747 20791
rect 11747 20757 11756 20791
rect 11704 20748 11756 20757
rect 12256 20791 12308 20800
rect 12256 20757 12265 20791
rect 12265 20757 12299 20791
rect 12299 20757 12308 20791
rect 12256 20748 12308 20757
rect 12348 20748 12400 20800
rect 12992 20748 13044 20800
rect 14096 20748 14148 20800
rect 15384 20816 15436 20868
rect 15660 20816 15712 20868
rect 20444 21088 20496 21140
rect 20628 21088 20680 21140
rect 22284 21088 22336 21140
rect 22560 21088 22612 21140
rect 23480 21088 23532 21140
rect 20168 21020 20220 21072
rect 21732 21020 21784 21072
rect 16488 20884 16540 20936
rect 16948 20884 17000 20936
rect 17684 20884 17736 20936
rect 16672 20816 16724 20868
rect 20076 20927 20128 20936
rect 20076 20893 20085 20927
rect 20085 20893 20119 20927
rect 20119 20893 20128 20927
rect 20076 20884 20128 20893
rect 20352 20884 20404 20936
rect 20720 20927 20772 20936
rect 20720 20893 20729 20927
rect 20729 20893 20763 20927
rect 20763 20893 20772 20927
rect 20720 20884 20772 20893
rect 21548 20927 21600 20936
rect 21548 20893 21557 20927
rect 21557 20893 21591 20927
rect 21591 20893 21600 20927
rect 21548 20884 21600 20893
rect 21732 20927 21784 20936
rect 21732 20893 21741 20927
rect 21741 20893 21775 20927
rect 21775 20893 21784 20927
rect 21732 20884 21784 20893
rect 18788 20816 18840 20868
rect 22284 20884 22336 20936
rect 22376 20927 22428 20936
rect 22376 20893 22385 20927
rect 22385 20893 22419 20927
rect 22419 20893 22428 20927
rect 22376 20884 22428 20893
rect 18880 20791 18932 20800
rect 18880 20757 18889 20791
rect 18889 20757 18923 20791
rect 18923 20757 18932 20791
rect 18880 20748 18932 20757
rect 22284 20791 22336 20800
rect 22284 20757 22293 20791
rect 22293 20757 22327 20791
rect 22327 20757 22336 20791
rect 22284 20748 22336 20757
rect 22744 20816 22796 20868
rect 22836 20816 22888 20868
rect 23572 20748 23624 20800
rect 9390 20646 9442 20698
rect 9454 20646 9506 20698
rect 9518 20646 9570 20698
rect 9582 20646 9634 20698
rect 9646 20646 9698 20698
rect 17831 20646 17883 20698
rect 17895 20646 17947 20698
rect 17959 20646 18011 20698
rect 18023 20646 18075 20698
rect 18087 20646 18139 20698
rect 26272 20646 26324 20698
rect 26336 20646 26388 20698
rect 26400 20646 26452 20698
rect 26464 20646 26516 20698
rect 26528 20646 26580 20698
rect 34713 20646 34765 20698
rect 34777 20646 34829 20698
rect 34841 20646 34893 20698
rect 34905 20646 34957 20698
rect 34969 20646 35021 20698
rect 8484 20544 8536 20596
rect 9220 20544 9272 20596
rect 10968 20544 11020 20596
rect 11060 20544 11112 20596
rect 8944 20408 8996 20460
rect 9312 20476 9364 20528
rect 13452 20544 13504 20596
rect 14188 20587 14240 20596
rect 14188 20553 14197 20587
rect 14197 20553 14231 20587
rect 14231 20553 14240 20587
rect 14188 20544 14240 20553
rect 14924 20544 14976 20596
rect 15200 20544 15252 20596
rect 15384 20544 15436 20596
rect 16396 20544 16448 20596
rect 9956 20408 10008 20460
rect 10048 20408 10100 20460
rect 12348 20476 12400 20528
rect 19340 20476 19392 20528
rect 12256 20408 12308 20460
rect 12532 20408 12584 20460
rect 13084 20451 13136 20460
rect 13084 20417 13118 20451
rect 13118 20417 13136 20451
rect 13084 20408 13136 20417
rect 17132 20408 17184 20460
rect 20076 20451 20128 20460
rect 20076 20417 20085 20451
rect 20085 20417 20119 20451
rect 20119 20417 20128 20451
rect 20076 20408 20128 20417
rect 20720 20544 20772 20596
rect 21180 20544 21232 20596
rect 9312 20383 9364 20392
rect 9312 20349 9321 20383
rect 9321 20349 9355 20383
rect 9355 20349 9364 20383
rect 9312 20340 9364 20349
rect 14372 20383 14424 20392
rect 14372 20349 14381 20383
rect 14381 20349 14415 20383
rect 14415 20349 14424 20383
rect 14372 20340 14424 20349
rect 9220 20204 9272 20256
rect 11060 20204 11112 20256
rect 13820 20272 13872 20324
rect 14556 20272 14608 20324
rect 17224 20383 17276 20392
rect 17224 20349 17233 20383
rect 17233 20349 17267 20383
rect 17267 20349 17276 20383
rect 17224 20340 17276 20349
rect 20812 20476 20864 20528
rect 12440 20204 12492 20256
rect 12716 20247 12768 20256
rect 12716 20213 12725 20247
rect 12725 20213 12759 20247
rect 12759 20213 12768 20247
rect 12716 20204 12768 20213
rect 15016 20247 15068 20256
rect 15016 20213 15025 20247
rect 15025 20213 15059 20247
rect 15059 20213 15068 20247
rect 15016 20204 15068 20213
rect 17776 20204 17828 20256
rect 20260 20247 20312 20256
rect 20260 20213 20269 20247
rect 20269 20213 20303 20247
rect 20303 20213 20312 20247
rect 20260 20204 20312 20213
rect 20536 20247 20588 20256
rect 20536 20213 20545 20247
rect 20545 20213 20579 20247
rect 20579 20213 20588 20247
rect 20536 20204 20588 20213
rect 21824 20408 21876 20460
rect 22192 20408 22244 20460
rect 22284 20408 22336 20460
rect 21916 20383 21968 20392
rect 21916 20349 21925 20383
rect 21925 20349 21959 20383
rect 21959 20349 21968 20383
rect 21916 20340 21968 20349
rect 22744 20476 22796 20528
rect 23572 20519 23624 20528
rect 23572 20485 23581 20519
rect 23581 20485 23615 20519
rect 23615 20485 23624 20519
rect 23572 20476 23624 20485
rect 23204 20451 23256 20460
rect 23204 20417 23213 20451
rect 23213 20417 23247 20451
rect 23247 20417 23256 20451
rect 23204 20408 23256 20417
rect 20812 20272 20864 20324
rect 21548 20272 21600 20324
rect 21916 20204 21968 20256
rect 22468 20204 22520 20256
rect 33140 20204 33192 20256
rect 5170 20102 5222 20154
rect 5234 20102 5286 20154
rect 5298 20102 5350 20154
rect 5362 20102 5414 20154
rect 5426 20102 5478 20154
rect 13611 20102 13663 20154
rect 13675 20102 13727 20154
rect 13739 20102 13791 20154
rect 13803 20102 13855 20154
rect 13867 20102 13919 20154
rect 22052 20102 22104 20154
rect 22116 20102 22168 20154
rect 22180 20102 22232 20154
rect 22244 20102 22296 20154
rect 22308 20102 22360 20154
rect 30493 20102 30545 20154
rect 30557 20102 30609 20154
rect 30621 20102 30673 20154
rect 30685 20102 30737 20154
rect 30749 20102 30801 20154
rect 10048 20000 10100 20052
rect 9312 19864 9364 19916
rect 11704 20000 11756 20052
rect 11888 19932 11940 19984
rect 13084 20000 13136 20052
rect 14556 20000 14608 20052
rect 9772 19839 9824 19848
rect 9772 19805 9781 19839
rect 9781 19805 9815 19839
rect 9815 19805 9824 19839
rect 9772 19796 9824 19805
rect 10692 19796 10744 19848
rect 12716 19839 12768 19848
rect 12716 19805 12734 19839
rect 12734 19805 12768 19839
rect 12716 19796 12768 19805
rect 13176 19796 13228 19848
rect 13268 19839 13320 19848
rect 13268 19805 13277 19839
rect 13277 19805 13311 19839
rect 13311 19805 13320 19839
rect 13268 19796 13320 19805
rect 15016 19796 15068 19848
rect 15292 20000 15344 20052
rect 15660 20043 15712 20052
rect 15660 20009 15669 20043
rect 15669 20009 15703 20043
rect 15703 20009 15712 20043
rect 15660 20000 15712 20009
rect 17224 20000 17276 20052
rect 19616 20000 19668 20052
rect 20352 20000 20404 20052
rect 20536 20000 20588 20052
rect 20812 20043 20864 20052
rect 20812 20009 20821 20043
rect 20821 20009 20855 20043
rect 20855 20009 20864 20043
rect 20812 20000 20864 20009
rect 20996 20000 21048 20052
rect 21732 20043 21784 20052
rect 21732 20009 21741 20043
rect 21741 20009 21775 20043
rect 21775 20009 21784 20043
rect 21732 20000 21784 20009
rect 22468 20000 22520 20052
rect 22652 20043 22704 20052
rect 22652 20009 22661 20043
rect 22661 20009 22695 20043
rect 22695 20009 22704 20043
rect 22652 20000 22704 20009
rect 23204 20000 23256 20052
rect 16396 19839 16448 19848
rect 16396 19805 16405 19839
rect 16405 19805 16439 19839
rect 16439 19805 16448 19839
rect 16396 19796 16448 19805
rect 17132 19864 17184 19916
rect 17776 19796 17828 19848
rect 22376 19864 22428 19916
rect 21088 19839 21140 19848
rect 21088 19805 21097 19839
rect 21097 19805 21131 19839
rect 21131 19805 21140 19839
rect 21088 19796 21140 19805
rect 9956 19728 10008 19780
rect 10600 19728 10652 19780
rect 7656 19660 7708 19712
rect 12808 19660 12860 19712
rect 18420 19728 18472 19780
rect 20260 19728 20312 19780
rect 21824 19796 21876 19848
rect 21916 19839 21968 19848
rect 21916 19805 21925 19839
rect 21925 19805 21959 19839
rect 21959 19805 21968 19839
rect 21916 19796 21968 19805
rect 21180 19660 21232 19712
rect 22284 19771 22336 19780
rect 22284 19737 22293 19771
rect 22293 19737 22327 19771
rect 22327 19737 22336 19771
rect 33140 19839 33192 19848
rect 33140 19805 33149 19839
rect 33149 19805 33183 19839
rect 33183 19805 33192 19839
rect 33140 19796 33192 19805
rect 22284 19728 22336 19737
rect 34612 19728 34664 19780
rect 22652 19660 22704 19712
rect 9390 19558 9442 19610
rect 9454 19558 9506 19610
rect 9518 19558 9570 19610
rect 9582 19558 9634 19610
rect 9646 19558 9698 19610
rect 17831 19558 17883 19610
rect 17895 19558 17947 19610
rect 17959 19558 18011 19610
rect 18023 19558 18075 19610
rect 18087 19558 18139 19610
rect 26272 19558 26324 19610
rect 26336 19558 26388 19610
rect 26400 19558 26452 19610
rect 26464 19558 26516 19610
rect 26528 19558 26580 19610
rect 34713 19558 34765 19610
rect 34777 19558 34829 19610
rect 34841 19558 34893 19610
rect 34905 19558 34957 19610
rect 34969 19558 35021 19610
rect 10600 19499 10652 19508
rect 10600 19465 10609 19499
rect 10609 19465 10643 19499
rect 10643 19465 10652 19499
rect 10600 19456 10652 19465
rect 10692 19456 10744 19508
rect 12440 19456 12492 19508
rect 14372 19456 14424 19508
rect 14464 19456 14516 19508
rect 16396 19456 16448 19508
rect 18420 19499 18472 19508
rect 18420 19465 18429 19499
rect 18429 19465 18463 19499
rect 18463 19465 18472 19499
rect 18420 19456 18472 19465
rect 18880 19456 18932 19508
rect 20720 19456 20772 19508
rect 21548 19456 21600 19508
rect 22284 19456 22336 19508
rect 11060 19320 11112 19372
rect 11888 19320 11940 19372
rect 12348 19320 12400 19372
rect 14556 19431 14608 19440
rect 14556 19397 14565 19431
rect 14565 19397 14599 19431
rect 14599 19397 14608 19431
rect 14556 19388 14608 19397
rect 14924 19320 14976 19372
rect 18696 19320 18748 19372
rect 18788 19363 18840 19372
rect 18788 19329 18797 19363
rect 18797 19329 18831 19363
rect 18831 19329 18840 19363
rect 18788 19320 18840 19329
rect 19616 19363 19668 19372
rect 19616 19329 19625 19363
rect 19625 19329 19659 19363
rect 19659 19329 19668 19363
rect 19616 19320 19668 19329
rect 14096 19252 14148 19304
rect 20904 19252 20956 19304
rect 5170 19014 5222 19066
rect 5234 19014 5286 19066
rect 5298 19014 5350 19066
rect 5362 19014 5414 19066
rect 5426 19014 5478 19066
rect 13611 19014 13663 19066
rect 13675 19014 13727 19066
rect 13739 19014 13791 19066
rect 13803 19014 13855 19066
rect 13867 19014 13919 19066
rect 22052 19014 22104 19066
rect 22116 19014 22168 19066
rect 22180 19014 22232 19066
rect 22244 19014 22296 19066
rect 22308 19014 22360 19066
rect 30493 19014 30545 19066
rect 30557 19014 30609 19066
rect 30621 19014 30673 19066
rect 30685 19014 30737 19066
rect 30749 19014 30801 19066
rect 9390 18470 9442 18522
rect 9454 18470 9506 18522
rect 9518 18470 9570 18522
rect 9582 18470 9634 18522
rect 9646 18470 9698 18522
rect 17831 18470 17883 18522
rect 17895 18470 17947 18522
rect 17959 18470 18011 18522
rect 18023 18470 18075 18522
rect 18087 18470 18139 18522
rect 26272 18470 26324 18522
rect 26336 18470 26388 18522
rect 26400 18470 26452 18522
rect 26464 18470 26516 18522
rect 26528 18470 26580 18522
rect 34713 18470 34765 18522
rect 34777 18470 34829 18522
rect 34841 18470 34893 18522
rect 34905 18470 34957 18522
rect 34969 18470 35021 18522
rect 5170 17926 5222 17978
rect 5234 17926 5286 17978
rect 5298 17926 5350 17978
rect 5362 17926 5414 17978
rect 5426 17926 5478 17978
rect 13611 17926 13663 17978
rect 13675 17926 13727 17978
rect 13739 17926 13791 17978
rect 13803 17926 13855 17978
rect 13867 17926 13919 17978
rect 22052 17926 22104 17978
rect 22116 17926 22168 17978
rect 22180 17926 22232 17978
rect 22244 17926 22296 17978
rect 22308 17926 22360 17978
rect 30493 17926 30545 17978
rect 30557 17926 30609 17978
rect 30621 17926 30673 17978
rect 30685 17926 30737 17978
rect 30749 17926 30801 17978
rect 9390 17382 9442 17434
rect 9454 17382 9506 17434
rect 9518 17382 9570 17434
rect 9582 17382 9634 17434
rect 9646 17382 9698 17434
rect 17831 17382 17883 17434
rect 17895 17382 17947 17434
rect 17959 17382 18011 17434
rect 18023 17382 18075 17434
rect 18087 17382 18139 17434
rect 26272 17382 26324 17434
rect 26336 17382 26388 17434
rect 26400 17382 26452 17434
rect 26464 17382 26516 17434
rect 26528 17382 26580 17434
rect 34713 17382 34765 17434
rect 34777 17382 34829 17434
rect 34841 17382 34893 17434
rect 34905 17382 34957 17434
rect 34969 17382 35021 17434
rect 5170 16838 5222 16890
rect 5234 16838 5286 16890
rect 5298 16838 5350 16890
rect 5362 16838 5414 16890
rect 5426 16838 5478 16890
rect 13611 16838 13663 16890
rect 13675 16838 13727 16890
rect 13739 16838 13791 16890
rect 13803 16838 13855 16890
rect 13867 16838 13919 16890
rect 22052 16838 22104 16890
rect 22116 16838 22168 16890
rect 22180 16838 22232 16890
rect 22244 16838 22296 16890
rect 22308 16838 22360 16890
rect 30493 16838 30545 16890
rect 30557 16838 30609 16890
rect 30621 16838 30673 16890
rect 30685 16838 30737 16890
rect 30749 16838 30801 16890
rect 9390 16294 9442 16346
rect 9454 16294 9506 16346
rect 9518 16294 9570 16346
rect 9582 16294 9634 16346
rect 9646 16294 9698 16346
rect 17831 16294 17883 16346
rect 17895 16294 17947 16346
rect 17959 16294 18011 16346
rect 18023 16294 18075 16346
rect 18087 16294 18139 16346
rect 26272 16294 26324 16346
rect 26336 16294 26388 16346
rect 26400 16294 26452 16346
rect 26464 16294 26516 16346
rect 26528 16294 26580 16346
rect 34713 16294 34765 16346
rect 34777 16294 34829 16346
rect 34841 16294 34893 16346
rect 34905 16294 34957 16346
rect 34969 16294 35021 16346
rect 5170 15750 5222 15802
rect 5234 15750 5286 15802
rect 5298 15750 5350 15802
rect 5362 15750 5414 15802
rect 5426 15750 5478 15802
rect 13611 15750 13663 15802
rect 13675 15750 13727 15802
rect 13739 15750 13791 15802
rect 13803 15750 13855 15802
rect 13867 15750 13919 15802
rect 22052 15750 22104 15802
rect 22116 15750 22168 15802
rect 22180 15750 22232 15802
rect 22244 15750 22296 15802
rect 22308 15750 22360 15802
rect 30493 15750 30545 15802
rect 30557 15750 30609 15802
rect 30621 15750 30673 15802
rect 30685 15750 30737 15802
rect 30749 15750 30801 15802
rect 9390 15206 9442 15258
rect 9454 15206 9506 15258
rect 9518 15206 9570 15258
rect 9582 15206 9634 15258
rect 9646 15206 9698 15258
rect 17831 15206 17883 15258
rect 17895 15206 17947 15258
rect 17959 15206 18011 15258
rect 18023 15206 18075 15258
rect 18087 15206 18139 15258
rect 26272 15206 26324 15258
rect 26336 15206 26388 15258
rect 26400 15206 26452 15258
rect 26464 15206 26516 15258
rect 26528 15206 26580 15258
rect 34713 15206 34765 15258
rect 34777 15206 34829 15258
rect 34841 15206 34893 15258
rect 34905 15206 34957 15258
rect 34969 15206 35021 15258
rect 5170 14662 5222 14714
rect 5234 14662 5286 14714
rect 5298 14662 5350 14714
rect 5362 14662 5414 14714
rect 5426 14662 5478 14714
rect 13611 14662 13663 14714
rect 13675 14662 13727 14714
rect 13739 14662 13791 14714
rect 13803 14662 13855 14714
rect 13867 14662 13919 14714
rect 22052 14662 22104 14714
rect 22116 14662 22168 14714
rect 22180 14662 22232 14714
rect 22244 14662 22296 14714
rect 22308 14662 22360 14714
rect 30493 14662 30545 14714
rect 30557 14662 30609 14714
rect 30621 14662 30673 14714
rect 30685 14662 30737 14714
rect 30749 14662 30801 14714
rect 1584 14603 1636 14612
rect 1584 14569 1593 14603
rect 1593 14569 1627 14603
rect 1627 14569 1636 14603
rect 1584 14560 1636 14569
rect 940 14356 992 14408
rect 9390 14118 9442 14170
rect 9454 14118 9506 14170
rect 9518 14118 9570 14170
rect 9582 14118 9634 14170
rect 9646 14118 9698 14170
rect 17831 14118 17883 14170
rect 17895 14118 17947 14170
rect 17959 14118 18011 14170
rect 18023 14118 18075 14170
rect 18087 14118 18139 14170
rect 26272 14118 26324 14170
rect 26336 14118 26388 14170
rect 26400 14118 26452 14170
rect 26464 14118 26516 14170
rect 26528 14118 26580 14170
rect 34713 14118 34765 14170
rect 34777 14118 34829 14170
rect 34841 14118 34893 14170
rect 34905 14118 34957 14170
rect 34969 14118 35021 14170
rect 5170 13574 5222 13626
rect 5234 13574 5286 13626
rect 5298 13574 5350 13626
rect 5362 13574 5414 13626
rect 5426 13574 5478 13626
rect 13611 13574 13663 13626
rect 13675 13574 13727 13626
rect 13739 13574 13791 13626
rect 13803 13574 13855 13626
rect 13867 13574 13919 13626
rect 22052 13574 22104 13626
rect 22116 13574 22168 13626
rect 22180 13574 22232 13626
rect 22244 13574 22296 13626
rect 22308 13574 22360 13626
rect 30493 13574 30545 13626
rect 30557 13574 30609 13626
rect 30621 13574 30673 13626
rect 30685 13574 30737 13626
rect 30749 13574 30801 13626
rect 24032 13132 24084 13184
rect 35164 13132 35216 13184
rect 9390 13030 9442 13082
rect 9454 13030 9506 13082
rect 9518 13030 9570 13082
rect 9582 13030 9634 13082
rect 9646 13030 9698 13082
rect 17831 13030 17883 13082
rect 17895 13030 17947 13082
rect 17959 13030 18011 13082
rect 18023 13030 18075 13082
rect 18087 13030 18139 13082
rect 26272 13030 26324 13082
rect 26336 13030 26388 13082
rect 26400 13030 26452 13082
rect 26464 13030 26516 13082
rect 26528 13030 26580 13082
rect 34713 13030 34765 13082
rect 34777 13030 34829 13082
rect 34841 13030 34893 13082
rect 34905 13030 34957 13082
rect 34969 13030 35021 13082
rect 5170 12486 5222 12538
rect 5234 12486 5286 12538
rect 5298 12486 5350 12538
rect 5362 12486 5414 12538
rect 5426 12486 5478 12538
rect 13611 12486 13663 12538
rect 13675 12486 13727 12538
rect 13739 12486 13791 12538
rect 13803 12486 13855 12538
rect 13867 12486 13919 12538
rect 22052 12486 22104 12538
rect 22116 12486 22168 12538
rect 22180 12486 22232 12538
rect 22244 12486 22296 12538
rect 22308 12486 22360 12538
rect 30493 12486 30545 12538
rect 30557 12486 30609 12538
rect 30621 12486 30673 12538
rect 30685 12486 30737 12538
rect 30749 12486 30801 12538
rect 9390 11942 9442 11994
rect 9454 11942 9506 11994
rect 9518 11942 9570 11994
rect 9582 11942 9634 11994
rect 9646 11942 9698 11994
rect 17831 11942 17883 11994
rect 17895 11942 17947 11994
rect 17959 11942 18011 11994
rect 18023 11942 18075 11994
rect 18087 11942 18139 11994
rect 26272 11942 26324 11994
rect 26336 11942 26388 11994
rect 26400 11942 26452 11994
rect 26464 11942 26516 11994
rect 26528 11942 26580 11994
rect 34713 11942 34765 11994
rect 34777 11942 34829 11994
rect 34841 11942 34893 11994
rect 34905 11942 34957 11994
rect 34969 11942 35021 11994
rect 5170 11398 5222 11450
rect 5234 11398 5286 11450
rect 5298 11398 5350 11450
rect 5362 11398 5414 11450
rect 5426 11398 5478 11450
rect 13611 11398 13663 11450
rect 13675 11398 13727 11450
rect 13739 11398 13791 11450
rect 13803 11398 13855 11450
rect 13867 11398 13919 11450
rect 22052 11398 22104 11450
rect 22116 11398 22168 11450
rect 22180 11398 22232 11450
rect 22244 11398 22296 11450
rect 22308 11398 22360 11450
rect 30493 11398 30545 11450
rect 30557 11398 30609 11450
rect 30621 11398 30673 11450
rect 30685 11398 30737 11450
rect 30749 11398 30801 11450
rect 9390 10854 9442 10906
rect 9454 10854 9506 10906
rect 9518 10854 9570 10906
rect 9582 10854 9634 10906
rect 9646 10854 9698 10906
rect 17831 10854 17883 10906
rect 17895 10854 17947 10906
rect 17959 10854 18011 10906
rect 18023 10854 18075 10906
rect 18087 10854 18139 10906
rect 26272 10854 26324 10906
rect 26336 10854 26388 10906
rect 26400 10854 26452 10906
rect 26464 10854 26516 10906
rect 26528 10854 26580 10906
rect 34713 10854 34765 10906
rect 34777 10854 34829 10906
rect 34841 10854 34893 10906
rect 34905 10854 34957 10906
rect 34969 10854 35021 10906
rect 5170 10310 5222 10362
rect 5234 10310 5286 10362
rect 5298 10310 5350 10362
rect 5362 10310 5414 10362
rect 5426 10310 5478 10362
rect 13611 10310 13663 10362
rect 13675 10310 13727 10362
rect 13739 10310 13791 10362
rect 13803 10310 13855 10362
rect 13867 10310 13919 10362
rect 22052 10310 22104 10362
rect 22116 10310 22168 10362
rect 22180 10310 22232 10362
rect 22244 10310 22296 10362
rect 22308 10310 22360 10362
rect 30493 10310 30545 10362
rect 30557 10310 30609 10362
rect 30621 10310 30673 10362
rect 30685 10310 30737 10362
rect 30749 10310 30801 10362
rect 9390 9766 9442 9818
rect 9454 9766 9506 9818
rect 9518 9766 9570 9818
rect 9582 9766 9634 9818
rect 9646 9766 9698 9818
rect 17831 9766 17883 9818
rect 17895 9766 17947 9818
rect 17959 9766 18011 9818
rect 18023 9766 18075 9818
rect 18087 9766 18139 9818
rect 26272 9766 26324 9818
rect 26336 9766 26388 9818
rect 26400 9766 26452 9818
rect 26464 9766 26516 9818
rect 26528 9766 26580 9818
rect 34713 9766 34765 9818
rect 34777 9766 34829 9818
rect 34841 9766 34893 9818
rect 34905 9766 34957 9818
rect 34969 9766 35021 9818
rect 5170 9222 5222 9274
rect 5234 9222 5286 9274
rect 5298 9222 5350 9274
rect 5362 9222 5414 9274
rect 5426 9222 5478 9274
rect 13611 9222 13663 9274
rect 13675 9222 13727 9274
rect 13739 9222 13791 9274
rect 13803 9222 13855 9274
rect 13867 9222 13919 9274
rect 22052 9222 22104 9274
rect 22116 9222 22168 9274
rect 22180 9222 22232 9274
rect 22244 9222 22296 9274
rect 22308 9222 22360 9274
rect 30493 9222 30545 9274
rect 30557 9222 30609 9274
rect 30621 9222 30673 9274
rect 30685 9222 30737 9274
rect 30749 9222 30801 9274
rect 9390 8678 9442 8730
rect 9454 8678 9506 8730
rect 9518 8678 9570 8730
rect 9582 8678 9634 8730
rect 9646 8678 9698 8730
rect 17831 8678 17883 8730
rect 17895 8678 17947 8730
rect 17959 8678 18011 8730
rect 18023 8678 18075 8730
rect 18087 8678 18139 8730
rect 26272 8678 26324 8730
rect 26336 8678 26388 8730
rect 26400 8678 26452 8730
rect 26464 8678 26516 8730
rect 26528 8678 26580 8730
rect 34713 8678 34765 8730
rect 34777 8678 34829 8730
rect 34841 8678 34893 8730
rect 34905 8678 34957 8730
rect 34969 8678 35021 8730
rect 5170 8134 5222 8186
rect 5234 8134 5286 8186
rect 5298 8134 5350 8186
rect 5362 8134 5414 8186
rect 5426 8134 5478 8186
rect 13611 8134 13663 8186
rect 13675 8134 13727 8186
rect 13739 8134 13791 8186
rect 13803 8134 13855 8186
rect 13867 8134 13919 8186
rect 22052 8134 22104 8186
rect 22116 8134 22168 8186
rect 22180 8134 22232 8186
rect 22244 8134 22296 8186
rect 22308 8134 22360 8186
rect 30493 8134 30545 8186
rect 30557 8134 30609 8186
rect 30621 8134 30673 8186
rect 30685 8134 30737 8186
rect 30749 8134 30801 8186
rect 9390 7590 9442 7642
rect 9454 7590 9506 7642
rect 9518 7590 9570 7642
rect 9582 7590 9634 7642
rect 9646 7590 9698 7642
rect 17831 7590 17883 7642
rect 17895 7590 17947 7642
rect 17959 7590 18011 7642
rect 18023 7590 18075 7642
rect 18087 7590 18139 7642
rect 26272 7590 26324 7642
rect 26336 7590 26388 7642
rect 26400 7590 26452 7642
rect 26464 7590 26516 7642
rect 26528 7590 26580 7642
rect 34713 7590 34765 7642
rect 34777 7590 34829 7642
rect 34841 7590 34893 7642
rect 34905 7590 34957 7642
rect 34969 7590 35021 7642
rect 1400 7191 1452 7200
rect 1400 7157 1409 7191
rect 1409 7157 1443 7191
rect 1443 7157 1452 7191
rect 1400 7148 1452 7157
rect 5170 7046 5222 7098
rect 5234 7046 5286 7098
rect 5298 7046 5350 7098
rect 5362 7046 5414 7098
rect 5426 7046 5478 7098
rect 13611 7046 13663 7098
rect 13675 7046 13727 7098
rect 13739 7046 13791 7098
rect 13803 7046 13855 7098
rect 13867 7046 13919 7098
rect 22052 7046 22104 7098
rect 22116 7046 22168 7098
rect 22180 7046 22232 7098
rect 22244 7046 22296 7098
rect 22308 7046 22360 7098
rect 30493 7046 30545 7098
rect 30557 7046 30609 7098
rect 30621 7046 30673 7098
rect 30685 7046 30737 7098
rect 30749 7046 30801 7098
rect 9390 6502 9442 6554
rect 9454 6502 9506 6554
rect 9518 6502 9570 6554
rect 9582 6502 9634 6554
rect 9646 6502 9698 6554
rect 17831 6502 17883 6554
rect 17895 6502 17947 6554
rect 17959 6502 18011 6554
rect 18023 6502 18075 6554
rect 18087 6502 18139 6554
rect 26272 6502 26324 6554
rect 26336 6502 26388 6554
rect 26400 6502 26452 6554
rect 26464 6502 26516 6554
rect 26528 6502 26580 6554
rect 34713 6502 34765 6554
rect 34777 6502 34829 6554
rect 34841 6502 34893 6554
rect 34905 6502 34957 6554
rect 34969 6502 35021 6554
rect 5170 5958 5222 6010
rect 5234 5958 5286 6010
rect 5298 5958 5350 6010
rect 5362 5958 5414 6010
rect 5426 5958 5478 6010
rect 13611 5958 13663 6010
rect 13675 5958 13727 6010
rect 13739 5958 13791 6010
rect 13803 5958 13855 6010
rect 13867 5958 13919 6010
rect 22052 5958 22104 6010
rect 22116 5958 22168 6010
rect 22180 5958 22232 6010
rect 22244 5958 22296 6010
rect 22308 5958 22360 6010
rect 30493 5958 30545 6010
rect 30557 5958 30609 6010
rect 30621 5958 30673 6010
rect 30685 5958 30737 6010
rect 30749 5958 30801 6010
rect 34520 5627 34572 5636
rect 34520 5593 34529 5627
rect 34529 5593 34563 5627
rect 34563 5593 34572 5627
rect 34520 5584 34572 5593
rect 9390 5414 9442 5466
rect 9454 5414 9506 5466
rect 9518 5414 9570 5466
rect 9582 5414 9634 5466
rect 9646 5414 9698 5466
rect 17831 5414 17883 5466
rect 17895 5414 17947 5466
rect 17959 5414 18011 5466
rect 18023 5414 18075 5466
rect 18087 5414 18139 5466
rect 26272 5414 26324 5466
rect 26336 5414 26388 5466
rect 26400 5414 26452 5466
rect 26464 5414 26516 5466
rect 26528 5414 26580 5466
rect 34713 5414 34765 5466
rect 34777 5414 34829 5466
rect 34841 5414 34893 5466
rect 34905 5414 34957 5466
rect 34969 5414 35021 5466
rect 5170 4870 5222 4922
rect 5234 4870 5286 4922
rect 5298 4870 5350 4922
rect 5362 4870 5414 4922
rect 5426 4870 5478 4922
rect 13611 4870 13663 4922
rect 13675 4870 13727 4922
rect 13739 4870 13791 4922
rect 13803 4870 13855 4922
rect 13867 4870 13919 4922
rect 22052 4870 22104 4922
rect 22116 4870 22168 4922
rect 22180 4870 22232 4922
rect 22244 4870 22296 4922
rect 22308 4870 22360 4922
rect 30493 4870 30545 4922
rect 30557 4870 30609 4922
rect 30621 4870 30673 4922
rect 30685 4870 30737 4922
rect 30749 4870 30801 4922
rect 9390 4326 9442 4378
rect 9454 4326 9506 4378
rect 9518 4326 9570 4378
rect 9582 4326 9634 4378
rect 9646 4326 9698 4378
rect 17831 4326 17883 4378
rect 17895 4326 17947 4378
rect 17959 4326 18011 4378
rect 18023 4326 18075 4378
rect 18087 4326 18139 4378
rect 26272 4326 26324 4378
rect 26336 4326 26388 4378
rect 26400 4326 26452 4378
rect 26464 4326 26516 4378
rect 26528 4326 26580 4378
rect 34713 4326 34765 4378
rect 34777 4326 34829 4378
rect 34841 4326 34893 4378
rect 34905 4326 34957 4378
rect 34969 4326 35021 4378
rect 5170 3782 5222 3834
rect 5234 3782 5286 3834
rect 5298 3782 5350 3834
rect 5362 3782 5414 3834
rect 5426 3782 5478 3834
rect 13611 3782 13663 3834
rect 13675 3782 13727 3834
rect 13739 3782 13791 3834
rect 13803 3782 13855 3834
rect 13867 3782 13919 3834
rect 22052 3782 22104 3834
rect 22116 3782 22168 3834
rect 22180 3782 22232 3834
rect 22244 3782 22296 3834
rect 22308 3782 22360 3834
rect 30493 3782 30545 3834
rect 30557 3782 30609 3834
rect 30621 3782 30673 3834
rect 30685 3782 30737 3834
rect 30749 3782 30801 3834
rect 9390 3238 9442 3290
rect 9454 3238 9506 3290
rect 9518 3238 9570 3290
rect 9582 3238 9634 3290
rect 9646 3238 9698 3290
rect 17831 3238 17883 3290
rect 17895 3238 17947 3290
rect 17959 3238 18011 3290
rect 18023 3238 18075 3290
rect 18087 3238 18139 3290
rect 26272 3238 26324 3290
rect 26336 3238 26388 3290
rect 26400 3238 26452 3290
rect 26464 3238 26516 3290
rect 26528 3238 26580 3290
rect 34713 3238 34765 3290
rect 34777 3238 34829 3290
rect 34841 3238 34893 3290
rect 34905 3238 34957 3290
rect 34969 3238 35021 3290
rect 5170 2694 5222 2746
rect 5234 2694 5286 2746
rect 5298 2694 5350 2746
rect 5362 2694 5414 2746
rect 5426 2694 5478 2746
rect 13611 2694 13663 2746
rect 13675 2694 13727 2746
rect 13739 2694 13791 2746
rect 13803 2694 13855 2746
rect 13867 2694 13919 2746
rect 22052 2694 22104 2746
rect 22116 2694 22168 2746
rect 22180 2694 22232 2746
rect 22244 2694 22296 2746
rect 22308 2694 22360 2746
rect 30493 2694 30545 2746
rect 30557 2694 30609 2746
rect 30621 2694 30673 2746
rect 30685 2694 30737 2746
rect 30749 2694 30801 2746
rect 20720 2499 20772 2508
rect 20720 2465 20729 2499
rect 20729 2465 20763 2499
rect 20763 2465 20772 2499
rect 20720 2456 20772 2465
rect 13636 2431 13688 2440
rect 13636 2397 13645 2431
rect 13645 2397 13679 2431
rect 13679 2397 13688 2431
rect 13636 2388 13688 2397
rect 20260 2431 20312 2440
rect 20260 2397 20269 2431
rect 20269 2397 20303 2431
rect 20303 2397 20312 2431
rect 20260 2388 20312 2397
rect 20 2252 72 2304
rect 6552 2295 6604 2304
rect 6552 2261 6561 2295
rect 6561 2261 6595 2295
rect 6595 2261 6604 2295
rect 6552 2252 6604 2261
rect 27160 2295 27212 2304
rect 27160 2261 27169 2295
rect 27169 2261 27203 2295
rect 27203 2261 27212 2295
rect 27160 2252 27212 2261
rect 34244 2295 34296 2304
rect 34244 2261 34253 2295
rect 34253 2261 34287 2295
rect 34287 2261 34296 2295
rect 34244 2252 34296 2261
rect 9390 2150 9442 2202
rect 9454 2150 9506 2202
rect 9518 2150 9570 2202
rect 9582 2150 9634 2202
rect 9646 2150 9698 2202
rect 17831 2150 17883 2202
rect 17895 2150 17947 2202
rect 17959 2150 18011 2202
rect 18023 2150 18075 2202
rect 18087 2150 18139 2202
rect 26272 2150 26324 2202
rect 26336 2150 26388 2202
rect 26400 2150 26452 2202
rect 26464 2150 26516 2202
rect 26528 2150 26580 2202
rect 34713 2150 34765 2202
rect 34777 2150 34829 2202
rect 34841 2150 34893 2202
rect 34905 2150 34957 2202
rect 34969 2150 35021 2202
<< metal2 >>
rect 1278 41200 1390 42000
rect 8362 41200 8474 42000
rect 14802 41200 14914 42000
rect 21886 41200 21998 42000
rect 28970 41200 29082 42000
rect 35410 41200 35522 42000
rect 1320 38962 1348 41200
rect 5170 39740 5478 39749
rect 5170 39738 5176 39740
rect 5232 39738 5256 39740
rect 5312 39738 5336 39740
rect 5392 39738 5416 39740
rect 5472 39738 5478 39740
rect 5232 39686 5234 39738
rect 5414 39686 5416 39738
rect 5170 39684 5176 39686
rect 5232 39684 5256 39686
rect 5312 39684 5336 39686
rect 5392 39684 5416 39686
rect 5472 39684 5478 39686
rect 5170 39675 5478 39684
rect 8404 39438 8432 41200
rect 13611 39740 13919 39749
rect 13611 39738 13617 39740
rect 13673 39738 13697 39740
rect 13753 39738 13777 39740
rect 13833 39738 13857 39740
rect 13913 39738 13919 39740
rect 13673 39686 13675 39738
rect 13855 39686 13857 39738
rect 13611 39684 13617 39686
rect 13673 39684 13697 39686
rect 13753 39684 13777 39686
rect 13833 39684 13857 39686
rect 13913 39684 13919 39686
rect 13611 39675 13919 39684
rect 14844 39438 14872 41200
rect 18328 39636 18380 39642
rect 18328 39578 18380 39584
rect 16396 39500 16448 39506
rect 16396 39442 16448 39448
rect 3056 39432 3108 39438
rect 3056 39374 3108 39380
rect 8392 39432 8444 39438
rect 8392 39374 8444 39380
rect 14832 39432 14884 39438
rect 14832 39374 14884 39380
rect 3068 39098 3096 39374
rect 16120 39364 16172 39370
rect 16120 39306 16172 39312
rect 4896 39296 4948 39302
rect 4896 39238 4948 39244
rect 8484 39296 8536 39302
rect 8484 39238 8536 39244
rect 13912 39296 13964 39302
rect 13912 39238 13964 39244
rect 15292 39296 15344 39302
rect 15292 39238 15344 39244
rect 15384 39296 15436 39302
rect 15384 39238 15436 39244
rect 3056 39092 3108 39098
rect 3056 39034 3108 39040
rect 1308 38956 1360 38962
rect 1308 38898 1360 38904
rect 4908 38350 4936 39238
rect 5170 38652 5478 38661
rect 5170 38650 5176 38652
rect 5232 38650 5256 38652
rect 5312 38650 5336 38652
rect 5392 38650 5416 38652
rect 5472 38650 5478 38652
rect 5232 38598 5234 38650
rect 5414 38598 5416 38650
rect 5170 38596 5176 38598
rect 5232 38596 5256 38598
rect 5312 38596 5336 38598
rect 5392 38596 5416 38598
rect 5472 38596 5478 38598
rect 5170 38587 5478 38596
rect 8496 38350 8524 39238
rect 9390 39196 9698 39205
rect 9390 39194 9396 39196
rect 9452 39194 9476 39196
rect 9532 39194 9556 39196
rect 9612 39194 9636 39196
rect 9692 39194 9698 39196
rect 9452 39142 9454 39194
rect 9634 39142 9636 39194
rect 9390 39140 9396 39142
rect 9452 39140 9476 39142
rect 9532 39140 9556 39142
rect 9612 39140 9636 39142
rect 9692 39140 9698 39142
rect 9390 39131 9698 39140
rect 13924 39098 13952 39238
rect 13912 39092 13964 39098
rect 13912 39034 13964 39040
rect 14096 38888 14148 38894
rect 14096 38830 14148 38836
rect 13611 38652 13919 38661
rect 13611 38650 13617 38652
rect 13673 38650 13697 38652
rect 13753 38650 13777 38652
rect 13833 38650 13857 38652
rect 13913 38650 13919 38652
rect 13673 38598 13675 38650
rect 13855 38598 13857 38650
rect 13611 38596 13617 38598
rect 13673 38596 13697 38598
rect 13753 38596 13777 38598
rect 13833 38596 13857 38598
rect 13913 38596 13919 38598
rect 13611 38587 13919 38596
rect 14108 38350 14136 38830
rect 15304 38554 15332 39238
rect 15396 38962 15424 39238
rect 15384 38956 15436 38962
rect 15384 38898 15436 38904
rect 15292 38548 15344 38554
rect 15292 38490 15344 38496
rect 4896 38344 4948 38350
rect 4896 38286 4948 38292
rect 7472 38344 7524 38350
rect 7472 38286 7524 38292
rect 8392 38344 8444 38350
rect 8392 38286 8444 38292
rect 8484 38344 8536 38350
rect 8484 38286 8536 38292
rect 14096 38344 14148 38350
rect 14096 38286 14148 38292
rect 6920 38208 6972 38214
rect 6920 38150 6972 38156
rect 6000 37800 6052 37806
rect 6000 37742 6052 37748
rect 5170 37564 5478 37573
rect 5170 37562 5176 37564
rect 5232 37562 5256 37564
rect 5312 37562 5336 37564
rect 5392 37562 5416 37564
rect 5472 37562 5478 37564
rect 5232 37510 5234 37562
rect 5414 37510 5416 37562
rect 5170 37508 5176 37510
rect 5232 37508 5256 37510
rect 5312 37508 5336 37510
rect 5392 37508 5416 37510
rect 5472 37508 5478 37510
rect 5170 37499 5478 37508
rect 5170 36476 5478 36485
rect 5170 36474 5176 36476
rect 5232 36474 5256 36476
rect 5312 36474 5336 36476
rect 5392 36474 5416 36476
rect 5472 36474 5478 36476
rect 5232 36422 5234 36474
rect 5414 36422 5416 36474
rect 5170 36420 5176 36422
rect 5232 36420 5256 36422
rect 5312 36420 5336 36422
rect 5392 36420 5416 36422
rect 5472 36420 5478 36422
rect 5170 36411 5478 36420
rect 940 36168 992 36174
rect 938 36136 940 36145
rect 992 36136 994 36145
rect 938 36071 994 36080
rect 5170 35388 5478 35397
rect 5170 35386 5176 35388
rect 5232 35386 5256 35388
rect 5312 35386 5336 35388
rect 5392 35386 5416 35388
rect 5472 35386 5478 35388
rect 5232 35334 5234 35386
rect 5414 35334 5416 35386
rect 5170 35332 5176 35334
rect 5232 35332 5256 35334
rect 5312 35332 5336 35334
rect 5392 35332 5416 35334
rect 5472 35332 5478 35334
rect 5170 35323 5478 35332
rect 5170 34300 5478 34309
rect 5170 34298 5176 34300
rect 5232 34298 5256 34300
rect 5312 34298 5336 34300
rect 5392 34298 5416 34300
rect 5472 34298 5478 34300
rect 5232 34246 5234 34298
rect 5414 34246 5416 34298
rect 5170 34244 5176 34246
rect 5232 34244 5256 34246
rect 5312 34244 5336 34246
rect 5392 34244 5416 34246
rect 5472 34244 5478 34246
rect 5170 34235 5478 34244
rect 5170 33212 5478 33221
rect 5170 33210 5176 33212
rect 5232 33210 5256 33212
rect 5312 33210 5336 33212
rect 5392 33210 5416 33212
rect 5472 33210 5478 33212
rect 5232 33158 5234 33210
rect 5414 33158 5416 33210
rect 5170 33156 5176 33158
rect 5232 33156 5256 33158
rect 5312 33156 5336 33158
rect 5392 33156 5416 33158
rect 5472 33156 5478 33158
rect 5170 33147 5478 33156
rect 5170 32124 5478 32133
rect 5170 32122 5176 32124
rect 5232 32122 5256 32124
rect 5312 32122 5336 32124
rect 5392 32122 5416 32124
rect 5472 32122 5478 32124
rect 5232 32070 5234 32122
rect 5414 32070 5416 32122
rect 5170 32068 5176 32070
rect 5232 32068 5256 32070
rect 5312 32068 5336 32070
rect 5392 32068 5416 32070
rect 5472 32068 5478 32070
rect 5170 32059 5478 32068
rect 5170 31036 5478 31045
rect 5170 31034 5176 31036
rect 5232 31034 5256 31036
rect 5312 31034 5336 31036
rect 5392 31034 5416 31036
rect 5472 31034 5478 31036
rect 5232 30982 5234 31034
rect 5414 30982 5416 31034
rect 5170 30980 5176 30982
rect 5232 30980 5256 30982
rect 5312 30980 5336 30982
rect 5392 30980 5416 30982
rect 5472 30980 5478 30982
rect 5170 30971 5478 30980
rect 5170 29948 5478 29957
rect 5170 29946 5176 29948
rect 5232 29946 5256 29948
rect 5312 29946 5336 29948
rect 5392 29946 5416 29948
rect 5472 29946 5478 29948
rect 5232 29894 5234 29946
rect 5414 29894 5416 29946
rect 5170 29892 5176 29894
rect 5232 29892 5256 29894
rect 5312 29892 5336 29894
rect 5392 29892 5416 29894
rect 5472 29892 5478 29894
rect 5170 29883 5478 29892
rect 6012 29714 6040 37742
rect 6932 36174 6960 38150
rect 7288 37664 7340 37670
rect 7288 37606 7340 37612
rect 7300 37330 7328 37606
rect 7288 37324 7340 37330
rect 7288 37266 7340 37272
rect 7484 36786 7512 38286
rect 8404 37806 8432 38286
rect 8668 38208 8720 38214
rect 8668 38150 8720 38156
rect 8680 38010 8708 38150
rect 9390 38108 9698 38117
rect 9390 38106 9396 38108
rect 9452 38106 9476 38108
rect 9532 38106 9556 38108
rect 9612 38106 9636 38108
rect 9692 38106 9698 38108
rect 9452 38054 9454 38106
rect 9634 38054 9636 38106
rect 9390 38052 9396 38054
rect 9452 38052 9476 38054
rect 9532 38052 9556 38054
rect 9612 38052 9636 38054
rect 9692 38052 9698 38054
rect 9390 38043 9698 38052
rect 8668 38004 8720 38010
rect 8668 37946 8720 37952
rect 10508 37868 10560 37874
rect 10508 37810 10560 37816
rect 10692 37868 10744 37874
rect 10692 37810 10744 37816
rect 10784 37868 10836 37874
rect 10784 37810 10836 37816
rect 11152 37868 11204 37874
rect 11152 37810 11204 37816
rect 11704 37868 11756 37874
rect 11704 37810 11756 37816
rect 14004 37868 14056 37874
rect 14004 37810 14056 37816
rect 8392 37800 8444 37806
rect 8392 37742 8444 37748
rect 9036 37664 9088 37670
rect 9036 37606 9088 37612
rect 10140 37664 10192 37670
rect 10140 37606 10192 37612
rect 8852 37256 8904 37262
rect 8852 37198 8904 37204
rect 8024 37188 8076 37194
rect 8024 37130 8076 37136
rect 8036 36922 8064 37130
rect 8024 36916 8076 36922
rect 8024 36858 8076 36864
rect 8864 36786 8892 37198
rect 9048 36854 9076 37606
rect 10152 37194 10180 37606
rect 10140 37188 10192 37194
rect 10140 37130 10192 37136
rect 9128 37120 9180 37126
rect 9128 37062 9180 37068
rect 9036 36848 9088 36854
rect 9036 36790 9088 36796
rect 7472 36780 7524 36786
rect 7472 36722 7524 36728
rect 8852 36780 8904 36786
rect 8852 36722 8904 36728
rect 8576 36712 8628 36718
rect 8576 36654 8628 36660
rect 7656 36576 7708 36582
rect 7656 36518 7708 36524
rect 6920 36168 6972 36174
rect 6920 36110 6972 36116
rect 7380 33448 7432 33454
rect 7380 33390 7432 33396
rect 7392 31890 7420 33390
rect 7380 31884 7432 31890
rect 7380 31826 7432 31832
rect 6920 30660 6972 30666
rect 6920 30602 6972 30608
rect 6552 30252 6604 30258
rect 6552 30194 6604 30200
rect 6564 29850 6592 30194
rect 6932 30190 6960 30602
rect 6920 30184 6972 30190
rect 6920 30126 6972 30132
rect 6552 29844 6604 29850
rect 6552 29786 6604 29792
rect 6000 29708 6052 29714
rect 6000 29650 6052 29656
rect 1400 29164 1452 29170
rect 1400 29106 1452 29112
rect 1584 29164 1636 29170
rect 1584 29106 1636 29112
rect 1412 28937 1440 29106
rect 1398 28928 1454 28937
rect 1398 28863 1454 28872
rect 940 21956 992 21962
rect 940 21898 992 21904
rect 952 21865 980 21898
rect 938 21856 994 21865
rect 938 21791 994 21800
rect 1596 14618 1624 29106
rect 6012 29034 6040 29650
rect 6092 29640 6144 29646
rect 6092 29582 6144 29588
rect 7380 29640 7432 29646
rect 7380 29582 7432 29588
rect 6104 29306 6132 29582
rect 6092 29300 6144 29306
rect 6092 29242 6144 29248
rect 7392 29170 7420 29582
rect 6644 29164 6696 29170
rect 6644 29106 6696 29112
rect 7380 29164 7432 29170
rect 7380 29106 7432 29112
rect 6000 29028 6052 29034
rect 6000 28970 6052 28976
rect 6184 28960 6236 28966
rect 6184 28902 6236 28908
rect 5170 28860 5478 28869
rect 5170 28858 5176 28860
rect 5232 28858 5256 28860
rect 5312 28858 5336 28860
rect 5392 28858 5416 28860
rect 5472 28858 5478 28860
rect 5232 28806 5234 28858
rect 5414 28806 5416 28858
rect 5170 28804 5176 28806
rect 5232 28804 5256 28806
rect 5312 28804 5336 28806
rect 5392 28804 5416 28806
rect 5472 28804 5478 28806
rect 5170 28795 5478 28804
rect 6196 28558 6224 28902
rect 6656 28762 6684 29106
rect 6644 28756 6696 28762
rect 6644 28698 6696 28704
rect 6184 28552 6236 28558
rect 6184 28494 6236 28500
rect 7196 28416 7248 28422
rect 7196 28358 7248 28364
rect 7208 28218 7236 28358
rect 7196 28212 7248 28218
rect 7196 28154 7248 28160
rect 7392 28014 7420 29106
rect 7472 28416 7524 28422
rect 7472 28358 7524 28364
rect 7484 28082 7512 28358
rect 7472 28076 7524 28082
rect 7472 28018 7524 28024
rect 7380 28008 7432 28014
rect 7380 27950 7432 27956
rect 7196 27872 7248 27878
rect 7196 27814 7248 27820
rect 5170 27772 5478 27781
rect 5170 27770 5176 27772
rect 5232 27770 5256 27772
rect 5312 27770 5336 27772
rect 5392 27770 5416 27772
rect 5472 27770 5478 27772
rect 5232 27718 5234 27770
rect 5414 27718 5416 27770
rect 5170 27716 5176 27718
rect 5232 27716 5256 27718
rect 5312 27716 5336 27718
rect 5392 27716 5416 27718
rect 5472 27716 5478 27718
rect 5170 27707 5478 27716
rect 7208 27470 7236 27814
rect 7392 27470 7420 27950
rect 7196 27464 7248 27470
rect 7196 27406 7248 27412
rect 7380 27464 7432 27470
rect 7380 27406 7432 27412
rect 5170 26684 5478 26693
rect 5170 26682 5176 26684
rect 5232 26682 5256 26684
rect 5312 26682 5336 26684
rect 5392 26682 5416 26684
rect 5472 26682 5478 26684
rect 5232 26630 5234 26682
rect 5414 26630 5416 26682
rect 5170 26628 5176 26630
rect 5232 26628 5256 26630
rect 5312 26628 5336 26630
rect 5392 26628 5416 26630
rect 5472 26628 5478 26630
rect 5170 26619 5478 26628
rect 5170 25596 5478 25605
rect 5170 25594 5176 25596
rect 5232 25594 5256 25596
rect 5312 25594 5336 25596
rect 5392 25594 5416 25596
rect 5472 25594 5478 25596
rect 5232 25542 5234 25594
rect 5414 25542 5416 25594
rect 5170 25540 5176 25542
rect 5232 25540 5256 25542
rect 5312 25540 5336 25542
rect 5392 25540 5416 25542
rect 5472 25540 5478 25542
rect 5170 25531 5478 25540
rect 5170 24508 5478 24517
rect 5170 24506 5176 24508
rect 5232 24506 5256 24508
rect 5312 24506 5336 24508
rect 5392 24506 5416 24508
rect 5472 24506 5478 24508
rect 5232 24454 5234 24506
rect 5414 24454 5416 24506
rect 5170 24452 5176 24454
rect 5232 24452 5256 24454
rect 5312 24452 5336 24454
rect 5392 24452 5416 24454
rect 5472 24452 5478 24454
rect 5170 24443 5478 24452
rect 5170 23420 5478 23429
rect 5170 23418 5176 23420
rect 5232 23418 5256 23420
rect 5312 23418 5336 23420
rect 5392 23418 5416 23420
rect 5472 23418 5478 23420
rect 5232 23366 5234 23418
rect 5414 23366 5416 23418
rect 5170 23364 5176 23366
rect 5232 23364 5256 23366
rect 5312 23364 5336 23366
rect 5392 23364 5416 23366
rect 5472 23364 5478 23366
rect 5170 23355 5478 23364
rect 5170 22332 5478 22341
rect 5170 22330 5176 22332
rect 5232 22330 5256 22332
rect 5312 22330 5336 22332
rect 5392 22330 5416 22332
rect 5472 22330 5478 22332
rect 5232 22278 5234 22330
rect 5414 22278 5416 22330
rect 5170 22276 5176 22278
rect 5232 22276 5256 22278
rect 5312 22276 5336 22278
rect 5392 22276 5416 22278
rect 5472 22276 5478 22278
rect 5170 22267 5478 22276
rect 5170 21244 5478 21253
rect 5170 21242 5176 21244
rect 5232 21242 5256 21244
rect 5312 21242 5336 21244
rect 5392 21242 5416 21244
rect 5472 21242 5478 21244
rect 5232 21190 5234 21242
rect 5414 21190 5416 21242
rect 5170 21188 5176 21190
rect 5232 21188 5256 21190
rect 5312 21188 5336 21190
rect 5392 21188 5416 21190
rect 5472 21188 5478 21190
rect 5170 21179 5478 21188
rect 5170 20156 5478 20165
rect 5170 20154 5176 20156
rect 5232 20154 5256 20156
rect 5312 20154 5336 20156
rect 5392 20154 5416 20156
rect 5472 20154 5478 20156
rect 5232 20102 5234 20154
rect 5414 20102 5416 20154
rect 5170 20100 5176 20102
rect 5232 20100 5256 20102
rect 5312 20100 5336 20102
rect 5392 20100 5416 20102
rect 5472 20100 5478 20102
rect 5170 20091 5478 20100
rect 7668 19718 7696 36518
rect 8588 36378 8616 36654
rect 8576 36372 8628 36378
rect 8576 36314 8628 36320
rect 8864 35698 8892 36722
rect 9140 36378 9168 37062
rect 9390 37020 9698 37029
rect 9390 37018 9396 37020
rect 9452 37018 9476 37020
rect 9532 37018 9556 37020
rect 9612 37018 9636 37020
rect 9692 37018 9698 37020
rect 9452 36966 9454 37018
rect 9634 36966 9636 37018
rect 9390 36964 9396 36966
rect 9452 36964 9476 36966
rect 9532 36964 9556 36966
rect 9612 36964 9636 36966
rect 9692 36964 9698 36966
rect 9390 36955 9698 36964
rect 10048 36780 10100 36786
rect 10048 36722 10100 36728
rect 9128 36372 9180 36378
rect 9128 36314 9180 36320
rect 9772 36032 9824 36038
rect 9772 35974 9824 35980
rect 9956 36032 10008 36038
rect 9956 35974 10008 35980
rect 9390 35932 9698 35941
rect 9390 35930 9396 35932
rect 9452 35930 9476 35932
rect 9532 35930 9556 35932
rect 9612 35930 9636 35932
rect 9692 35930 9698 35932
rect 9452 35878 9454 35930
rect 9634 35878 9636 35930
rect 9390 35876 9396 35878
rect 9452 35876 9476 35878
rect 9532 35876 9556 35878
rect 9612 35876 9636 35878
rect 9692 35876 9698 35878
rect 9390 35867 9698 35876
rect 9784 35834 9812 35974
rect 9772 35828 9824 35834
rect 9772 35770 9824 35776
rect 8760 35692 8812 35698
rect 8760 35634 8812 35640
rect 8852 35692 8904 35698
rect 8852 35634 8904 35640
rect 8772 35290 8800 35634
rect 9312 35624 9364 35630
rect 9312 35566 9364 35572
rect 8760 35284 8812 35290
rect 8760 35226 8812 35232
rect 9324 35154 9352 35566
rect 9312 35148 9364 35154
rect 9312 35090 9364 35096
rect 9968 35086 9996 35974
rect 9956 35080 10008 35086
rect 9956 35022 10008 35028
rect 10060 35018 10088 36722
rect 10232 36576 10284 36582
rect 10232 36518 10284 36524
rect 10244 36378 10272 36518
rect 10232 36372 10284 36378
rect 10232 36314 10284 36320
rect 10048 35012 10100 35018
rect 10048 34954 10100 34960
rect 9390 34844 9698 34853
rect 9390 34842 9396 34844
rect 9452 34842 9476 34844
rect 9532 34842 9556 34844
rect 9612 34842 9636 34844
rect 9692 34842 9698 34844
rect 9452 34790 9454 34842
rect 9634 34790 9636 34842
rect 9390 34788 9396 34790
rect 9452 34788 9476 34790
rect 9532 34788 9556 34790
rect 9612 34788 9636 34790
rect 9692 34788 9698 34790
rect 9390 34779 9698 34788
rect 10060 34746 10088 34954
rect 10048 34740 10100 34746
rect 10048 34682 10100 34688
rect 9220 34604 9272 34610
rect 9956 34604 10008 34610
rect 9220 34546 9272 34552
rect 9692 34564 9956 34592
rect 8576 34536 8628 34542
rect 8576 34478 8628 34484
rect 8392 34128 8444 34134
rect 8392 34070 8444 34076
rect 8300 33856 8352 33862
rect 8300 33798 8352 33804
rect 8312 33658 8340 33798
rect 8300 33652 8352 33658
rect 8300 33594 8352 33600
rect 7932 33040 7984 33046
rect 7932 32982 7984 32988
rect 7840 32768 7892 32774
rect 7840 32710 7892 32716
rect 7852 32434 7880 32710
rect 7944 32434 7972 32982
rect 8300 32836 8352 32842
rect 8300 32778 8352 32784
rect 7840 32428 7892 32434
rect 7840 32370 7892 32376
rect 7932 32428 7984 32434
rect 7932 32370 7984 32376
rect 8116 32428 8168 32434
rect 8116 32370 8168 32376
rect 8024 31748 8076 31754
rect 8024 31690 8076 31696
rect 8036 31482 8064 31690
rect 8024 31476 8076 31482
rect 8024 31418 8076 31424
rect 8128 30938 8156 32370
rect 8312 31328 8340 32778
rect 8404 32366 8432 34070
rect 8484 33992 8536 33998
rect 8484 33934 8536 33940
rect 8496 33114 8524 33934
rect 8484 33108 8536 33114
rect 8484 33050 8536 33056
rect 8588 32910 8616 34478
rect 8944 34400 8996 34406
rect 8944 34342 8996 34348
rect 8760 34060 8812 34066
rect 8760 34002 8812 34008
rect 8772 33318 8800 34002
rect 8956 33998 8984 34342
rect 9232 34202 9260 34546
rect 9692 34474 9720 34564
rect 9956 34546 10008 34552
rect 10048 34604 10100 34610
rect 10048 34546 10100 34552
rect 9680 34468 9732 34474
rect 9680 34410 9732 34416
rect 9220 34196 9272 34202
rect 9220 34138 9272 34144
rect 8944 33992 8996 33998
rect 8944 33934 8996 33940
rect 8852 33924 8904 33930
rect 8852 33866 8904 33872
rect 9772 33924 9824 33930
rect 9772 33866 9824 33872
rect 8760 33312 8812 33318
rect 8760 33254 8812 33260
rect 8772 33046 8800 33254
rect 8760 33040 8812 33046
rect 8760 32982 8812 32988
rect 8576 32904 8628 32910
rect 8576 32846 8628 32852
rect 8484 32496 8536 32502
rect 8484 32438 8536 32444
rect 8392 32360 8444 32366
rect 8392 32302 8444 32308
rect 8496 31482 8524 32438
rect 8864 32366 8892 33866
rect 9220 33856 9272 33862
rect 9220 33798 9272 33804
rect 9232 32910 9260 33798
rect 9390 33756 9698 33765
rect 9390 33754 9396 33756
rect 9452 33754 9476 33756
rect 9532 33754 9556 33756
rect 9612 33754 9636 33756
rect 9692 33754 9698 33756
rect 9452 33702 9454 33754
rect 9634 33702 9636 33754
rect 9390 33700 9396 33702
rect 9452 33700 9476 33702
rect 9532 33700 9556 33702
rect 9612 33700 9636 33702
rect 9692 33700 9698 33702
rect 9390 33691 9698 33700
rect 9312 33652 9364 33658
rect 9312 33594 9364 33600
rect 9036 32904 9088 32910
rect 9036 32846 9088 32852
rect 9220 32904 9272 32910
rect 9220 32846 9272 32852
rect 8852 32360 8904 32366
rect 8852 32302 8904 32308
rect 8864 32026 8892 32302
rect 8944 32224 8996 32230
rect 8944 32166 8996 32172
rect 8852 32020 8904 32026
rect 8852 31962 8904 31968
rect 8864 31634 8892 31962
rect 8772 31606 8892 31634
rect 8484 31476 8536 31482
rect 8484 31418 8536 31424
rect 8772 31346 8800 31606
rect 8956 31414 8984 32166
rect 9048 31822 9076 32846
rect 9128 32836 9180 32842
rect 9128 32778 9180 32784
rect 9140 32502 9168 32778
rect 9128 32496 9180 32502
rect 9128 32438 9180 32444
rect 9324 32434 9352 33594
rect 9784 32774 9812 33866
rect 10060 33658 10088 34546
rect 10520 34406 10548 37810
rect 10600 36712 10652 36718
rect 10600 36654 10652 36660
rect 10612 36378 10640 36654
rect 10600 36372 10652 36378
rect 10600 36314 10652 36320
rect 10704 36106 10732 37810
rect 10796 36242 10824 37810
rect 11060 37800 11112 37806
rect 11060 37742 11112 37748
rect 10876 37664 10928 37670
rect 10876 37606 10928 37612
rect 10888 36718 10916 37606
rect 11072 37466 11100 37742
rect 11060 37460 11112 37466
rect 11060 37402 11112 37408
rect 10876 36712 10928 36718
rect 10876 36654 10928 36660
rect 10784 36236 10836 36242
rect 10784 36178 10836 36184
rect 10692 36100 10744 36106
rect 10692 36042 10744 36048
rect 10796 35222 10824 36178
rect 10888 36174 10916 36654
rect 11164 36242 11192 37810
rect 11520 37664 11572 37670
rect 11520 37606 11572 37612
rect 11532 37194 11560 37606
rect 11520 37188 11572 37194
rect 11520 37130 11572 37136
rect 11244 36576 11296 36582
rect 11244 36518 11296 36524
rect 11152 36236 11204 36242
rect 11152 36178 11204 36184
rect 10876 36168 10928 36174
rect 10876 36110 10928 36116
rect 11164 35834 11192 36178
rect 11152 35828 11204 35834
rect 11152 35770 11204 35776
rect 10784 35216 10836 35222
rect 10784 35158 10836 35164
rect 11256 35086 11284 36518
rect 11716 36378 11744 37810
rect 11980 37800 12032 37806
rect 11980 37742 12032 37748
rect 11704 36372 11756 36378
rect 11704 36314 11756 36320
rect 11992 36174 12020 37742
rect 12992 37732 13044 37738
rect 12992 37674 13044 37680
rect 12624 37664 12676 37670
rect 12624 37606 12676 37612
rect 12900 37664 12952 37670
rect 12900 37606 12952 37612
rect 12440 37120 12492 37126
rect 12440 37062 12492 37068
rect 12452 36922 12480 37062
rect 12440 36916 12492 36922
rect 12440 36858 12492 36864
rect 12532 36712 12584 36718
rect 12532 36654 12584 36660
rect 12440 36576 12492 36582
rect 12440 36518 12492 36524
rect 11980 36168 12032 36174
rect 11980 36110 12032 36116
rect 11796 35828 11848 35834
rect 11796 35770 11848 35776
rect 11612 35556 11664 35562
rect 11612 35498 11664 35504
rect 11624 35086 11652 35498
rect 11704 35488 11756 35494
rect 11704 35430 11756 35436
rect 11244 35080 11296 35086
rect 11244 35022 11296 35028
rect 11336 35080 11388 35086
rect 11520 35080 11572 35086
rect 11336 35022 11388 35028
rect 11518 35048 11520 35057
rect 11612 35080 11664 35086
rect 11572 35048 11574 35057
rect 11348 34746 11376 35022
rect 11612 35022 11664 35028
rect 11518 34983 11574 34992
rect 11244 34740 11296 34746
rect 11244 34682 11296 34688
rect 11336 34740 11388 34746
rect 11336 34682 11388 34688
rect 10784 34536 10836 34542
rect 10784 34478 10836 34484
rect 10508 34400 10560 34406
rect 10508 34342 10560 34348
rect 10416 33924 10468 33930
rect 10416 33866 10468 33872
rect 10048 33652 10100 33658
rect 10048 33594 10100 33600
rect 10048 33108 10100 33114
rect 10048 33050 10100 33056
rect 9772 32768 9824 32774
rect 9772 32710 9824 32716
rect 9390 32668 9698 32677
rect 9390 32666 9396 32668
rect 9452 32666 9476 32668
rect 9532 32666 9556 32668
rect 9612 32666 9636 32668
rect 9692 32666 9698 32668
rect 9452 32614 9454 32666
rect 9634 32614 9636 32666
rect 9390 32612 9396 32614
rect 9452 32612 9476 32614
rect 9532 32612 9556 32614
rect 9612 32612 9636 32614
rect 9692 32612 9698 32614
rect 9390 32603 9698 32612
rect 9864 32496 9916 32502
rect 9864 32438 9916 32444
rect 9954 32464 10010 32473
rect 9312 32428 9364 32434
rect 9312 32370 9364 32376
rect 9680 32428 9732 32434
rect 9680 32370 9732 32376
rect 9220 32292 9272 32298
rect 9220 32234 9272 32240
rect 9232 31822 9260 32234
rect 9692 32026 9720 32370
rect 9876 32230 9904 32438
rect 10060 32434 10088 33050
rect 10324 32768 10376 32774
rect 10324 32710 10376 32716
rect 10230 32600 10286 32609
rect 10230 32535 10232 32544
rect 10284 32535 10286 32544
rect 10232 32506 10284 32512
rect 9954 32399 9956 32408
rect 10008 32399 10010 32408
rect 10048 32428 10100 32434
rect 9956 32370 10008 32376
rect 10048 32370 10100 32376
rect 9864 32224 9916 32230
rect 9864 32166 9916 32172
rect 9680 32020 9732 32026
rect 9680 31962 9732 31968
rect 10336 31958 10364 32710
rect 10324 31952 10376 31958
rect 10324 31894 10376 31900
rect 9036 31816 9088 31822
rect 9036 31758 9088 31764
rect 9220 31816 9272 31822
rect 9220 31758 9272 31764
rect 8944 31408 8996 31414
rect 8944 31350 8996 31356
rect 8484 31340 8536 31346
rect 8312 31300 8484 31328
rect 8484 31282 8536 31288
rect 8760 31340 8812 31346
rect 8760 31282 8812 31288
rect 8116 30932 8168 30938
rect 8116 30874 8168 30880
rect 8944 30728 8996 30734
rect 9048 30716 9076 31758
rect 9390 31580 9698 31589
rect 9390 31578 9396 31580
rect 9452 31578 9476 31580
rect 9532 31578 9556 31580
rect 9612 31578 9636 31580
rect 9692 31578 9698 31580
rect 9452 31526 9454 31578
rect 9634 31526 9636 31578
rect 9390 31524 9396 31526
rect 9452 31524 9476 31526
rect 9532 31524 9556 31526
rect 9612 31524 9636 31526
rect 9692 31524 9698 31526
rect 9390 31515 9698 31524
rect 10232 31340 10284 31346
rect 10232 31282 10284 31288
rect 10048 31136 10100 31142
rect 10048 31078 10100 31084
rect 8996 30688 9076 30716
rect 8944 30670 8996 30676
rect 8956 30258 8984 30670
rect 9864 30660 9916 30666
rect 9864 30602 9916 30608
rect 9390 30492 9698 30501
rect 9390 30490 9396 30492
rect 9452 30490 9476 30492
rect 9532 30490 9556 30492
rect 9612 30490 9636 30492
rect 9692 30490 9698 30492
rect 9452 30438 9454 30490
rect 9634 30438 9636 30490
rect 9390 30436 9396 30438
rect 9452 30436 9476 30438
rect 9532 30436 9556 30438
rect 9612 30436 9636 30438
rect 9692 30436 9698 30438
rect 9390 30427 9698 30436
rect 8116 30252 8168 30258
rect 8116 30194 8168 30200
rect 8944 30252 8996 30258
rect 8944 30194 8996 30200
rect 9404 30252 9456 30258
rect 9404 30194 9456 30200
rect 7932 30048 7984 30054
rect 7932 29990 7984 29996
rect 7944 29646 7972 29990
rect 7932 29640 7984 29646
rect 7932 29582 7984 29588
rect 8128 29306 8156 30194
rect 9416 29714 9444 30194
rect 9876 29850 9904 30602
rect 10060 30326 10088 31078
rect 10244 30394 10272 31282
rect 10428 30666 10456 33866
rect 10796 33114 10824 34478
rect 10876 33856 10928 33862
rect 10876 33798 10928 33804
rect 10784 33108 10836 33114
rect 10784 33050 10836 33056
rect 10506 32600 10562 32609
rect 10796 32570 10824 33050
rect 10506 32535 10562 32544
rect 10784 32564 10836 32570
rect 10520 32434 10548 32535
rect 10784 32506 10836 32512
rect 10600 32496 10652 32502
rect 10692 32496 10744 32502
rect 10600 32438 10652 32444
rect 10690 32464 10692 32473
rect 10744 32464 10746 32473
rect 10508 32428 10560 32434
rect 10508 32370 10560 32376
rect 10612 32230 10640 32438
rect 10888 32434 10916 33798
rect 11256 33658 11284 34682
rect 11624 34610 11652 35022
rect 11716 34610 11744 35430
rect 11808 35086 11836 35770
rect 11888 35692 11940 35698
rect 11888 35634 11940 35640
rect 11796 35080 11848 35086
rect 11796 35022 11848 35028
rect 11612 34604 11664 34610
rect 11612 34546 11664 34552
rect 11704 34604 11756 34610
rect 11704 34546 11756 34552
rect 11704 34468 11756 34474
rect 11704 34410 11756 34416
rect 11716 33930 11744 34410
rect 11808 34406 11836 35022
rect 11900 34649 11928 35634
rect 12452 35630 12480 36518
rect 12544 36378 12572 36654
rect 12532 36372 12584 36378
rect 12532 36314 12584 36320
rect 12636 36242 12664 37606
rect 12912 37194 12940 37606
rect 12900 37188 12952 37194
rect 12900 37130 12952 37136
rect 12900 36780 12952 36786
rect 12900 36722 12952 36728
rect 12716 36712 12768 36718
rect 12716 36654 12768 36660
rect 12624 36236 12676 36242
rect 12624 36178 12676 36184
rect 12728 36106 12756 36654
rect 12912 36378 12940 36722
rect 13004 36378 13032 37674
rect 13611 37564 13919 37573
rect 13611 37562 13617 37564
rect 13673 37562 13697 37564
rect 13753 37562 13777 37564
rect 13833 37562 13857 37564
rect 13913 37562 13919 37564
rect 13673 37510 13675 37562
rect 13855 37510 13857 37562
rect 13611 37508 13617 37510
rect 13673 37508 13697 37510
rect 13753 37508 13777 37510
rect 13833 37508 13857 37510
rect 13913 37508 13919 37510
rect 13611 37499 13919 37508
rect 14016 37466 14044 37810
rect 14108 37806 14136 38286
rect 15396 37942 15424 38898
rect 16132 38894 16160 39306
rect 16408 39098 16436 39442
rect 17500 39432 17552 39438
rect 17500 39374 17552 39380
rect 17592 39432 17644 39438
rect 17592 39374 17644 39380
rect 18236 39432 18288 39438
rect 18236 39374 18288 39380
rect 17040 39296 17092 39302
rect 17040 39238 17092 39244
rect 17316 39296 17368 39302
rect 17316 39238 17368 39244
rect 17052 39098 17080 39238
rect 16396 39092 16448 39098
rect 16396 39034 16448 39040
rect 17040 39092 17092 39098
rect 17040 39034 17092 39040
rect 16120 38888 16172 38894
rect 16120 38830 16172 38836
rect 15752 38752 15804 38758
rect 15752 38694 15804 38700
rect 15764 38350 15792 38694
rect 15752 38344 15804 38350
rect 15752 38286 15804 38292
rect 15568 38208 15620 38214
rect 15568 38150 15620 38156
rect 15384 37936 15436 37942
rect 15384 37878 15436 37884
rect 14464 37868 14516 37874
rect 14464 37810 14516 37816
rect 14096 37800 14148 37806
rect 14096 37742 14148 37748
rect 14004 37460 14056 37466
rect 14004 37402 14056 37408
rect 14108 37262 14136 37742
rect 14476 37466 14504 37810
rect 14464 37460 14516 37466
rect 14464 37402 14516 37408
rect 14096 37256 14148 37262
rect 14096 37198 14148 37204
rect 14372 37256 14424 37262
rect 14372 37198 14424 37204
rect 13084 37188 13136 37194
rect 13084 37130 13136 37136
rect 12900 36372 12952 36378
rect 12900 36314 12952 36320
rect 12992 36372 13044 36378
rect 12992 36314 13044 36320
rect 12716 36100 12768 36106
rect 12716 36042 12768 36048
rect 12532 36032 12584 36038
rect 12532 35974 12584 35980
rect 12544 35834 12572 35974
rect 12532 35828 12584 35834
rect 12532 35770 12584 35776
rect 12440 35624 12492 35630
rect 12440 35566 12492 35572
rect 12624 35012 12676 35018
rect 12624 34954 12676 34960
rect 12256 34944 12308 34950
rect 12308 34892 12572 34898
rect 12256 34886 12572 34892
rect 12268 34870 12572 34886
rect 12544 34746 12572 34870
rect 12532 34740 12584 34746
rect 12532 34682 12584 34688
rect 11886 34640 11942 34649
rect 11886 34575 11942 34584
rect 11796 34400 11848 34406
rect 11796 34342 11848 34348
rect 12164 34400 12216 34406
rect 12164 34342 12216 34348
rect 11980 33992 12032 33998
rect 11980 33934 12032 33940
rect 11704 33924 11756 33930
rect 11704 33866 11756 33872
rect 11244 33652 11296 33658
rect 11244 33594 11296 33600
rect 11520 33312 11572 33318
rect 11520 33254 11572 33260
rect 11532 32910 11560 33254
rect 11520 32904 11572 32910
rect 11440 32864 11520 32892
rect 11336 32768 11388 32774
rect 11336 32710 11388 32716
rect 11152 32496 11204 32502
rect 11152 32438 11204 32444
rect 10690 32399 10746 32408
rect 10876 32428 10928 32434
rect 10876 32370 10928 32376
rect 10600 32224 10652 32230
rect 10600 32166 10652 32172
rect 11164 32026 11192 32438
rect 11060 32020 11112 32026
rect 11060 31962 11112 31968
rect 11152 32020 11204 32026
rect 11152 31962 11204 31968
rect 11072 31346 11100 31962
rect 11348 31754 11376 32710
rect 11440 32230 11468 32864
rect 11520 32846 11572 32852
rect 11520 32768 11572 32774
rect 11520 32710 11572 32716
rect 11532 32570 11560 32710
rect 11520 32564 11572 32570
rect 11520 32506 11572 32512
rect 11428 32224 11480 32230
rect 11428 32166 11480 32172
rect 11336 31748 11388 31754
rect 11336 31690 11388 31696
rect 11060 31340 11112 31346
rect 11060 31282 11112 31288
rect 11612 31340 11664 31346
rect 11612 31282 11664 31288
rect 11796 31340 11848 31346
rect 11796 31282 11848 31288
rect 10508 31272 10560 31278
rect 10508 31214 10560 31220
rect 10520 30938 10548 31214
rect 11152 31136 11204 31142
rect 11152 31078 11204 31084
rect 10508 30932 10560 30938
rect 10508 30874 10560 30880
rect 10416 30660 10468 30666
rect 10416 30602 10468 30608
rect 10232 30388 10284 30394
rect 10232 30330 10284 30336
rect 10048 30320 10100 30326
rect 10048 30262 10100 30268
rect 9864 29844 9916 29850
rect 9864 29786 9916 29792
rect 10232 29776 10284 29782
rect 10232 29718 10284 29724
rect 8852 29708 8904 29714
rect 8852 29650 8904 29656
rect 9404 29708 9456 29714
rect 9404 29650 9456 29656
rect 8484 29504 8536 29510
rect 8484 29446 8536 29452
rect 8116 29300 8168 29306
rect 8116 29242 8168 29248
rect 8116 29164 8168 29170
rect 8116 29106 8168 29112
rect 8128 28558 8156 29106
rect 8496 29102 8524 29446
rect 8864 29238 8892 29650
rect 9312 29640 9364 29646
rect 9312 29582 9364 29588
rect 8944 29504 8996 29510
rect 8944 29446 8996 29452
rect 8956 29306 8984 29446
rect 9324 29306 9352 29582
rect 9390 29404 9698 29413
rect 9390 29402 9396 29404
rect 9452 29402 9476 29404
rect 9532 29402 9556 29404
rect 9612 29402 9636 29404
rect 9692 29402 9698 29404
rect 9452 29350 9454 29402
rect 9634 29350 9636 29402
rect 9390 29348 9396 29350
rect 9452 29348 9476 29350
rect 9532 29348 9556 29350
rect 9612 29348 9636 29350
rect 9692 29348 9698 29350
rect 9390 29339 9698 29348
rect 8944 29300 8996 29306
rect 8944 29242 8996 29248
rect 9312 29300 9364 29306
rect 9312 29242 9364 29248
rect 9772 29300 9824 29306
rect 9772 29242 9824 29248
rect 8852 29232 8904 29238
rect 8852 29174 8904 29180
rect 9220 29232 9272 29238
rect 9220 29174 9272 29180
rect 8484 29096 8536 29102
rect 8484 29038 8536 29044
rect 8300 28960 8352 28966
rect 8300 28902 8352 28908
rect 8312 28626 8340 28902
rect 8300 28620 8352 28626
rect 8300 28562 8352 28568
rect 8496 28558 8524 29038
rect 8116 28552 8168 28558
rect 8116 28494 8168 28500
rect 8208 28552 8260 28558
rect 8208 28494 8260 28500
rect 8484 28552 8536 28558
rect 8484 28494 8536 28500
rect 8220 28218 8248 28494
rect 8208 28212 8260 28218
rect 8208 28154 8260 28160
rect 8864 27130 8892 29174
rect 8944 28620 8996 28626
rect 8944 28562 8996 28568
rect 8956 27946 8984 28562
rect 9232 28490 9260 29174
rect 9324 29034 9352 29242
rect 9496 29164 9548 29170
rect 9496 29106 9548 29112
rect 9312 29028 9364 29034
rect 9312 28970 9364 28976
rect 9324 28762 9352 28970
rect 9312 28756 9364 28762
rect 9312 28698 9364 28704
rect 9508 28626 9536 29106
rect 9496 28620 9548 28626
rect 9496 28562 9548 28568
rect 9220 28484 9272 28490
rect 9220 28426 9272 28432
rect 9036 28416 9088 28422
rect 9036 28358 9088 28364
rect 8944 27940 8996 27946
rect 8944 27882 8996 27888
rect 8852 27124 8904 27130
rect 8852 27066 8904 27072
rect 9048 26994 9076 28358
rect 9232 28082 9260 28426
rect 9390 28316 9698 28325
rect 9390 28314 9396 28316
rect 9452 28314 9476 28316
rect 9532 28314 9556 28316
rect 9612 28314 9636 28316
rect 9692 28314 9698 28316
rect 9452 28262 9454 28314
rect 9634 28262 9636 28314
rect 9390 28260 9396 28262
rect 9452 28260 9476 28262
rect 9532 28260 9556 28262
rect 9612 28260 9636 28262
rect 9692 28260 9698 28262
rect 9390 28251 9698 28260
rect 9220 28076 9272 28082
rect 9220 28018 9272 28024
rect 9232 27674 9260 28018
rect 9220 27668 9272 27674
rect 9220 27610 9272 27616
rect 9784 27402 9812 29242
rect 10048 29164 10100 29170
rect 10048 29106 10100 29112
rect 9956 29028 10008 29034
rect 9956 28970 10008 28976
rect 9864 28620 9916 28626
rect 9864 28562 9916 28568
rect 9876 28014 9904 28562
rect 9968 28558 9996 28970
rect 9956 28552 10008 28558
rect 9956 28494 10008 28500
rect 9956 28416 10008 28422
rect 9956 28358 10008 28364
rect 9968 28218 9996 28358
rect 9956 28212 10008 28218
rect 9956 28154 10008 28160
rect 9864 28008 9916 28014
rect 9864 27950 9916 27956
rect 9876 27470 9904 27950
rect 9864 27464 9916 27470
rect 9864 27406 9916 27412
rect 9772 27396 9824 27402
rect 9772 27338 9824 27344
rect 9390 27228 9698 27237
rect 9390 27226 9396 27228
rect 9452 27226 9476 27228
rect 9532 27226 9556 27228
rect 9612 27226 9636 27228
rect 9692 27226 9698 27228
rect 9452 27174 9454 27226
rect 9634 27174 9636 27226
rect 9390 27172 9396 27174
rect 9452 27172 9476 27174
rect 9532 27172 9556 27174
rect 9612 27172 9636 27174
rect 9692 27172 9698 27174
rect 9390 27163 9698 27172
rect 9036 26988 9088 26994
rect 9036 26930 9088 26936
rect 9876 26382 9904 27406
rect 10060 27130 10088 29106
rect 10244 28966 10272 29718
rect 10324 29164 10376 29170
rect 10324 29106 10376 29112
rect 10232 28960 10284 28966
rect 10232 28902 10284 28908
rect 10244 28558 10272 28902
rect 10336 28558 10364 29106
rect 10232 28552 10284 28558
rect 10232 28494 10284 28500
rect 10324 28552 10376 28558
rect 10324 28494 10376 28500
rect 10048 27124 10100 27130
rect 10048 27066 10100 27072
rect 8300 26376 8352 26382
rect 8300 26318 8352 26324
rect 9864 26376 9916 26382
rect 9864 26318 9916 26324
rect 8312 26042 8340 26318
rect 9390 26140 9698 26149
rect 9390 26138 9396 26140
rect 9452 26138 9476 26140
rect 9532 26138 9556 26140
rect 9612 26138 9636 26140
rect 9692 26138 9698 26140
rect 9452 26086 9454 26138
rect 9634 26086 9636 26138
rect 9390 26084 9396 26086
rect 9452 26084 9476 26086
rect 9532 26084 9556 26086
rect 9612 26084 9636 26086
rect 9692 26084 9698 26086
rect 9390 26075 9698 26084
rect 8300 26036 8352 26042
rect 8300 25978 8352 25984
rect 10428 25906 10456 30602
rect 11164 30122 11192 31078
rect 11520 30252 11572 30258
rect 11520 30194 11572 30200
rect 11152 30116 11204 30122
rect 11152 30058 11204 30064
rect 10968 30048 11020 30054
rect 10968 29990 11020 29996
rect 10980 29782 11008 29990
rect 10968 29776 11020 29782
rect 10968 29718 11020 29724
rect 10692 29504 10744 29510
rect 10692 29446 10744 29452
rect 10784 29504 10836 29510
rect 10784 29446 10836 29452
rect 10508 28960 10560 28966
rect 10508 28902 10560 28908
rect 10600 28960 10652 28966
rect 10600 28902 10652 28908
rect 10520 28762 10548 28902
rect 10508 28756 10560 28762
rect 10508 28698 10560 28704
rect 10612 28422 10640 28902
rect 10704 28762 10732 29446
rect 10796 29170 10824 29446
rect 10784 29164 10836 29170
rect 10784 29106 10836 29112
rect 10692 28756 10744 28762
rect 10692 28698 10744 28704
rect 10796 28558 10824 29106
rect 10876 29096 10928 29102
rect 10876 29038 10928 29044
rect 10980 29050 11008 29718
rect 11532 29306 11560 30194
rect 11520 29300 11572 29306
rect 11520 29242 11572 29248
rect 11244 29096 11296 29102
rect 10980 29044 11244 29050
rect 10980 29038 11296 29044
rect 10888 28558 10916 29038
rect 10980 29022 11284 29038
rect 11624 28762 11652 31282
rect 11704 30048 11756 30054
rect 11704 29990 11756 29996
rect 11612 28756 11664 28762
rect 11612 28698 11664 28704
rect 11716 28558 11744 29990
rect 11808 29306 11836 31282
rect 11992 29850 12020 33934
rect 12176 33862 12204 34342
rect 12544 34082 12572 34682
rect 12452 34054 12572 34082
rect 12164 33856 12216 33862
rect 12164 33798 12216 33804
rect 12256 33856 12308 33862
rect 12256 33798 12308 33804
rect 12176 33590 12204 33798
rect 12164 33584 12216 33590
rect 12164 33526 12216 33532
rect 12268 32978 12296 33798
rect 12256 32972 12308 32978
rect 12256 32914 12308 32920
rect 12256 31884 12308 31890
rect 12256 31826 12308 31832
rect 12072 30592 12124 30598
rect 12072 30534 12124 30540
rect 11980 29844 12032 29850
rect 11980 29786 12032 29792
rect 11796 29300 11848 29306
rect 11796 29242 11848 29248
rect 11992 28994 12020 29786
rect 12084 29646 12112 30534
rect 12072 29640 12124 29646
rect 12072 29582 12124 29588
rect 12164 29640 12216 29646
rect 12164 29582 12216 29588
rect 11900 28966 12020 28994
rect 11796 28960 11848 28966
rect 11796 28902 11848 28908
rect 10784 28552 10836 28558
rect 10784 28494 10836 28500
rect 10876 28552 10928 28558
rect 10876 28494 10928 28500
rect 11704 28552 11756 28558
rect 11704 28494 11756 28500
rect 10600 28416 10652 28422
rect 10600 28358 10652 28364
rect 10612 28218 10640 28358
rect 10600 28212 10652 28218
rect 10600 28154 10652 28160
rect 10888 27674 10916 28494
rect 11520 28484 11572 28490
rect 11520 28426 11572 28432
rect 11532 28218 11560 28426
rect 11704 28416 11756 28422
rect 11704 28358 11756 28364
rect 11520 28212 11572 28218
rect 11520 28154 11572 28160
rect 10876 27668 10928 27674
rect 10876 27610 10928 27616
rect 11716 27062 11744 28358
rect 11808 28082 11836 28902
rect 11900 28218 11928 28966
rect 12176 28762 12204 29582
rect 12268 29238 12296 31826
rect 12348 31680 12400 31686
rect 12348 31622 12400 31628
rect 12360 31346 12388 31622
rect 12452 31346 12480 34054
rect 12532 33992 12584 33998
rect 12532 33934 12584 33940
rect 12544 33114 12572 33934
rect 12636 33522 12664 34954
rect 12728 34950 12756 36042
rect 13096 36038 13124 37130
rect 13268 37120 13320 37126
rect 13268 37062 13320 37068
rect 13280 36922 13308 37062
rect 13268 36916 13320 36922
rect 13268 36858 13320 36864
rect 13176 36576 13228 36582
rect 13176 36518 13228 36524
rect 13084 36032 13136 36038
rect 13084 35974 13136 35980
rect 13188 35834 13216 36518
rect 13280 36378 13308 36858
rect 13452 36712 13504 36718
rect 13452 36654 13504 36660
rect 13360 36576 13412 36582
rect 13360 36518 13412 36524
rect 13372 36378 13400 36518
rect 13268 36372 13320 36378
rect 13268 36314 13320 36320
rect 13360 36372 13412 36378
rect 13360 36314 13412 36320
rect 13464 35834 13492 36654
rect 13611 36476 13919 36485
rect 13611 36474 13617 36476
rect 13673 36474 13697 36476
rect 13753 36474 13777 36476
rect 13833 36474 13857 36476
rect 13913 36474 13919 36476
rect 13673 36422 13675 36474
rect 13855 36422 13857 36474
rect 13611 36420 13617 36422
rect 13673 36420 13697 36422
rect 13753 36420 13777 36422
rect 13833 36420 13857 36422
rect 13913 36420 13919 36422
rect 13611 36411 13919 36420
rect 14108 36174 14136 37198
rect 14384 36922 14412 37198
rect 15396 37126 15424 37878
rect 15580 37398 15608 38150
rect 16132 37738 16160 38830
rect 17040 38752 17092 38758
rect 17040 38694 17092 38700
rect 17052 38350 17080 38694
rect 17040 38344 17092 38350
rect 17040 38286 17092 38292
rect 16120 37732 16172 37738
rect 16120 37674 16172 37680
rect 15568 37392 15620 37398
rect 15568 37334 15620 37340
rect 17052 37126 17080 38286
rect 17224 37664 17276 37670
rect 17224 37606 17276 37612
rect 15384 37120 15436 37126
rect 15384 37062 15436 37068
rect 16304 37120 16356 37126
rect 16304 37062 16356 37068
rect 16948 37120 17000 37126
rect 16948 37062 17000 37068
rect 17040 37120 17092 37126
rect 17040 37062 17092 37068
rect 14372 36916 14424 36922
rect 14372 36858 14424 36864
rect 14648 36576 14700 36582
rect 14648 36518 14700 36524
rect 14660 36174 14688 36518
rect 14096 36168 14148 36174
rect 14096 36110 14148 36116
rect 14648 36168 14700 36174
rect 14648 36110 14700 36116
rect 13636 36032 13688 36038
rect 13636 35974 13688 35980
rect 14556 36032 14608 36038
rect 14556 35974 14608 35980
rect 13648 35834 13676 35974
rect 13176 35828 13228 35834
rect 13176 35770 13228 35776
rect 13452 35828 13504 35834
rect 13452 35770 13504 35776
rect 13636 35828 13688 35834
rect 13636 35770 13688 35776
rect 12992 35692 13044 35698
rect 12992 35634 13044 35640
rect 14096 35692 14148 35698
rect 14096 35634 14148 35640
rect 13004 35494 13032 35634
rect 13360 35624 13412 35630
rect 13360 35566 13412 35572
rect 13084 35556 13136 35562
rect 13084 35498 13136 35504
rect 12992 35488 13044 35494
rect 12992 35430 13044 35436
rect 12900 35148 12952 35154
rect 13004 35136 13032 35430
rect 12952 35108 13032 35136
rect 12900 35090 12952 35096
rect 12716 34944 12768 34950
rect 12716 34886 12768 34892
rect 12992 34740 13044 34746
rect 12992 34682 13044 34688
rect 13004 34610 13032 34682
rect 13096 34678 13124 35498
rect 13372 34746 13400 35566
rect 13611 35388 13919 35397
rect 13611 35386 13617 35388
rect 13673 35386 13697 35388
rect 13753 35386 13777 35388
rect 13833 35386 13857 35388
rect 13913 35386 13919 35388
rect 13673 35334 13675 35386
rect 13855 35334 13857 35386
rect 13611 35332 13617 35334
rect 13673 35332 13697 35334
rect 13753 35332 13777 35334
rect 13833 35332 13857 35334
rect 13913 35332 13919 35334
rect 13611 35323 13919 35332
rect 14004 35080 14056 35086
rect 14004 35022 14056 35028
rect 13360 34740 13412 34746
rect 13360 34682 13412 34688
rect 13084 34672 13136 34678
rect 13084 34614 13136 34620
rect 12992 34604 13044 34610
rect 12992 34546 13044 34552
rect 13096 34134 13124 34614
rect 13360 34400 13412 34406
rect 13360 34342 13412 34348
rect 13084 34128 13136 34134
rect 13084 34070 13136 34076
rect 13372 34082 13400 34342
rect 13611 34300 13919 34309
rect 13611 34298 13617 34300
rect 13673 34298 13697 34300
rect 13753 34298 13777 34300
rect 13833 34298 13857 34300
rect 13913 34298 13919 34300
rect 13673 34246 13675 34298
rect 13855 34246 13857 34298
rect 13611 34244 13617 34246
rect 13673 34244 13697 34246
rect 13753 34244 13777 34246
rect 13833 34244 13857 34246
rect 13913 34244 13919 34246
rect 13611 34235 13919 34244
rect 13372 34066 13492 34082
rect 13372 34060 13504 34066
rect 13372 34054 13452 34060
rect 13452 34002 13504 34008
rect 12624 33516 12676 33522
rect 12624 33458 12676 33464
rect 13360 33448 13412 33454
rect 13360 33390 13412 33396
rect 12716 33312 12768 33318
rect 12716 33254 12768 33260
rect 13084 33312 13136 33318
rect 13084 33254 13136 33260
rect 12532 33108 12584 33114
rect 12532 33050 12584 33056
rect 12728 32774 12756 33254
rect 13096 32910 13124 33254
rect 13084 32904 13136 32910
rect 13084 32846 13136 32852
rect 12716 32768 12768 32774
rect 12716 32710 12768 32716
rect 12728 32230 12756 32710
rect 13372 32570 13400 33390
rect 13464 33266 13492 34002
rect 14016 33998 14044 35022
rect 14108 34474 14136 35634
rect 14568 35562 14596 35974
rect 14556 35556 14608 35562
rect 14556 35498 14608 35504
rect 14568 35154 14596 35498
rect 14740 35488 14792 35494
rect 14740 35430 14792 35436
rect 14556 35148 14608 35154
rect 14556 35090 14608 35096
rect 14752 34610 14780 35430
rect 15016 35012 15068 35018
rect 15016 34954 15068 34960
rect 15028 34746 15056 34954
rect 15108 34944 15160 34950
rect 15108 34886 15160 34892
rect 15016 34740 15068 34746
rect 15016 34682 15068 34688
rect 14740 34604 14792 34610
rect 14740 34546 14792 34552
rect 14096 34468 14148 34474
rect 14096 34410 14148 34416
rect 15120 34406 15148 34886
rect 15198 34640 15254 34649
rect 15198 34575 15254 34584
rect 14924 34400 14976 34406
rect 14924 34342 14976 34348
rect 15108 34400 15160 34406
rect 15108 34342 15160 34348
rect 14936 34202 14964 34342
rect 14096 34196 14148 34202
rect 14096 34138 14148 34144
rect 14924 34196 14976 34202
rect 14924 34138 14976 34144
rect 13820 33992 13872 33998
rect 13820 33934 13872 33940
rect 14004 33992 14056 33998
rect 14004 33934 14056 33940
rect 13728 33856 13780 33862
rect 13728 33798 13780 33804
rect 13740 33658 13768 33798
rect 13728 33652 13780 33658
rect 13728 33594 13780 33600
rect 13832 33590 13860 33934
rect 14004 33856 14056 33862
rect 14004 33798 14056 33804
rect 13820 33584 13872 33590
rect 13820 33526 13872 33532
rect 13544 33516 13596 33522
rect 13544 33458 13596 33464
rect 13556 33266 13584 33458
rect 13464 33238 13584 33266
rect 13360 32564 13412 32570
rect 13360 32506 13412 32512
rect 13464 32502 13492 33238
rect 13611 33212 13919 33221
rect 13611 33210 13617 33212
rect 13673 33210 13697 33212
rect 13753 33210 13777 33212
rect 13833 33210 13857 33212
rect 13913 33210 13919 33212
rect 13673 33158 13675 33210
rect 13855 33158 13857 33210
rect 13611 33156 13617 33158
rect 13673 33156 13697 33158
rect 13753 33156 13777 33158
rect 13833 33156 13857 33158
rect 13913 33156 13919 33158
rect 13611 33147 13919 33156
rect 14016 32570 14044 33798
rect 14108 33114 14136 34138
rect 14556 34060 14608 34066
rect 14556 34002 14608 34008
rect 14188 33924 14240 33930
rect 14188 33866 14240 33872
rect 14372 33924 14424 33930
rect 14372 33866 14424 33872
rect 14096 33108 14148 33114
rect 14096 33050 14148 33056
rect 14004 32564 14056 32570
rect 14004 32506 14056 32512
rect 13452 32496 13504 32502
rect 13452 32438 13504 32444
rect 12716 32224 12768 32230
rect 12716 32166 12768 32172
rect 12728 31822 12756 32166
rect 13464 31822 13492 32438
rect 14200 32434 14228 33866
rect 14280 33652 14332 33658
rect 14280 33594 14332 33600
rect 14292 32910 14320 33594
rect 14384 33318 14412 33866
rect 14464 33448 14516 33454
rect 14464 33390 14516 33396
rect 14372 33312 14424 33318
rect 14372 33254 14424 33260
rect 14476 32978 14504 33390
rect 14464 32972 14516 32978
rect 14464 32914 14516 32920
rect 14280 32904 14332 32910
rect 14280 32846 14332 32852
rect 14096 32428 14148 32434
rect 14016 32388 14096 32416
rect 14016 32337 14044 32388
rect 14096 32370 14148 32376
rect 14188 32428 14240 32434
rect 14188 32370 14240 32376
rect 14002 32328 14058 32337
rect 14002 32263 14058 32272
rect 14096 32292 14148 32298
rect 14096 32234 14148 32240
rect 13611 32124 13919 32133
rect 13611 32122 13617 32124
rect 13673 32122 13697 32124
rect 13753 32122 13777 32124
rect 13833 32122 13857 32124
rect 13913 32122 13919 32124
rect 13673 32070 13675 32122
rect 13855 32070 13857 32122
rect 13611 32068 13617 32070
rect 13673 32068 13697 32070
rect 13753 32068 13777 32070
rect 13833 32068 13857 32070
rect 13913 32068 13919 32070
rect 13611 32059 13919 32068
rect 14108 32026 14136 32234
rect 14096 32020 14148 32026
rect 14096 31962 14148 31968
rect 13820 31884 13872 31890
rect 13820 31826 13872 31832
rect 12716 31816 12768 31822
rect 12716 31758 12768 31764
rect 13452 31816 13504 31822
rect 13452 31758 13504 31764
rect 12348 31340 12400 31346
rect 12348 31282 12400 31288
rect 12440 31340 12492 31346
rect 12440 31282 12492 31288
rect 12728 31278 12756 31758
rect 13268 31680 13320 31686
rect 13268 31622 13320 31628
rect 13280 31414 13308 31622
rect 13832 31482 13860 31826
rect 14200 31822 14228 32370
rect 14280 32360 14332 32366
rect 14280 32302 14332 32308
rect 14096 31816 14148 31822
rect 14016 31764 14096 31770
rect 14016 31758 14148 31764
rect 14188 31816 14240 31822
rect 14188 31758 14240 31764
rect 14016 31742 14136 31758
rect 13820 31476 13872 31482
rect 13820 31418 13872 31424
rect 13268 31408 13320 31414
rect 13268 31350 13320 31356
rect 14016 31346 14044 31742
rect 13360 31340 13412 31346
rect 13360 31282 13412 31288
rect 14004 31340 14056 31346
rect 14004 31282 14056 31288
rect 12716 31272 12768 31278
rect 12716 31214 12768 31220
rect 12532 31136 12584 31142
rect 12532 31078 12584 31084
rect 12544 30734 12572 31078
rect 12728 30802 12756 31214
rect 12716 30796 12768 30802
rect 12716 30738 12768 30744
rect 12532 30728 12584 30734
rect 12532 30670 12584 30676
rect 12728 30258 12756 30738
rect 13372 30734 13400 31282
rect 14200 31142 14228 31758
rect 14292 31686 14320 32302
rect 14372 32224 14424 32230
rect 14372 32166 14424 32172
rect 14280 31680 14332 31686
rect 14280 31622 14332 31628
rect 14292 31414 14320 31622
rect 14280 31408 14332 31414
rect 14280 31350 14332 31356
rect 14384 31346 14412 32166
rect 14476 31346 14504 32914
rect 14568 32230 14596 34002
rect 14936 33522 14964 34138
rect 15016 33856 15068 33862
rect 15016 33798 15068 33804
rect 14740 33516 14792 33522
rect 14740 33458 14792 33464
rect 14924 33516 14976 33522
rect 14924 33458 14976 33464
rect 14752 33114 14780 33458
rect 14936 33402 14964 33458
rect 14844 33374 14964 33402
rect 14740 33108 14792 33114
rect 14740 33050 14792 33056
rect 14844 33017 14872 33374
rect 14924 33312 14976 33318
rect 14924 33254 14976 33260
rect 14830 33008 14886 33017
rect 14740 32972 14792 32978
rect 14830 32943 14886 32952
rect 14740 32914 14792 32920
rect 14648 32904 14700 32910
rect 14648 32846 14700 32852
rect 14660 32570 14688 32846
rect 14752 32570 14780 32914
rect 14832 32836 14884 32842
rect 14832 32778 14884 32784
rect 14844 32570 14872 32778
rect 14648 32564 14700 32570
rect 14648 32506 14700 32512
rect 14740 32564 14792 32570
rect 14740 32506 14792 32512
rect 14832 32564 14884 32570
rect 14832 32506 14884 32512
rect 14556 32224 14608 32230
rect 14556 32166 14608 32172
rect 14660 31958 14688 32506
rect 14738 32464 14794 32473
rect 14936 32450 14964 33254
rect 14844 32434 14964 32450
rect 15028 32434 15056 33798
rect 14738 32399 14794 32408
rect 14832 32428 14964 32434
rect 14648 31952 14700 31958
rect 14648 31894 14700 31900
rect 14556 31476 14608 31482
rect 14556 31418 14608 31424
rect 14372 31340 14424 31346
rect 14372 31282 14424 31288
rect 14464 31340 14516 31346
rect 14464 31282 14516 31288
rect 13452 31136 13504 31142
rect 13452 31078 13504 31084
rect 14188 31136 14240 31142
rect 14188 31078 14240 31084
rect 13464 30734 13492 31078
rect 13611 31036 13919 31045
rect 13611 31034 13617 31036
rect 13673 31034 13697 31036
rect 13753 31034 13777 31036
rect 13833 31034 13857 31036
rect 13913 31034 13919 31036
rect 13673 30982 13675 31034
rect 13855 30982 13857 31034
rect 13611 30980 13617 30982
rect 13673 30980 13697 30982
rect 13753 30980 13777 30982
rect 13833 30980 13857 30982
rect 13913 30980 13919 30982
rect 13611 30971 13919 30980
rect 13360 30728 13412 30734
rect 13360 30670 13412 30676
rect 13452 30728 13504 30734
rect 13452 30670 13504 30676
rect 12716 30252 12768 30258
rect 12716 30194 12768 30200
rect 12728 29850 12756 30194
rect 13268 30048 13320 30054
rect 13268 29990 13320 29996
rect 12716 29844 12768 29850
rect 12716 29786 12768 29792
rect 12440 29572 12492 29578
rect 12440 29514 12492 29520
rect 12348 29504 12400 29510
rect 12348 29446 12400 29452
rect 12256 29232 12308 29238
rect 12256 29174 12308 29180
rect 12164 28756 12216 28762
rect 12164 28698 12216 28704
rect 11888 28212 11940 28218
rect 11888 28154 11940 28160
rect 11796 28076 11848 28082
rect 11796 28018 11848 28024
rect 12268 27946 12296 29174
rect 12360 29034 12388 29446
rect 12348 29028 12400 29034
rect 12348 28970 12400 28976
rect 12360 28150 12388 28970
rect 12348 28144 12400 28150
rect 12348 28086 12400 28092
rect 12256 27940 12308 27946
rect 12256 27882 12308 27888
rect 12452 27538 12480 29514
rect 13280 29238 13308 29990
rect 13372 29646 13400 30670
rect 14200 30666 14228 31078
rect 14476 30734 14504 31282
rect 14464 30728 14516 30734
rect 14464 30670 14516 30676
rect 14568 30666 14596 31418
rect 14660 31346 14688 31894
rect 14752 31686 14780 32399
rect 14884 32422 14964 32428
rect 15016 32428 15068 32434
rect 14832 32370 14884 32376
rect 15016 32370 15068 32376
rect 14844 32026 14872 32370
rect 15120 32366 15148 34342
rect 15108 32360 15160 32366
rect 15108 32302 15160 32308
rect 14832 32020 14884 32026
rect 14832 31962 14884 31968
rect 14740 31680 14792 31686
rect 14740 31622 14792 31628
rect 14844 31346 15056 31362
rect 14648 31340 14700 31346
rect 14648 31282 14700 31288
rect 14844 31340 15068 31346
rect 14844 31334 15016 31340
rect 14648 31204 14700 31210
rect 14648 31146 14700 31152
rect 14188 30660 14240 30666
rect 14188 30602 14240 30608
rect 14556 30660 14608 30666
rect 14556 30602 14608 30608
rect 14096 30592 14148 30598
rect 14096 30534 14148 30540
rect 14280 30592 14332 30598
rect 14280 30534 14332 30540
rect 14108 30326 14136 30534
rect 14096 30320 14148 30326
rect 14096 30262 14148 30268
rect 14004 30184 14056 30190
rect 14292 30138 14320 30534
rect 14568 30190 14596 30602
rect 14660 30394 14688 31146
rect 14844 31090 14872 31334
rect 15016 31282 15068 31288
rect 14752 31062 14872 31090
rect 15016 31136 15068 31142
rect 15016 31078 15068 31084
rect 14752 30734 14780 31062
rect 15028 30870 15056 31078
rect 15016 30864 15068 30870
rect 15016 30806 15068 30812
rect 14740 30728 14792 30734
rect 14740 30670 14792 30676
rect 14648 30388 14700 30394
rect 14648 30330 14700 30336
rect 14056 30132 14320 30138
rect 14004 30126 14320 30132
rect 14556 30184 14608 30190
rect 14556 30126 14608 30132
rect 14016 30110 14320 30126
rect 14004 30048 14056 30054
rect 14004 29990 14056 29996
rect 13611 29948 13919 29957
rect 13611 29946 13617 29948
rect 13673 29946 13697 29948
rect 13753 29946 13777 29948
rect 13833 29946 13857 29948
rect 13913 29946 13919 29948
rect 13673 29894 13675 29946
rect 13855 29894 13857 29946
rect 13611 29892 13617 29894
rect 13673 29892 13697 29894
rect 13753 29892 13777 29894
rect 13833 29892 13857 29894
rect 13913 29892 13919 29894
rect 13611 29883 13919 29892
rect 13360 29640 13412 29646
rect 13360 29582 13412 29588
rect 13372 29306 13400 29582
rect 14016 29306 14044 29990
rect 14200 29306 14228 30110
rect 14740 30048 14792 30054
rect 14740 29990 14792 29996
rect 14752 29646 14780 29990
rect 14740 29640 14792 29646
rect 14740 29582 14792 29588
rect 14464 29504 14516 29510
rect 14464 29446 14516 29452
rect 14476 29306 14504 29446
rect 13360 29300 13412 29306
rect 13360 29242 13412 29248
rect 14004 29300 14056 29306
rect 14004 29242 14056 29248
rect 14188 29300 14240 29306
rect 14188 29242 14240 29248
rect 14464 29300 14516 29306
rect 14464 29242 14516 29248
rect 13268 29232 13320 29238
rect 13268 29174 13320 29180
rect 14740 29232 14792 29238
rect 14740 29174 14792 29180
rect 13176 29164 13228 29170
rect 13176 29106 13228 29112
rect 12716 28960 12768 28966
rect 12716 28902 12768 28908
rect 12900 28960 12952 28966
rect 12900 28902 12952 28908
rect 12728 28506 12756 28902
rect 12912 28626 12940 28902
rect 13188 28762 13216 29106
rect 13176 28756 13228 28762
rect 13176 28698 13228 28704
rect 12900 28620 12952 28626
rect 12900 28562 12952 28568
rect 12808 28552 12860 28558
rect 12728 28500 12808 28506
rect 12728 28494 12860 28500
rect 12728 28478 12848 28494
rect 12728 28082 12756 28478
rect 12716 28076 12768 28082
rect 12716 28018 12768 28024
rect 12912 28014 12940 28562
rect 13188 28082 13216 28698
rect 13176 28076 13228 28082
rect 13176 28018 13228 28024
rect 13280 28014 13308 29174
rect 14372 29164 14424 29170
rect 14372 29106 14424 29112
rect 14096 29028 14148 29034
rect 14096 28970 14148 28976
rect 13611 28860 13919 28869
rect 13611 28858 13617 28860
rect 13673 28858 13697 28860
rect 13753 28858 13777 28860
rect 13833 28858 13857 28860
rect 13913 28858 13919 28860
rect 13673 28806 13675 28858
rect 13855 28806 13857 28858
rect 13611 28804 13617 28806
rect 13673 28804 13697 28806
rect 13753 28804 13777 28806
rect 13833 28804 13857 28806
rect 13913 28804 13919 28806
rect 13611 28795 13919 28804
rect 13360 28620 13412 28626
rect 13360 28562 13412 28568
rect 13372 28218 13400 28562
rect 13544 28552 13596 28558
rect 13544 28494 13596 28500
rect 13556 28218 13584 28494
rect 13912 28484 13964 28490
rect 13912 28426 13964 28432
rect 13360 28212 13412 28218
rect 13360 28154 13412 28160
rect 13544 28212 13596 28218
rect 13544 28154 13596 28160
rect 13924 28082 13952 28426
rect 13912 28076 13964 28082
rect 13912 28018 13964 28024
rect 12900 28008 12952 28014
rect 12900 27950 12952 27956
rect 13268 28008 13320 28014
rect 13268 27950 13320 27956
rect 13924 27928 13952 28018
rect 13924 27900 14044 27928
rect 13452 27872 13504 27878
rect 13452 27814 13504 27820
rect 12440 27532 12492 27538
rect 12440 27474 12492 27480
rect 13084 27532 13136 27538
rect 13084 27474 13136 27480
rect 12256 27464 12308 27470
rect 12256 27406 12308 27412
rect 11980 27124 12032 27130
rect 11980 27066 12032 27072
rect 11704 27056 11756 27062
rect 11704 26998 11756 27004
rect 11152 26988 11204 26994
rect 11152 26930 11204 26936
rect 10692 26308 10744 26314
rect 10692 26250 10744 26256
rect 10704 25974 10732 26250
rect 10692 25968 10744 25974
rect 10692 25910 10744 25916
rect 10416 25900 10468 25906
rect 10416 25842 10468 25848
rect 10232 25424 10284 25430
rect 10232 25366 10284 25372
rect 10140 25356 10192 25362
rect 10140 25298 10192 25304
rect 9390 25052 9698 25061
rect 9390 25050 9396 25052
rect 9452 25050 9476 25052
rect 9532 25050 9556 25052
rect 9612 25050 9636 25052
rect 9692 25050 9698 25052
rect 9452 24998 9454 25050
rect 9634 24998 9636 25050
rect 9390 24996 9396 24998
rect 9452 24996 9476 24998
rect 9532 24996 9556 24998
rect 9612 24996 9636 24998
rect 9692 24996 9698 24998
rect 9390 24987 9698 24996
rect 10152 24818 10180 25298
rect 10244 24818 10272 25366
rect 10140 24812 10192 24818
rect 10140 24754 10192 24760
rect 10232 24812 10284 24818
rect 10232 24754 10284 24760
rect 10048 24608 10100 24614
rect 10048 24550 10100 24556
rect 10060 24410 10088 24550
rect 10048 24404 10100 24410
rect 10048 24346 10100 24352
rect 8944 24200 8996 24206
rect 8944 24142 8996 24148
rect 8956 22098 8984 24142
rect 9312 24132 9364 24138
rect 9312 24074 9364 24080
rect 9324 23866 9352 24074
rect 9390 23964 9698 23973
rect 9390 23962 9396 23964
rect 9452 23962 9476 23964
rect 9532 23962 9556 23964
rect 9612 23962 9636 23964
rect 9692 23962 9698 23964
rect 9452 23910 9454 23962
rect 9634 23910 9636 23962
rect 9390 23908 9396 23910
rect 9452 23908 9476 23910
rect 9532 23908 9556 23910
rect 9612 23908 9636 23910
rect 9692 23908 9698 23910
rect 9390 23899 9698 23908
rect 9312 23860 9364 23866
rect 9312 23802 9364 23808
rect 10152 23662 10180 24754
rect 10140 23656 10192 23662
rect 10140 23598 10192 23604
rect 9390 22876 9698 22885
rect 9390 22874 9396 22876
rect 9452 22874 9476 22876
rect 9532 22874 9556 22876
rect 9612 22874 9636 22876
rect 9692 22874 9698 22876
rect 9452 22822 9454 22874
rect 9634 22822 9636 22874
rect 9390 22820 9396 22822
rect 9452 22820 9476 22822
rect 9532 22820 9556 22822
rect 9612 22820 9636 22822
rect 9692 22820 9698 22822
rect 9390 22811 9698 22820
rect 9036 22704 9088 22710
rect 9036 22646 9088 22652
rect 8944 22092 8996 22098
rect 8944 22034 8996 22040
rect 8484 20936 8536 20942
rect 8484 20878 8536 20884
rect 8496 20602 8524 20878
rect 8484 20596 8536 20602
rect 8484 20538 8536 20544
rect 8956 20466 8984 22034
rect 9048 21350 9076 22646
rect 9864 22636 9916 22642
rect 9916 22596 9996 22624
rect 9864 22578 9916 22584
rect 9864 22432 9916 22438
rect 9864 22374 9916 22380
rect 9312 21956 9364 21962
rect 9312 21898 9364 21904
rect 9324 21690 9352 21898
rect 9390 21788 9698 21797
rect 9390 21786 9396 21788
rect 9452 21786 9476 21788
rect 9532 21786 9556 21788
rect 9612 21786 9636 21788
rect 9692 21786 9698 21788
rect 9452 21734 9454 21786
rect 9634 21734 9636 21786
rect 9390 21732 9396 21734
rect 9452 21732 9476 21734
rect 9532 21732 9556 21734
rect 9612 21732 9636 21734
rect 9692 21732 9698 21734
rect 9390 21723 9698 21732
rect 9312 21684 9364 21690
rect 9312 21626 9364 21632
rect 9876 21554 9904 22374
rect 9864 21548 9916 21554
rect 9864 21490 9916 21496
rect 9968 21350 9996 22596
rect 10232 22432 10284 22438
rect 10232 22374 10284 22380
rect 10244 21622 10272 22374
rect 10232 21616 10284 21622
rect 10232 21558 10284 21564
rect 9036 21344 9088 21350
rect 9036 21286 9088 21292
rect 9220 21344 9272 21350
rect 9220 21286 9272 21292
rect 9956 21344 10008 21350
rect 9956 21286 10008 21292
rect 9232 20602 9260 21286
rect 9772 21140 9824 21146
rect 9772 21082 9824 21088
rect 9312 20800 9364 20806
rect 9312 20742 9364 20748
rect 9220 20596 9272 20602
rect 9220 20538 9272 20544
rect 8944 20460 8996 20466
rect 8944 20402 8996 20408
rect 9232 20262 9260 20538
rect 9324 20534 9352 20742
rect 9390 20700 9698 20709
rect 9390 20698 9396 20700
rect 9452 20698 9476 20700
rect 9532 20698 9556 20700
rect 9612 20698 9636 20700
rect 9692 20698 9698 20700
rect 9452 20646 9454 20698
rect 9634 20646 9636 20698
rect 9390 20644 9396 20646
rect 9452 20644 9476 20646
rect 9532 20644 9556 20646
rect 9612 20644 9636 20646
rect 9692 20644 9698 20646
rect 9390 20635 9698 20644
rect 9312 20528 9364 20534
rect 9312 20470 9364 20476
rect 9312 20392 9364 20398
rect 9312 20334 9364 20340
rect 9220 20256 9272 20262
rect 9220 20198 9272 20204
rect 9324 19922 9352 20334
rect 9312 19916 9364 19922
rect 9312 19858 9364 19864
rect 9784 19854 9812 21082
rect 9968 20466 9996 21286
rect 10428 20942 10456 25842
rect 10600 25764 10652 25770
rect 10600 25706 10652 25712
rect 10612 25294 10640 25706
rect 10600 25288 10652 25294
rect 10600 25230 10652 25236
rect 10612 24954 10640 25230
rect 10968 25220 11020 25226
rect 10968 25162 11020 25168
rect 10600 24948 10652 24954
rect 10600 24890 10652 24896
rect 10980 24818 11008 25162
rect 11060 24948 11112 24954
rect 11060 24890 11112 24896
rect 11072 24818 11100 24890
rect 11164 24818 11192 26930
rect 11612 26784 11664 26790
rect 11612 26726 11664 26732
rect 11624 26586 11652 26726
rect 11612 26580 11664 26586
rect 11612 26522 11664 26528
rect 11992 26382 12020 27066
rect 12164 26988 12216 26994
rect 12164 26930 12216 26936
rect 12072 26852 12124 26858
rect 12072 26794 12124 26800
rect 12084 26450 12112 26794
rect 12176 26450 12204 26930
rect 12072 26444 12124 26450
rect 12072 26386 12124 26392
rect 12164 26444 12216 26450
rect 12164 26386 12216 26392
rect 11336 26376 11388 26382
rect 11336 26318 11388 26324
rect 11980 26376 12032 26382
rect 11980 26318 12032 26324
rect 11244 26240 11296 26246
rect 11244 26182 11296 26188
rect 11256 25906 11284 26182
rect 11244 25900 11296 25906
rect 11244 25842 11296 25848
rect 11348 25702 11376 26318
rect 11612 26240 11664 26246
rect 11612 26182 11664 26188
rect 11796 26240 11848 26246
rect 11796 26182 11848 26188
rect 11624 25906 11652 26182
rect 11612 25900 11664 25906
rect 11612 25842 11664 25848
rect 11336 25696 11388 25702
rect 11336 25638 11388 25644
rect 11244 25356 11296 25362
rect 11244 25298 11296 25304
rect 10508 24812 10560 24818
rect 10508 24754 10560 24760
rect 10600 24812 10652 24818
rect 10600 24754 10652 24760
rect 10968 24812 11020 24818
rect 10968 24754 11020 24760
rect 11060 24812 11112 24818
rect 11060 24754 11112 24760
rect 11152 24812 11204 24818
rect 11152 24754 11204 24760
rect 10520 24342 10548 24754
rect 10508 24336 10560 24342
rect 10508 24278 10560 24284
rect 10612 23322 10640 24754
rect 11256 24750 11284 25298
rect 11348 25294 11376 25638
rect 11336 25288 11388 25294
rect 11336 25230 11388 25236
rect 11428 25288 11480 25294
rect 11428 25230 11480 25236
rect 11244 24744 11296 24750
rect 11440 24698 11468 25230
rect 11520 25152 11572 25158
rect 11520 25094 11572 25100
rect 11244 24686 11296 24692
rect 11348 24670 11468 24698
rect 11348 24614 11376 24670
rect 11336 24608 11388 24614
rect 11164 24556 11336 24562
rect 11164 24550 11388 24556
rect 11164 24534 11376 24550
rect 10692 24336 10744 24342
rect 10692 24278 10744 24284
rect 10600 23316 10652 23322
rect 10600 23258 10652 23264
rect 10612 22094 10640 23258
rect 10704 23118 10732 24278
rect 11164 23866 11192 24534
rect 11244 24064 11296 24070
rect 11244 24006 11296 24012
rect 11256 23866 11284 24006
rect 11532 23866 11560 25094
rect 11152 23860 11204 23866
rect 11152 23802 11204 23808
rect 11244 23860 11296 23866
rect 11244 23802 11296 23808
rect 11520 23860 11572 23866
rect 11520 23802 11572 23808
rect 11520 23724 11572 23730
rect 11520 23666 11572 23672
rect 11244 23656 11296 23662
rect 11244 23598 11296 23604
rect 11060 23520 11112 23526
rect 11060 23462 11112 23468
rect 10692 23112 10744 23118
rect 10692 23054 10744 23060
rect 11072 22658 11100 23462
rect 11256 23322 11284 23598
rect 11244 23316 11296 23322
rect 11244 23258 11296 23264
rect 11256 22778 11284 23258
rect 11244 22772 11296 22778
rect 11244 22714 11296 22720
rect 11072 22630 11284 22658
rect 10784 22568 10836 22574
rect 10784 22510 10836 22516
rect 10796 22166 10824 22510
rect 11152 22432 11204 22438
rect 11152 22374 11204 22380
rect 10784 22160 10836 22166
rect 10784 22102 10836 22108
rect 10612 22066 10732 22094
rect 10704 21554 10732 22066
rect 10796 21554 10824 22102
rect 11164 22030 11192 22374
rect 11256 22030 11284 22630
rect 11532 22574 11560 23666
rect 11520 22568 11572 22574
rect 11520 22510 11572 22516
rect 11624 22094 11652 25842
rect 11704 24608 11756 24614
rect 11704 24550 11756 24556
rect 11716 23866 11744 24550
rect 11704 23860 11756 23866
rect 11704 23802 11756 23808
rect 11808 23644 11836 26182
rect 12084 25702 12112 26386
rect 11980 25696 12032 25702
rect 11980 25638 12032 25644
rect 12072 25696 12124 25702
rect 12072 25638 12124 25644
rect 11992 25362 12020 25638
rect 12084 25498 12112 25638
rect 12072 25492 12124 25498
rect 12072 25434 12124 25440
rect 12268 25378 12296 27406
rect 12452 27130 12480 27474
rect 12532 27464 12584 27470
rect 12532 27406 12584 27412
rect 12900 27464 12952 27470
rect 12900 27406 12952 27412
rect 12544 27130 12572 27406
rect 12624 27328 12676 27334
rect 12624 27270 12676 27276
rect 12440 27124 12492 27130
rect 12440 27066 12492 27072
rect 12532 27124 12584 27130
rect 12532 27066 12584 27072
rect 12348 26376 12400 26382
rect 12348 26318 12400 26324
rect 12360 25974 12388 26318
rect 12544 26194 12572 27066
rect 12636 26790 12664 27270
rect 12808 27056 12860 27062
rect 12808 26998 12860 27004
rect 12820 26790 12848 26998
rect 12624 26784 12676 26790
rect 12624 26726 12676 26732
rect 12808 26784 12860 26790
rect 12808 26726 12860 26732
rect 12636 26450 12664 26726
rect 12624 26444 12676 26450
rect 12624 26386 12676 26392
rect 12544 26166 12664 26194
rect 12348 25968 12400 25974
rect 12348 25910 12400 25916
rect 12636 25906 12664 26166
rect 12440 25900 12492 25906
rect 12440 25842 12492 25848
rect 12624 25900 12676 25906
rect 12624 25842 12676 25848
rect 12716 25900 12768 25906
rect 12716 25842 12768 25848
rect 12452 25378 12480 25842
rect 11888 25356 11940 25362
rect 11888 25298 11940 25304
rect 11980 25356 12032 25362
rect 11980 25298 12032 25304
rect 12268 25350 12480 25378
rect 11900 24614 11928 25298
rect 12268 25294 12296 25350
rect 12636 25294 12664 25842
rect 12728 25498 12756 25842
rect 12716 25492 12768 25498
rect 12716 25434 12768 25440
rect 12164 25288 12216 25294
rect 12164 25230 12216 25236
rect 12256 25288 12308 25294
rect 12256 25230 12308 25236
rect 12624 25288 12676 25294
rect 12624 25230 12676 25236
rect 11980 25220 12032 25226
rect 11980 25162 12032 25168
rect 11992 24954 12020 25162
rect 12176 24954 12204 25230
rect 12268 24954 12296 25230
rect 11980 24948 12032 24954
rect 11980 24890 12032 24896
rect 12164 24948 12216 24954
rect 12164 24890 12216 24896
rect 12256 24948 12308 24954
rect 12256 24890 12308 24896
rect 12532 24744 12584 24750
rect 12532 24686 12584 24692
rect 11888 24608 11940 24614
rect 11888 24550 11940 24556
rect 12544 24410 12572 24686
rect 12532 24404 12584 24410
rect 12532 24346 12584 24352
rect 12716 24200 12768 24206
rect 12716 24142 12768 24148
rect 12164 24064 12216 24070
rect 12164 24006 12216 24012
rect 11888 23656 11940 23662
rect 11808 23616 11888 23644
rect 11888 23598 11940 23604
rect 11900 23526 11928 23598
rect 11888 23520 11940 23526
rect 11888 23462 11940 23468
rect 12176 23118 12204 24006
rect 12728 23866 12756 24142
rect 12716 23860 12768 23866
rect 12716 23802 12768 23808
rect 12164 23112 12216 23118
rect 12164 23054 12216 23060
rect 12532 23112 12584 23118
rect 12532 23054 12584 23060
rect 12440 22432 12492 22438
rect 12440 22374 12492 22380
rect 12452 22166 12480 22374
rect 12440 22160 12492 22166
rect 12440 22102 12492 22108
rect 11532 22066 11652 22094
rect 11980 22092 12032 22098
rect 11532 22030 11560 22066
rect 11980 22034 12032 22040
rect 10968 22024 11020 22030
rect 10968 21966 11020 21972
rect 11152 22024 11204 22030
rect 11152 21966 11204 21972
rect 11244 22024 11296 22030
rect 11244 21966 11296 21972
rect 11520 22024 11572 22030
rect 11520 21966 11572 21972
rect 10980 21690 11008 21966
rect 11164 21690 11192 21966
rect 11888 21888 11940 21894
rect 11888 21830 11940 21836
rect 11900 21690 11928 21830
rect 10968 21684 11020 21690
rect 10968 21626 11020 21632
rect 11152 21684 11204 21690
rect 11152 21626 11204 21632
rect 11888 21684 11940 21690
rect 11888 21626 11940 21632
rect 10692 21548 10744 21554
rect 10692 21490 10744 21496
rect 10784 21548 10836 21554
rect 10784 21490 10836 21496
rect 10968 21548 11020 21554
rect 10968 21490 11020 21496
rect 11888 21548 11940 21554
rect 11992 21536 12020 22034
rect 12072 22024 12124 22030
rect 12072 21966 12124 21972
rect 12084 21554 12112 21966
rect 12348 21888 12400 21894
rect 12348 21830 12400 21836
rect 11940 21508 12020 21536
rect 12072 21548 12124 21554
rect 11888 21490 11940 21496
rect 12072 21490 12124 21496
rect 10980 21010 11008 21490
rect 10968 21004 11020 21010
rect 10968 20946 11020 20952
rect 10416 20936 10468 20942
rect 10416 20878 10468 20884
rect 10980 20602 11008 20946
rect 11060 20800 11112 20806
rect 11060 20742 11112 20748
rect 11704 20800 11756 20806
rect 11704 20742 11756 20748
rect 11072 20602 11100 20742
rect 10968 20596 11020 20602
rect 10968 20538 11020 20544
rect 11060 20596 11112 20602
rect 11060 20538 11112 20544
rect 9956 20460 10008 20466
rect 9956 20402 10008 20408
rect 10048 20460 10100 20466
rect 10048 20402 10100 20408
rect 9772 19848 9824 19854
rect 9772 19790 9824 19796
rect 9968 19786 9996 20402
rect 10060 20058 10088 20402
rect 11060 20256 11112 20262
rect 11060 20198 11112 20204
rect 10048 20052 10100 20058
rect 10048 19994 10100 20000
rect 10692 19848 10744 19854
rect 10692 19790 10744 19796
rect 9956 19780 10008 19786
rect 9956 19722 10008 19728
rect 10600 19780 10652 19786
rect 10600 19722 10652 19728
rect 7656 19712 7708 19718
rect 7656 19654 7708 19660
rect 9390 19612 9698 19621
rect 9390 19610 9396 19612
rect 9452 19610 9476 19612
rect 9532 19610 9556 19612
rect 9612 19610 9636 19612
rect 9692 19610 9698 19612
rect 9452 19558 9454 19610
rect 9634 19558 9636 19610
rect 9390 19556 9396 19558
rect 9452 19556 9476 19558
rect 9532 19556 9556 19558
rect 9612 19556 9636 19558
rect 9692 19556 9698 19558
rect 9390 19547 9698 19556
rect 10612 19514 10640 19722
rect 10704 19514 10732 19790
rect 10600 19508 10652 19514
rect 10600 19450 10652 19456
rect 10692 19508 10744 19514
rect 10692 19450 10744 19456
rect 11072 19378 11100 20198
rect 11716 20058 11744 20742
rect 11704 20052 11756 20058
rect 11704 19994 11756 20000
rect 11900 19990 11928 21490
rect 12360 20806 12388 21830
rect 12452 21554 12480 22102
rect 12440 21548 12492 21554
rect 12440 21490 12492 21496
rect 12544 20874 12572 23054
rect 12820 22642 12848 26726
rect 12912 26586 12940 27406
rect 12992 26784 13044 26790
rect 12992 26726 13044 26732
rect 12900 26580 12952 26586
rect 12900 26522 12952 26528
rect 13004 26382 13032 26726
rect 12992 26376 13044 26382
rect 12992 26318 13044 26324
rect 13004 25906 13032 26318
rect 12992 25900 13044 25906
rect 12912 25860 12992 25888
rect 12912 25362 12940 25860
rect 12992 25842 13044 25848
rect 12900 25356 12952 25362
rect 12900 25298 12952 25304
rect 12992 24812 13044 24818
rect 12992 24754 13044 24760
rect 13004 24206 13032 24754
rect 12992 24200 13044 24206
rect 12992 24142 13044 24148
rect 12900 24064 12952 24070
rect 12900 24006 12952 24012
rect 12912 23050 12940 24006
rect 13004 23730 13032 24142
rect 12992 23724 13044 23730
rect 12992 23666 13044 23672
rect 12900 23044 12952 23050
rect 12900 22986 12952 22992
rect 13096 22642 13124 27474
rect 13360 26988 13412 26994
rect 13360 26930 13412 26936
rect 13268 25968 13320 25974
rect 13268 25910 13320 25916
rect 13176 25900 13228 25906
rect 13176 25842 13228 25848
rect 13188 25702 13216 25842
rect 13176 25696 13228 25702
rect 13176 25638 13228 25644
rect 13188 25294 13216 25638
rect 13280 25378 13308 25910
rect 13372 25498 13400 26930
rect 13464 26466 13492 27814
rect 13611 27772 13919 27781
rect 13611 27770 13617 27772
rect 13673 27770 13697 27772
rect 13753 27770 13777 27772
rect 13833 27770 13857 27772
rect 13913 27770 13919 27772
rect 13673 27718 13675 27770
rect 13855 27718 13857 27770
rect 13611 27716 13617 27718
rect 13673 27716 13697 27718
rect 13753 27716 13777 27718
rect 13833 27716 13857 27718
rect 13913 27716 13919 27718
rect 13611 27707 13919 27716
rect 13544 27328 13596 27334
rect 13544 27270 13596 27276
rect 13912 27328 13964 27334
rect 13912 27270 13964 27276
rect 13556 27130 13584 27270
rect 13924 27130 13952 27270
rect 13544 27124 13596 27130
rect 13544 27066 13596 27072
rect 13912 27124 13964 27130
rect 13912 27066 13964 27072
rect 14016 26994 14044 27900
rect 14108 27470 14136 28970
rect 14384 28762 14412 29106
rect 14752 29034 14780 29174
rect 14740 29028 14792 29034
rect 14740 28970 14792 28976
rect 14372 28756 14424 28762
rect 14372 28698 14424 28704
rect 14280 28416 14332 28422
rect 14280 28358 14332 28364
rect 14188 28076 14240 28082
rect 14188 28018 14240 28024
rect 14200 27674 14228 28018
rect 14188 27668 14240 27674
rect 14188 27610 14240 27616
rect 14096 27464 14148 27470
rect 14096 27406 14148 27412
rect 14004 26988 14056 26994
rect 14004 26930 14056 26936
rect 13611 26684 13919 26693
rect 13611 26682 13617 26684
rect 13673 26682 13697 26684
rect 13753 26682 13777 26684
rect 13833 26682 13857 26684
rect 13913 26682 13919 26684
rect 13673 26630 13675 26682
rect 13855 26630 13857 26682
rect 13611 26628 13617 26630
rect 13673 26628 13697 26630
rect 13753 26628 13777 26630
rect 13833 26628 13857 26630
rect 13913 26628 13919 26630
rect 13611 26619 13919 26628
rect 13464 26438 13584 26466
rect 13452 26376 13504 26382
rect 13452 26318 13504 26324
rect 13464 25498 13492 26318
rect 13556 25906 13584 26438
rect 14292 26382 14320 28358
rect 15028 27452 15056 30806
rect 15108 30728 15160 30734
rect 15108 30670 15160 30676
rect 15120 30394 15148 30670
rect 15108 30388 15160 30394
rect 15108 30330 15160 30336
rect 15212 28490 15240 34575
rect 15396 34406 15424 37062
rect 15936 36712 15988 36718
rect 15936 36654 15988 36660
rect 15948 36378 15976 36654
rect 15936 36372 15988 36378
rect 15936 36314 15988 36320
rect 15476 36304 15528 36310
rect 15476 36246 15528 36252
rect 15488 36145 15516 36246
rect 15474 36136 15530 36145
rect 15474 36071 15530 36080
rect 16212 36032 16264 36038
rect 16212 35974 16264 35980
rect 16028 35692 16080 35698
rect 16028 35634 16080 35640
rect 16040 34746 16068 35634
rect 16120 35488 16172 35494
rect 16120 35430 16172 35436
rect 16132 35290 16160 35430
rect 16120 35284 16172 35290
rect 16120 35226 16172 35232
rect 16132 34746 16160 35226
rect 16224 34746 16252 35974
rect 16316 35562 16344 37062
rect 16960 36242 16988 37062
rect 17052 36854 17080 37062
rect 17040 36848 17092 36854
rect 17040 36790 17092 36796
rect 16764 36236 16816 36242
rect 16764 36178 16816 36184
rect 16948 36236 17000 36242
rect 16948 36178 17000 36184
rect 16488 36032 16540 36038
rect 16488 35974 16540 35980
rect 16672 36032 16724 36038
rect 16672 35974 16724 35980
rect 16304 35556 16356 35562
rect 16304 35498 16356 35504
rect 16316 35170 16344 35498
rect 16316 35142 16436 35170
rect 16304 35080 16356 35086
rect 16304 35022 16356 35028
rect 16316 34746 16344 35022
rect 16028 34740 16080 34746
rect 16028 34682 16080 34688
rect 16120 34740 16172 34746
rect 16120 34682 16172 34688
rect 16212 34740 16264 34746
rect 16212 34682 16264 34688
rect 16304 34740 16356 34746
rect 16304 34682 16356 34688
rect 15658 34640 15714 34649
rect 16408 34610 16436 35142
rect 16500 34649 16528 35974
rect 16684 35834 16712 35974
rect 16672 35828 16724 35834
rect 16672 35770 16724 35776
rect 16776 35766 16804 36178
rect 17236 36174 17264 37606
rect 17328 37466 17356 39238
rect 17408 37800 17460 37806
rect 17408 37742 17460 37748
rect 17316 37460 17368 37466
rect 17316 37402 17368 37408
rect 17420 37346 17448 37742
rect 17512 37738 17540 39374
rect 17604 38350 17632 39374
rect 17831 39196 18139 39205
rect 17831 39194 17837 39196
rect 17893 39194 17917 39196
rect 17973 39194 17997 39196
rect 18053 39194 18077 39196
rect 18133 39194 18139 39196
rect 17893 39142 17895 39194
rect 18075 39142 18077 39194
rect 17831 39140 17837 39142
rect 17893 39140 17917 39142
rect 17973 39140 17997 39142
rect 18053 39140 18077 39142
rect 18133 39140 18139 39142
rect 17831 39131 18139 39140
rect 18248 38554 18276 39374
rect 18236 38548 18288 38554
rect 18236 38490 18288 38496
rect 17592 38344 17644 38350
rect 17592 38286 17644 38292
rect 18236 38344 18288 38350
rect 18236 38286 18288 38292
rect 17831 38108 18139 38117
rect 17831 38106 17837 38108
rect 17893 38106 17917 38108
rect 17973 38106 17997 38108
rect 18053 38106 18077 38108
rect 18133 38106 18139 38108
rect 17893 38054 17895 38106
rect 18075 38054 18077 38106
rect 17831 38052 17837 38054
rect 17893 38052 17917 38054
rect 17973 38052 17997 38054
rect 18053 38052 18077 38054
rect 18133 38052 18139 38054
rect 17831 38043 18139 38052
rect 17684 38004 17736 38010
rect 17684 37946 17736 37952
rect 17592 37868 17644 37874
rect 17592 37810 17644 37816
rect 17500 37732 17552 37738
rect 17500 37674 17552 37680
rect 17328 37318 17448 37346
rect 17328 37262 17356 37318
rect 17604 37262 17632 37810
rect 17696 37466 17724 37946
rect 18052 37936 18104 37942
rect 18052 37878 18104 37884
rect 17868 37800 17920 37806
rect 17868 37742 17920 37748
rect 17776 37732 17828 37738
rect 17776 37674 17828 37680
rect 17684 37460 17736 37466
rect 17684 37402 17736 37408
rect 17788 37398 17816 37674
rect 17880 37466 17908 37742
rect 17868 37460 17920 37466
rect 17868 37402 17920 37408
rect 17776 37392 17828 37398
rect 17776 37334 17828 37340
rect 18064 37330 18092 37878
rect 18144 37664 18196 37670
rect 18144 37606 18196 37612
rect 18052 37324 18104 37330
rect 18052 37266 18104 37272
rect 18156 37262 18184 37606
rect 17316 37256 17368 37262
rect 17316 37198 17368 37204
rect 17592 37256 17644 37262
rect 17592 37198 17644 37204
rect 18144 37256 18196 37262
rect 18144 37198 18196 37204
rect 17328 36922 17356 37198
rect 18248 37194 18276 38286
rect 18236 37188 18288 37194
rect 18236 37130 18288 37136
rect 18340 37126 18368 39578
rect 21928 39506 21956 41200
rect 22052 39740 22360 39749
rect 22052 39738 22058 39740
rect 22114 39738 22138 39740
rect 22194 39738 22218 39740
rect 22274 39738 22298 39740
rect 22354 39738 22360 39740
rect 22114 39686 22116 39738
rect 22296 39686 22298 39738
rect 22052 39684 22058 39686
rect 22114 39684 22138 39686
rect 22194 39684 22218 39686
rect 22274 39684 22298 39686
rect 22354 39684 22360 39686
rect 22052 39675 22360 39684
rect 22836 39568 22888 39574
rect 22836 39510 22888 39516
rect 21916 39500 21968 39506
rect 21916 39442 21968 39448
rect 19156 39364 19208 39370
rect 19156 39306 19208 39312
rect 22744 39364 22796 39370
rect 22744 39306 22796 39312
rect 18512 38752 18564 38758
rect 18512 38694 18564 38700
rect 18524 38418 18552 38694
rect 18512 38412 18564 38418
rect 18512 38354 18564 38360
rect 18420 38208 18472 38214
rect 18420 38150 18472 38156
rect 17684 37120 17736 37126
rect 17684 37062 17736 37068
rect 18328 37120 18380 37126
rect 18328 37062 18380 37068
rect 17316 36916 17368 36922
rect 17316 36858 17368 36864
rect 17696 36854 17724 37062
rect 17831 37020 18139 37029
rect 17831 37018 17837 37020
rect 17893 37018 17917 37020
rect 17973 37018 17997 37020
rect 18053 37018 18077 37020
rect 18133 37018 18139 37020
rect 17893 36966 17895 37018
rect 18075 36966 18077 37018
rect 17831 36964 17837 36966
rect 17893 36964 17917 36966
rect 17973 36964 17997 36966
rect 18053 36964 18077 36966
rect 18133 36964 18139 36966
rect 17831 36955 18139 36964
rect 17684 36848 17736 36854
rect 17684 36790 17736 36796
rect 17316 36304 17368 36310
rect 17316 36246 17368 36252
rect 17224 36168 17276 36174
rect 17224 36110 17276 36116
rect 17328 35766 17356 36246
rect 17500 36168 17552 36174
rect 17500 36110 17552 36116
rect 16764 35760 16816 35766
rect 16764 35702 16816 35708
rect 17316 35760 17368 35766
rect 17316 35702 17368 35708
rect 17224 35488 17276 35494
rect 17224 35430 17276 35436
rect 17236 35290 17264 35430
rect 17224 35284 17276 35290
rect 17224 35226 17276 35232
rect 17224 35148 17276 35154
rect 17224 35090 17276 35096
rect 16856 34944 16908 34950
rect 16856 34886 16908 34892
rect 16868 34746 16896 34886
rect 17236 34746 17264 35090
rect 16856 34740 16908 34746
rect 16856 34682 16908 34688
rect 17224 34740 17276 34746
rect 17224 34682 17276 34688
rect 16486 34640 16542 34649
rect 15658 34575 15660 34584
rect 15712 34575 15714 34584
rect 16396 34604 16448 34610
rect 15660 34546 15712 34552
rect 16486 34575 16542 34584
rect 16396 34546 16448 34552
rect 15844 34536 15896 34542
rect 15844 34478 15896 34484
rect 15292 34400 15344 34406
rect 15292 34342 15344 34348
rect 15384 34400 15436 34406
rect 15384 34342 15436 34348
rect 15304 33998 15332 34342
rect 15292 33992 15344 33998
rect 15292 33934 15344 33940
rect 15292 32360 15344 32366
rect 15290 32328 15292 32337
rect 15344 32328 15346 32337
rect 15396 32314 15424 34342
rect 15856 33658 15884 34478
rect 17328 34474 17356 35702
rect 17408 35284 17460 35290
rect 17408 35226 17460 35232
rect 17316 34468 17368 34474
rect 17316 34410 17368 34416
rect 15936 33856 15988 33862
rect 15936 33798 15988 33804
rect 16948 33856 17000 33862
rect 16948 33798 17000 33804
rect 15844 33652 15896 33658
rect 15844 33594 15896 33600
rect 15476 33516 15528 33522
rect 15476 33458 15528 33464
rect 15488 33046 15516 33458
rect 15752 33448 15804 33454
rect 15752 33390 15804 33396
rect 15660 33380 15712 33386
rect 15660 33322 15712 33328
rect 15568 33312 15620 33318
rect 15568 33254 15620 33260
rect 15476 33040 15528 33046
rect 15476 32982 15528 32988
rect 15476 32836 15528 32842
rect 15476 32778 15528 32784
rect 15488 32570 15516 32778
rect 15476 32564 15528 32570
rect 15476 32506 15528 32512
rect 15580 32434 15608 33254
rect 15672 32978 15700 33322
rect 15764 32978 15792 33390
rect 15660 32972 15712 32978
rect 15660 32914 15712 32920
rect 15752 32972 15804 32978
rect 15752 32914 15804 32920
rect 15672 32570 15700 32914
rect 15660 32564 15712 32570
rect 15660 32506 15712 32512
rect 15764 32434 15792 32914
rect 15568 32428 15620 32434
rect 15568 32370 15620 32376
rect 15752 32428 15804 32434
rect 15752 32370 15804 32376
rect 15844 32360 15896 32366
rect 15396 32286 15792 32314
rect 15844 32302 15896 32308
rect 15290 32263 15346 32272
rect 15660 32224 15712 32230
rect 15660 32166 15712 32172
rect 15672 31754 15700 32166
rect 15580 31726 15700 31754
rect 15476 31680 15528 31686
rect 15476 31622 15528 31628
rect 15384 30728 15436 30734
rect 15384 30670 15436 30676
rect 15292 30592 15344 30598
rect 15292 30534 15344 30540
rect 15304 29646 15332 30534
rect 15396 29850 15424 30670
rect 15488 30258 15516 31622
rect 15580 31210 15608 31726
rect 15568 31204 15620 31210
rect 15568 31146 15620 31152
rect 15660 31136 15712 31142
rect 15660 31078 15712 31084
rect 15476 30252 15528 30258
rect 15476 30194 15528 30200
rect 15568 30252 15620 30258
rect 15568 30194 15620 30200
rect 15580 29850 15608 30194
rect 15384 29844 15436 29850
rect 15384 29786 15436 29792
rect 15568 29844 15620 29850
rect 15568 29786 15620 29792
rect 15476 29708 15528 29714
rect 15476 29650 15528 29656
rect 15292 29640 15344 29646
rect 15292 29582 15344 29588
rect 15200 28484 15252 28490
rect 15200 28426 15252 28432
rect 15384 28484 15436 28490
rect 15384 28426 15436 28432
rect 15396 28218 15424 28426
rect 15384 28212 15436 28218
rect 15384 28154 15436 28160
rect 15292 27872 15344 27878
rect 15292 27814 15344 27820
rect 15304 27470 15332 27814
rect 14936 27424 15056 27452
rect 15292 27464 15344 27470
rect 14280 26376 14332 26382
rect 14280 26318 14332 26324
rect 14648 26376 14700 26382
rect 14648 26318 14700 26324
rect 13544 25900 13596 25906
rect 13544 25842 13596 25848
rect 14188 25900 14240 25906
rect 14188 25842 14240 25848
rect 13611 25596 13919 25605
rect 13611 25594 13617 25596
rect 13673 25594 13697 25596
rect 13753 25594 13777 25596
rect 13833 25594 13857 25596
rect 13913 25594 13919 25596
rect 13673 25542 13675 25594
rect 13855 25542 13857 25594
rect 13611 25540 13617 25542
rect 13673 25540 13697 25542
rect 13753 25540 13777 25542
rect 13833 25540 13857 25542
rect 13913 25540 13919 25542
rect 13611 25531 13919 25540
rect 13360 25492 13412 25498
rect 13360 25434 13412 25440
rect 13452 25492 13504 25498
rect 13452 25434 13504 25440
rect 13728 25492 13780 25498
rect 13728 25434 13780 25440
rect 13280 25350 13400 25378
rect 13176 25288 13228 25294
rect 13176 25230 13228 25236
rect 13188 24750 13216 25230
rect 13372 25158 13400 25350
rect 13360 25152 13412 25158
rect 13360 25094 13412 25100
rect 13372 24818 13400 25094
rect 13740 24818 13768 25434
rect 14200 25226 14228 25842
rect 14556 25696 14608 25702
rect 14556 25638 14608 25644
rect 14568 25430 14596 25638
rect 14556 25424 14608 25430
rect 14556 25366 14608 25372
rect 14188 25220 14240 25226
rect 14464 25220 14516 25226
rect 14240 25180 14320 25208
rect 14188 25162 14240 25168
rect 13360 24812 13412 24818
rect 13360 24754 13412 24760
rect 13728 24812 13780 24818
rect 13728 24754 13780 24760
rect 14004 24812 14056 24818
rect 14004 24754 14056 24760
rect 14188 24812 14240 24818
rect 14188 24754 14240 24760
rect 13176 24744 13228 24750
rect 13176 24686 13228 24692
rect 13188 24410 13216 24686
rect 13176 24404 13228 24410
rect 13176 24346 13228 24352
rect 13372 24070 13400 24754
rect 13611 24508 13919 24517
rect 13611 24506 13617 24508
rect 13673 24506 13697 24508
rect 13753 24506 13777 24508
rect 13833 24506 13857 24508
rect 13913 24506 13919 24508
rect 13673 24454 13675 24506
rect 13855 24454 13857 24506
rect 13611 24452 13617 24454
rect 13673 24452 13697 24454
rect 13753 24452 13777 24454
rect 13833 24452 13857 24454
rect 13913 24452 13919 24454
rect 13611 24443 13919 24452
rect 14016 24410 14044 24754
rect 14096 24676 14148 24682
rect 14096 24618 14148 24624
rect 14108 24410 14136 24618
rect 14004 24404 14056 24410
rect 14004 24346 14056 24352
rect 14096 24404 14148 24410
rect 14096 24346 14148 24352
rect 14200 24290 14228 24754
rect 14292 24682 14320 25180
rect 14464 25162 14516 25168
rect 14372 25152 14424 25158
rect 14372 25094 14424 25100
rect 14280 24676 14332 24682
rect 14280 24618 14332 24624
rect 14016 24274 14228 24290
rect 14384 24274 14412 25094
rect 14476 24886 14504 25162
rect 14464 24880 14516 24886
rect 14464 24822 14516 24828
rect 14556 24812 14608 24818
rect 14556 24754 14608 24760
rect 14568 24342 14596 24754
rect 14556 24336 14608 24342
rect 14556 24278 14608 24284
rect 14004 24268 14228 24274
rect 14056 24262 14228 24268
rect 14372 24268 14424 24274
rect 14004 24210 14056 24216
rect 14372 24210 14424 24216
rect 13452 24200 13504 24206
rect 13452 24142 13504 24148
rect 14280 24200 14332 24206
rect 14280 24142 14332 24148
rect 13360 24064 13412 24070
rect 13360 24006 13412 24012
rect 13464 23866 13492 24142
rect 13728 24132 13780 24138
rect 13728 24074 13780 24080
rect 13740 23866 13768 24074
rect 14292 23866 14320 24142
rect 13452 23860 13504 23866
rect 13452 23802 13504 23808
rect 13728 23860 13780 23866
rect 13728 23802 13780 23808
rect 14280 23860 14332 23866
rect 14280 23802 14332 23808
rect 13726 23760 13782 23769
rect 13176 23724 13228 23730
rect 14384 23730 14412 24210
rect 14464 24132 14516 24138
rect 14464 24074 14516 24080
rect 14476 23866 14504 24074
rect 14464 23860 14516 23866
rect 14464 23802 14516 23808
rect 13726 23695 13728 23704
rect 13176 23666 13228 23672
rect 13780 23695 13782 23704
rect 14188 23724 14240 23730
rect 13728 23666 13780 23672
rect 14188 23666 14240 23672
rect 14372 23724 14424 23730
rect 14372 23666 14424 23672
rect 13188 23526 13216 23666
rect 13176 23520 13228 23526
rect 13176 23462 13228 23468
rect 13611 23420 13919 23429
rect 13611 23418 13617 23420
rect 13673 23418 13697 23420
rect 13753 23418 13777 23420
rect 13833 23418 13857 23420
rect 13913 23418 13919 23420
rect 13673 23366 13675 23418
rect 13855 23366 13857 23418
rect 13611 23364 13617 23366
rect 13673 23364 13697 23366
rect 13753 23364 13777 23366
rect 13833 23364 13857 23366
rect 13913 23364 13919 23366
rect 13611 23355 13919 23364
rect 14200 23322 14228 23666
rect 14464 23520 14516 23526
rect 14464 23462 14516 23468
rect 14476 23322 14504 23462
rect 14188 23316 14240 23322
rect 14188 23258 14240 23264
rect 14464 23316 14516 23322
rect 14464 23258 14516 23264
rect 14096 23248 14148 23254
rect 14096 23190 14148 23196
rect 13544 23112 13596 23118
rect 13544 23054 13596 23060
rect 13452 22704 13504 22710
rect 13452 22646 13504 22652
rect 12808 22636 12860 22642
rect 12808 22578 12860 22584
rect 13084 22636 13136 22642
rect 13084 22578 13136 22584
rect 13096 22234 13124 22578
rect 13176 22500 13228 22506
rect 13176 22442 13228 22448
rect 13084 22228 13136 22234
rect 13084 22170 13136 22176
rect 12624 22024 12676 22030
rect 12624 21966 12676 21972
rect 12636 21690 12664 21966
rect 12716 21888 12768 21894
rect 12716 21830 12768 21836
rect 12992 21888 13044 21894
rect 12992 21830 13044 21836
rect 12624 21684 12676 21690
rect 12624 21626 12676 21632
rect 12624 21548 12676 21554
rect 12728 21536 12756 21830
rect 13004 21690 13032 21830
rect 12992 21684 13044 21690
rect 12992 21626 13044 21632
rect 13188 21536 13216 22442
rect 13268 22432 13320 22438
rect 13268 22374 13320 22380
rect 13360 22432 13412 22438
rect 13360 22374 13412 22380
rect 13280 22098 13308 22374
rect 13268 22092 13320 22098
rect 13268 22034 13320 22040
rect 13268 21548 13320 21554
rect 12676 21508 12756 21536
rect 13004 21508 13268 21536
rect 12624 21490 12676 21496
rect 12636 20924 12664 21490
rect 12808 20936 12860 20942
rect 12636 20896 12808 20924
rect 12808 20878 12860 20884
rect 12532 20868 12584 20874
rect 12532 20810 12584 20816
rect 12256 20800 12308 20806
rect 12256 20742 12308 20748
rect 12348 20800 12400 20806
rect 12348 20742 12400 20748
rect 12268 20466 12296 20742
rect 12348 20528 12400 20534
rect 12348 20470 12400 20476
rect 12256 20460 12308 20466
rect 12256 20402 12308 20408
rect 11888 19984 11940 19990
rect 11888 19926 11940 19932
rect 11900 19378 11928 19926
rect 12360 19378 12388 20470
rect 12544 20466 12572 20810
rect 12532 20460 12584 20466
rect 12532 20402 12584 20408
rect 12440 20256 12492 20262
rect 12440 20198 12492 20204
rect 12716 20256 12768 20262
rect 12716 20198 12768 20204
rect 12452 19514 12480 20198
rect 12728 19854 12756 20198
rect 12716 19848 12768 19854
rect 12716 19790 12768 19796
rect 12820 19718 12848 20878
rect 13004 20806 13032 21508
rect 13268 21490 13320 21496
rect 13372 21434 13400 22374
rect 13464 21486 13492 22646
rect 13556 22574 13584 23054
rect 14108 22642 14136 23190
rect 14200 22778 14228 23258
rect 14568 22778 14596 24278
rect 14660 23866 14688 26318
rect 14832 26308 14884 26314
rect 14936 26296 14964 27424
rect 15292 27406 15344 27412
rect 15488 27062 15516 29650
rect 15672 29646 15700 31078
rect 15764 30938 15792 32286
rect 15856 32026 15884 32302
rect 15844 32020 15896 32026
rect 15844 31962 15896 31968
rect 15948 31906 15976 33798
rect 16960 33522 16988 33798
rect 16120 33516 16172 33522
rect 16120 33458 16172 33464
rect 16580 33516 16632 33522
rect 16580 33458 16632 33464
rect 16856 33516 16908 33522
rect 16856 33458 16908 33464
rect 16948 33516 17000 33522
rect 16948 33458 17000 33464
rect 17132 33516 17184 33522
rect 17132 33458 17184 33464
rect 16132 33114 16160 33458
rect 16212 33448 16264 33454
rect 16212 33390 16264 33396
rect 16120 33108 16172 33114
rect 16120 33050 16172 33056
rect 16224 32910 16252 33390
rect 16304 33312 16356 33318
rect 16304 33254 16356 33260
rect 16212 32904 16264 32910
rect 16212 32846 16264 32852
rect 16212 32768 16264 32774
rect 16212 32710 16264 32716
rect 15856 31878 15976 31906
rect 16224 31890 16252 32710
rect 16316 32434 16344 33254
rect 16592 32881 16620 33458
rect 16868 33114 16896 33458
rect 16856 33108 16908 33114
rect 16856 33050 16908 33056
rect 16578 32872 16634 32881
rect 17144 32842 17172 33458
rect 17316 33380 17368 33386
rect 17316 33322 17368 33328
rect 16578 32807 16634 32816
rect 17132 32836 17184 32842
rect 16592 32570 16620 32807
rect 17132 32778 17184 32784
rect 16580 32564 16632 32570
rect 16580 32506 16632 32512
rect 17144 32434 17172 32778
rect 17328 32434 17356 33322
rect 17420 33046 17448 35226
rect 17512 34134 17540 36110
rect 17696 35698 17724 36790
rect 17868 36236 17920 36242
rect 17868 36178 17920 36184
rect 17880 36106 17908 36178
rect 17868 36100 17920 36106
rect 17868 36042 17920 36048
rect 18432 36038 18460 38150
rect 18524 37874 18552 38354
rect 19168 37942 19196 39306
rect 20536 39296 20588 39302
rect 20536 39238 20588 39244
rect 21456 39296 21508 39302
rect 21456 39238 21508 39244
rect 20548 39098 20576 39238
rect 21468 39098 21496 39238
rect 20536 39092 20588 39098
rect 20536 39034 20588 39040
rect 21456 39092 21508 39098
rect 21456 39034 21508 39040
rect 21640 39092 21692 39098
rect 21640 39034 21692 39040
rect 19340 38888 19392 38894
rect 19340 38830 19392 38836
rect 19352 38350 19380 38830
rect 21272 38412 21324 38418
rect 21272 38354 21324 38360
rect 19340 38344 19392 38350
rect 19340 38286 19392 38292
rect 19156 37936 19208 37942
rect 19156 37878 19208 37884
rect 19248 37936 19300 37942
rect 19248 37878 19300 37884
rect 18512 37868 18564 37874
rect 18512 37810 18564 37816
rect 18604 37868 18656 37874
rect 18604 37810 18656 37816
rect 18616 36786 18644 37810
rect 19064 37188 19116 37194
rect 19064 37130 19116 37136
rect 18604 36780 18656 36786
rect 18604 36722 18656 36728
rect 19076 36378 19104 37130
rect 19064 36372 19116 36378
rect 19064 36314 19116 36320
rect 19168 36242 19196 37878
rect 19260 37466 19288 37878
rect 19352 37806 19380 38286
rect 20720 38276 20772 38282
rect 20720 38218 20772 38224
rect 20732 38010 20760 38218
rect 21284 38010 21312 38354
rect 20720 38004 20772 38010
rect 20720 37946 20772 37952
rect 21272 38004 21324 38010
rect 21272 37946 21324 37952
rect 21548 38004 21600 38010
rect 21548 37946 21600 37952
rect 21560 37874 21588 37946
rect 21652 37874 21680 39034
rect 21824 38752 21876 38758
rect 21824 38694 21876 38700
rect 21836 38418 21864 38694
rect 22052 38652 22360 38661
rect 22052 38650 22058 38652
rect 22114 38650 22138 38652
rect 22194 38650 22218 38652
rect 22274 38650 22298 38652
rect 22354 38650 22360 38652
rect 22114 38598 22116 38650
rect 22296 38598 22298 38650
rect 22052 38596 22058 38598
rect 22114 38596 22138 38598
rect 22194 38596 22218 38598
rect 22274 38596 22298 38598
rect 22354 38596 22360 38598
rect 22052 38587 22360 38596
rect 22756 38554 22784 39306
rect 22848 38554 22876 39510
rect 23112 39432 23164 39438
rect 23112 39374 23164 39380
rect 22744 38548 22796 38554
rect 22744 38490 22796 38496
rect 22836 38548 22888 38554
rect 22836 38490 22888 38496
rect 21824 38412 21876 38418
rect 21824 38354 21876 38360
rect 21836 38026 21864 38354
rect 22560 38208 22612 38214
rect 22560 38150 22612 38156
rect 22652 38208 22704 38214
rect 22652 38150 22704 38156
rect 21836 38010 21956 38026
rect 21836 38004 21968 38010
rect 21836 37998 21916 38004
rect 21916 37946 21968 37952
rect 20536 37868 20588 37874
rect 20536 37810 20588 37816
rect 21548 37868 21600 37874
rect 21548 37810 21600 37816
rect 21640 37868 21692 37874
rect 21640 37810 21692 37816
rect 19340 37800 19392 37806
rect 19340 37742 19392 37748
rect 19248 37460 19300 37466
rect 19248 37402 19300 37408
rect 19352 37262 19380 37742
rect 19432 37664 19484 37670
rect 19432 37606 19484 37612
rect 19340 37256 19392 37262
rect 19340 37198 19392 37204
rect 19352 36854 19380 37198
rect 19340 36848 19392 36854
rect 19340 36790 19392 36796
rect 19444 36718 19472 37606
rect 20548 37194 20576 37810
rect 21180 37664 21232 37670
rect 21180 37606 21232 37612
rect 22376 37664 22428 37670
rect 22376 37606 22428 37612
rect 21192 37466 21220 37606
rect 22052 37564 22360 37573
rect 22052 37562 22058 37564
rect 22114 37562 22138 37564
rect 22194 37562 22218 37564
rect 22274 37562 22298 37564
rect 22354 37562 22360 37564
rect 22114 37510 22116 37562
rect 22296 37510 22298 37562
rect 22052 37508 22058 37510
rect 22114 37508 22138 37510
rect 22194 37508 22218 37510
rect 22274 37508 22298 37510
rect 22354 37508 22360 37510
rect 22052 37499 22360 37508
rect 21180 37460 21232 37466
rect 21180 37402 21232 37408
rect 20628 37256 20680 37262
rect 20628 37198 20680 37204
rect 20720 37256 20772 37262
rect 20720 37198 20772 37204
rect 21916 37256 21968 37262
rect 21916 37198 21968 37204
rect 20536 37188 20588 37194
rect 20536 37130 20588 37136
rect 20548 36922 20576 37130
rect 20536 36916 20588 36922
rect 20536 36858 20588 36864
rect 19984 36780 20036 36786
rect 19984 36722 20036 36728
rect 19432 36712 19484 36718
rect 19432 36654 19484 36660
rect 18604 36236 18656 36242
rect 18604 36178 18656 36184
rect 19156 36236 19208 36242
rect 19156 36178 19208 36184
rect 18510 36136 18566 36145
rect 18510 36071 18566 36080
rect 18420 36032 18472 36038
rect 18420 35974 18472 35980
rect 17831 35932 18139 35941
rect 17831 35930 17837 35932
rect 17893 35930 17917 35932
rect 17973 35930 17997 35932
rect 18053 35930 18077 35932
rect 18133 35930 18139 35932
rect 17893 35878 17895 35930
rect 18075 35878 18077 35930
rect 17831 35876 17837 35878
rect 17893 35876 17917 35878
rect 17973 35876 17997 35878
rect 18053 35876 18077 35878
rect 18133 35876 18139 35878
rect 17831 35867 18139 35876
rect 17684 35692 17736 35698
rect 17684 35634 17736 35640
rect 17684 35080 17736 35086
rect 17684 35022 17736 35028
rect 18420 35080 18472 35086
rect 18420 35022 18472 35028
rect 17696 34202 17724 35022
rect 17831 34844 18139 34853
rect 17831 34842 17837 34844
rect 17893 34842 17917 34844
rect 17973 34842 17997 34844
rect 18053 34842 18077 34844
rect 18133 34842 18139 34844
rect 17893 34790 17895 34842
rect 18075 34790 18077 34842
rect 17831 34788 17837 34790
rect 17893 34788 17917 34790
rect 17973 34788 17997 34790
rect 18053 34788 18077 34790
rect 18133 34788 18139 34790
rect 17831 34779 18139 34788
rect 18432 34678 18460 35022
rect 18420 34672 18472 34678
rect 18420 34614 18472 34620
rect 17684 34196 17736 34202
rect 17684 34138 17736 34144
rect 17500 34128 17552 34134
rect 17500 34070 17552 34076
rect 18524 34082 18552 36071
rect 18616 34202 18644 36178
rect 18696 36168 18748 36174
rect 18696 36110 18748 36116
rect 19892 36168 19944 36174
rect 19892 36110 19944 36116
rect 18708 35834 18736 36110
rect 18696 35828 18748 35834
rect 18696 35770 18748 35776
rect 18972 35760 19024 35766
rect 18972 35702 19024 35708
rect 18880 35216 18932 35222
rect 18708 35176 18880 35204
rect 18604 34196 18656 34202
rect 18604 34138 18656 34144
rect 18524 34054 18644 34082
rect 18708 34066 18736 35176
rect 18880 35158 18932 35164
rect 18880 34740 18932 34746
rect 18880 34682 18932 34688
rect 18786 34640 18842 34649
rect 18786 34575 18842 34584
rect 18236 33992 18288 33998
rect 18236 33934 18288 33940
rect 17831 33756 18139 33765
rect 17831 33754 17837 33756
rect 17893 33754 17917 33756
rect 17973 33754 17997 33756
rect 18053 33754 18077 33756
rect 18133 33754 18139 33756
rect 17893 33702 17895 33754
rect 18075 33702 18077 33754
rect 17831 33700 17837 33702
rect 17893 33700 17917 33702
rect 17973 33700 17997 33702
rect 18053 33700 18077 33702
rect 18133 33700 18139 33702
rect 17831 33691 18139 33700
rect 18248 33658 18276 33934
rect 18512 33856 18564 33862
rect 18512 33798 18564 33804
rect 18236 33652 18288 33658
rect 18236 33594 18288 33600
rect 18052 33516 18104 33522
rect 18052 33458 18104 33464
rect 18064 33114 18092 33458
rect 18524 33386 18552 33798
rect 18512 33380 18564 33386
rect 18512 33322 18564 33328
rect 18052 33108 18104 33114
rect 18052 33050 18104 33056
rect 17408 33040 17460 33046
rect 17408 32982 17460 32988
rect 17776 32904 17828 32910
rect 17696 32864 17776 32892
rect 17592 32836 17644 32842
rect 17592 32778 17644 32784
rect 17604 32473 17632 32778
rect 17590 32464 17646 32473
rect 16304 32428 16356 32434
rect 16304 32370 16356 32376
rect 17132 32428 17184 32434
rect 17132 32370 17184 32376
rect 17224 32428 17276 32434
rect 17224 32370 17276 32376
rect 17316 32428 17368 32434
rect 17590 32399 17646 32408
rect 17316 32370 17368 32376
rect 16856 32224 16908 32230
rect 16856 32166 16908 32172
rect 16212 31884 16264 31890
rect 15752 30932 15804 30938
rect 15752 30874 15804 30880
rect 15752 30048 15804 30054
rect 15752 29990 15804 29996
rect 15660 29640 15712 29646
rect 15660 29582 15712 29588
rect 15764 29186 15792 29990
rect 15856 29646 15884 31878
rect 16212 31826 16264 31832
rect 15936 31816 15988 31822
rect 15936 31758 15988 31764
rect 16672 31816 16724 31822
rect 16672 31758 16724 31764
rect 15948 30326 15976 31758
rect 16028 31136 16080 31142
rect 16028 31078 16080 31084
rect 15936 30320 15988 30326
rect 15936 30262 15988 30268
rect 16040 30122 16068 31078
rect 16028 30116 16080 30122
rect 16028 30058 16080 30064
rect 16580 30116 16632 30122
rect 16580 30058 16632 30064
rect 15844 29640 15896 29646
rect 15934 29608 15990 29617
rect 15896 29588 15934 29594
rect 15844 29582 15934 29588
rect 15856 29566 15934 29582
rect 15934 29543 15990 29552
rect 16592 29238 16620 30058
rect 16684 29850 16712 31758
rect 16764 31272 16816 31278
rect 16764 31214 16816 31220
rect 16776 30938 16804 31214
rect 16764 30932 16816 30938
rect 16764 30874 16816 30880
rect 16764 30252 16816 30258
rect 16764 30194 16816 30200
rect 16672 29844 16724 29850
rect 16672 29786 16724 29792
rect 16776 29306 16804 30194
rect 16868 30190 16896 32166
rect 17132 31952 17184 31958
rect 17132 31894 17184 31900
rect 17040 31816 17092 31822
rect 17040 31758 17092 31764
rect 16948 31748 17000 31754
rect 16948 31690 17000 31696
rect 16960 31414 16988 31690
rect 16948 31408 17000 31414
rect 16948 31350 17000 31356
rect 16960 30938 16988 31350
rect 16948 30932 17000 30938
rect 16948 30874 17000 30880
rect 16960 30394 16988 30874
rect 17052 30410 17080 31758
rect 17144 30954 17172 31894
rect 17236 31754 17264 32370
rect 17696 32366 17724 32864
rect 18144 32904 18196 32910
rect 17880 32881 18144 32892
rect 17776 32846 17828 32852
rect 17866 32872 18144 32881
rect 18196 32872 18198 32881
rect 17922 32864 18142 32872
rect 17866 32807 17922 32816
rect 18142 32807 18198 32816
rect 17831 32668 18139 32677
rect 17831 32666 17837 32668
rect 17893 32666 17917 32668
rect 17973 32666 17997 32668
rect 18053 32666 18077 32668
rect 18133 32666 18139 32668
rect 17893 32614 17895 32666
rect 18075 32614 18077 32666
rect 17831 32612 17837 32614
rect 17893 32612 17917 32614
rect 17973 32612 17997 32614
rect 18053 32612 18077 32614
rect 18133 32612 18139 32614
rect 17831 32603 18139 32612
rect 17684 32360 17736 32366
rect 17684 32302 17736 32308
rect 17776 32360 17828 32366
rect 18236 32360 18288 32366
rect 17776 32302 17828 32308
rect 18234 32328 18236 32337
rect 18288 32328 18290 32337
rect 17592 32224 17644 32230
rect 17592 32166 17644 32172
rect 17604 31754 17632 32166
rect 17696 31958 17724 32302
rect 17788 31958 17816 32302
rect 18234 32263 18290 32272
rect 18420 32020 18472 32026
rect 18420 31962 18472 31968
rect 17684 31952 17736 31958
rect 17684 31894 17736 31900
rect 17776 31952 17828 31958
rect 17776 31894 17828 31900
rect 18236 31952 18288 31958
rect 18236 31894 18288 31900
rect 17224 31748 17276 31754
rect 17604 31726 17724 31754
rect 17224 31690 17276 31696
rect 17236 31482 17264 31690
rect 17500 31680 17552 31686
rect 17500 31622 17552 31628
rect 17592 31680 17644 31686
rect 17592 31622 17644 31628
rect 17224 31476 17276 31482
rect 17224 31418 17276 31424
rect 17144 30926 17356 30954
rect 17512 30938 17540 31622
rect 17604 31482 17632 31622
rect 17592 31476 17644 31482
rect 17592 31418 17644 31424
rect 17696 31328 17724 31726
rect 17831 31580 18139 31589
rect 17831 31578 17837 31580
rect 17893 31578 17917 31580
rect 17973 31578 17997 31580
rect 18053 31578 18077 31580
rect 18133 31578 18139 31580
rect 17893 31526 17895 31578
rect 18075 31526 18077 31578
rect 17831 31524 17837 31526
rect 17893 31524 17917 31526
rect 17973 31524 17997 31526
rect 18053 31524 18077 31526
rect 18133 31524 18139 31526
rect 17831 31515 18139 31524
rect 18248 31346 18276 31894
rect 17868 31340 17920 31346
rect 17696 31300 17868 31328
rect 17868 31282 17920 31288
rect 18236 31340 18288 31346
rect 18236 31282 18288 31288
rect 16948 30388 17000 30394
rect 17052 30382 17172 30410
rect 16948 30330 17000 30336
rect 16948 30252 17000 30258
rect 16948 30194 17000 30200
rect 17040 30252 17092 30258
rect 17144 30240 17172 30382
rect 17224 30252 17276 30258
rect 17144 30212 17224 30240
rect 17040 30194 17092 30200
rect 17224 30194 17276 30200
rect 16856 30184 16908 30190
rect 16856 30126 16908 30132
rect 16960 29306 16988 30194
rect 17052 30138 17080 30194
rect 17328 30138 17356 30926
rect 17500 30932 17552 30938
rect 17500 30874 17552 30880
rect 17684 30932 17736 30938
rect 17684 30874 17736 30880
rect 17500 30592 17552 30598
rect 17500 30534 17552 30540
rect 17512 30258 17540 30534
rect 17696 30394 17724 30874
rect 18236 30728 18288 30734
rect 18236 30670 18288 30676
rect 17831 30492 18139 30501
rect 17831 30490 17837 30492
rect 17893 30490 17917 30492
rect 17973 30490 17997 30492
rect 18053 30490 18077 30492
rect 18133 30490 18139 30492
rect 17893 30438 17895 30490
rect 18075 30438 18077 30490
rect 17831 30436 17837 30438
rect 17893 30436 17917 30438
rect 17973 30436 17997 30438
rect 18053 30436 18077 30438
rect 18133 30436 18139 30438
rect 17831 30427 18139 30436
rect 17684 30388 17736 30394
rect 17684 30330 17736 30336
rect 17500 30252 17552 30258
rect 17500 30194 17552 30200
rect 17052 30110 17356 30138
rect 17132 30048 17184 30054
rect 17132 29990 17184 29996
rect 16764 29300 16816 29306
rect 16764 29242 16816 29248
rect 16948 29300 17000 29306
rect 16948 29242 17000 29248
rect 15672 29158 15792 29186
rect 16580 29232 16632 29238
rect 16580 29174 16632 29180
rect 16028 29164 16080 29170
rect 15672 29034 15700 29158
rect 16028 29106 16080 29112
rect 16212 29164 16264 29170
rect 16212 29106 16264 29112
rect 16856 29164 16908 29170
rect 16856 29106 16908 29112
rect 15660 29028 15712 29034
rect 15660 28970 15712 28976
rect 15752 29028 15804 29034
rect 15752 28970 15804 28976
rect 15672 27334 15700 28970
rect 15764 27470 15792 28970
rect 16040 28558 16068 29106
rect 16224 28966 16252 29106
rect 16672 29096 16724 29102
rect 16672 29038 16724 29044
rect 16212 28960 16264 28966
rect 16212 28902 16264 28908
rect 16028 28552 16080 28558
rect 16028 28494 16080 28500
rect 15936 28076 15988 28082
rect 15936 28018 15988 28024
rect 15948 27674 15976 28018
rect 16040 27674 16068 28494
rect 16224 28218 16252 28902
rect 16684 28694 16712 29038
rect 16764 28960 16816 28966
rect 16764 28902 16816 28908
rect 16672 28688 16724 28694
rect 16672 28630 16724 28636
rect 16776 28558 16804 28902
rect 16868 28762 16896 29106
rect 16856 28756 16908 28762
rect 16856 28698 16908 28704
rect 16672 28552 16724 28558
rect 16672 28494 16724 28500
rect 16764 28552 16816 28558
rect 16764 28494 16816 28500
rect 16212 28212 16264 28218
rect 16212 28154 16264 28160
rect 16684 28014 16712 28494
rect 16488 28008 16540 28014
rect 16488 27950 16540 27956
rect 16672 28008 16724 28014
rect 16672 27950 16724 27956
rect 15936 27668 15988 27674
rect 15936 27610 15988 27616
rect 16028 27668 16080 27674
rect 16028 27610 16080 27616
rect 15752 27464 15804 27470
rect 15752 27406 15804 27412
rect 15660 27328 15712 27334
rect 15660 27270 15712 27276
rect 16500 27130 16528 27950
rect 17144 27470 17172 29990
rect 18142 29608 18198 29617
rect 17868 29572 17920 29578
rect 18052 29572 18104 29578
rect 17920 29532 18052 29560
rect 17868 29514 17920 29520
rect 18142 29543 18144 29552
rect 18052 29514 18104 29520
rect 18196 29543 18198 29552
rect 18144 29514 18196 29520
rect 17831 29404 18139 29413
rect 17831 29402 17837 29404
rect 17893 29402 17917 29404
rect 17973 29402 17997 29404
rect 18053 29402 18077 29404
rect 18133 29402 18139 29404
rect 17893 29350 17895 29402
rect 18075 29350 18077 29402
rect 17831 29348 17837 29350
rect 17893 29348 17917 29350
rect 17973 29348 17997 29350
rect 18053 29348 18077 29350
rect 18133 29348 18139 29350
rect 17831 29339 18139 29348
rect 18052 29232 18104 29238
rect 17498 29200 17554 29209
rect 18052 29174 18104 29180
rect 17498 29135 17554 29144
rect 17684 29164 17736 29170
rect 17512 28966 17540 29135
rect 17684 29106 17736 29112
rect 17592 29096 17644 29102
rect 17592 29038 17644 29044
rect 17500 28960 17552 28966
rect 17500 28902 17552 28908
rect 17316 28620 17368 28626
rect 17316 28562 17368 28568
rect 17328 28422 17356 28562
rect 17512 28490 17540 28902
rect 17604 28762 17632 29038
rect 17696 28762 17724 29106
rect 17592 28756 17644 28762
rect 17592 28698 17644 28704
rect 17684 28756 17736 28762
rect 17684 28698 17736 28704
rect 18064 28626 18092 29174
rect 18248 28626 18276 30670
rect 18326 30424 18382 30433
rect 18326 30359 18382 30368
rect 18340 29510 18368 30359
rect 18432 29850 18460 31962
rect 18524 31754 18552 33322
rect 18616 32910 18644 34054
rect 18696 34060 18748 34066
rect 18696 34002 18748 34008
rect 18708 33402 18736 34002
rect 18800 33930 18828 34575
rect 18788 33924 18840 33930
rect 18788 33866 18840 33872
rect 18708 33374 18828 33402
rect 18696 33312 18748 33318
rect 18696 33254 18748 33260
rect 18604 32904 18656 32910
rect 18604 32846 18656 32852
rect 18616 31958 18644 32846
rect 18604 31952 18656 31958
rect 18604 31894 18656 31900
rect 18708 31822 18736 33254
rect 18800 32774 18828 33374
rect 18788 32768 18840 32774
rect 18788 32710 18840 32716
rect 18800 32570 18828 32710
rect 18788 32564 18840 32570
rect 18788 32506 18840 32512
rect 18788 32428 18840 32434
rect 18788 32370 18840 32376
rect 18800 32026 18828 32370
rect 18788 32020 18840 32026
rect 18788 31962 18840 31968
rect 18892 31822 18920 34682
rect 18984 34610 19012 35702
rect 19904 35290 19932 36110
rect 19892 35284 19944 35290
rect 19892 35226 19944 35232
rect 19064 35080 19116 35086
rect 19064 35022 19116 35028
rect 19154 35048 19210 35057
rect 19076 34746 19104 35022
rect 19154 34983 19210 34992
rect 19064 34740 19116 34746
rect 19064 34682 19116 34688
rect 19168 34678 19196 34983
rect 19340 34740 19392 34746
rect 19340 34682 19392 34688
rect 19156 34672 19208 34678
rect 19156 34614 19208 34620
rect 18972 34604 19024 34610
rect 18972 34546 19024 34552
rect 19156 33856 19208 33862
rect 19156 33798 19208 33804
rect 19168 33590 19196 33798
rect 19156 33584 19208 33590
rect 19156 33526 19208 33532
rect 19352 32774 19380 34682
rect 19524 34604 19576 34610
rect 19524 34546 19576 34552
rect 19536 33862 19564 34546
rect 19800 33992 19852 33998
rect 19800 33934 19852 33940
rect 19524 33856 19576 33862
rect 19524 33798 19576 33804
rect 19708 33856 19760 33862
rect 19708 33798 19760 33804
rect 19720 33658 19748 33798
rect 19812 33658 19840 33934
rect 19708 33652 19760 33658
rect 19708 33594 19760 33600
rect 19800 33652 19852 33658
rect 19800 33594 19852 33600
rect 19524 33380 19576 33386
rect 19444 33340 19524 33368
rect 19340 32768 19392 32774
rect 19340 32710 19392 32716
rect 19154 32464 19210 32473
rect 19154 32399 19210 32408
rect 19168 32298 19196 32399
rect 18972 32292 19024 32298
rect 18972 32234 19024 32240
rect 19156 32292 19208 32298
rect 19156 32234 19208 32240
rect 18984 31822 19012 32234
rect 18696 31816 18748 31822
rect 18696 31758 18748 31764
rect 18880 31816 18932 31822
rect 18880 31758 18932 31764
rect 18972 31816 19024 31822
rect 18972 31758 19024 31764
rect 18512 31748 18564 31754
rect 18512 31690 18564 31696
rect 18788 31748 18840 31754
rect 18788 31690 18840 31696
rect 18524 31414 18552 31690
rect 18512 31408 18564 31414
rect 18512 31350 18564 31356
rect 18696 30252 18748 30258
rect 18696 30194 18748 30200
rect 18420 29844 18472 29850
rect 18420 29786 18472 29792
rect 18512 29776 18564 29782
rect 18512 29718 18564 29724
rect 18420 29640 18472 29646
rect 18420 29582 18472 29588
rect 18328 29504 18380 29510
rect 18328 29446 18380 29452
rect 18052 28620 18104 28626
rect 18052 28562 18104 28568
rect 18236 28620 18288 28626
rect 18236 28562 18288 28568
rect 17500 28484 17552 28490
rect 17500 28426 17552 28432
rect 17316 28416 17368 28422
rect 17316 28358 17368 28364
rect 17408 28416 17460 28422
rect 17408 28358 17460 28364
rect 17132 27464 17184 27470
rect 17132 27406 17184 27412
rect 16488 27124 16540 27130
rect 16488 27066 16540 27072
rect 15476 27056 15528 27062
rect 15476 26998 15528 27004
rect 15660 26988 15712 26994
rect 15660 26930 15712 26936
rect 15016 26852 15068 26858
rect 15016 26794 15068 26800
rect 15028 26518 15056 26794
rect 15108 26784 15160 26790
rect 15108 26726 15160 26732
rect 15384 26784 15436 26790
rect 15384 26726 15436 26732
rect 15568 26784 15620 26790
rect 15568 26726 15620 26732
rect 15016 26512 15068 26518
rect 15016 26454 15068 26460
rect 14884 26268 14964 26296
rect 14832 26250 14884 26256
rect 14844 25974 14872 26250
rect 14832 25968 14884 25974
rect 14832 25910 14884 25916
rect 14832 25696 14884 25702
rect 14832 25638 14884 25644
rect 14844 25498 14872 25638
rect 14832 25492 14884 25498
rect 14832 25434 14884 25440
rect 14924 25288 14976 25294
rect 14924 25230 14976 25236
rect 14936 24954 14964 25230
rect 14924 24948 14976 24954
rect 14924 24890 14976 24896
rect 14832 24812 14884 24818
rect 14832 24754 14884 24760
rect 14844 24410 14872 24754
rect 14832 24404 14884 24410
rect 14832 24346 14884 24352
rect 14844 23866 14872 24346
rect 14648 23860 14700 23866
rect 14648 23802 14700 23808
rect 14832 23860 14884 23866
rect 14832 23802 14884 23808
rect 14740 23724 14792 23730
rect 14740 23666 14792 23672
rect 14924 23724 14976 23730
rect 14924 23666 14976 23672
rect 14648 23520 14700 23526
rect 14648 23462 14700 23468
rect 14660 23118 14688 23462
rect 14752 23186 14780 23666
rect 14740 23180 14792 23186
rect 14740 23122 14792 23128
rect 14648 23112 14700 23118
rect 14648 23054 14700 23060
rect 14188 22772 14240 22778
rect 14188 22714 14240 22720
rect 14556 22772 14608 22778
rect 14556 22714 14608 22720
rect 14096 22636 14148 22642
rect 14096 22578 14148 22584
rect 14832 22636 14884 22642
rect 14832 22578 14884 22584
rect 13544 22568 13596 22574
rect 13544 22510 13596 22516
rect 14648 22500 14700 22506
rect 14648 22442 14700 22448
rect 14280 22432 14332 22438
rect 14280 22374 14332 22380
rect 13611 22332 13919 22341
rect 13611 22330 13617 22332
rect 13673 22330 13697 22332
rect 13753 22330 13777 22332
rect 13833 22330 13857 22332
rect 13913 22330 13919 22332
rect 13673 22278 13675 22330
rect 13855 22278 13857 22330
rect 13611 22276 13617 22278
rect 13673 22276 13697 22278
rect 13753 22276 13777 22278
rect 13833 22276 13857 22278
rect 13913 22276 13919 22278
rect 13611 22267 13919 22276
rect 13820 22024 13872 22030
rect 14188 22024 14240 22030
rect 13820 21966 13872 21972
rect 14016 21972 14188 21978
rect 14016 21966 14240 21972
rect 13728 21888 13780 21894
rect 13728 21830 13780 21836
rect 13740 21690 13768 21830
rect 13728 21684 13780 21690
rect 13728 21626 13780 21632
rect 13544 21548 13596 21554
rect 13544 21490 13596 21496
rect 13280 21406 13400 21434
rect 13452 21480 13504 21486
rect 13452 21422 13504 21428
rect 13084 21344 13136 21350
rect 13084 21286 13136 21292
rect 13176 21344 13228 21350
rect 13176 21286 13228 21292
rect 13096 21146 13124 21286
rect 13188 21146 13216 21286
rect 13084 21140 13136 21146
rect 13084 21082 13136 21088
rect 13176 21140 13228 21146
rect 13176 21082 13228 21088
rect 12992 20800 13044 20806
rect 12992 20742 13044 20748
rect 13096 20618 13124 21082
rect 13096 20590 13216 20618
rect 13084 20460 13136 20466
rect 13084 20402 13136 20408
rect 13096 20058 13124 20402
rect 13084 20052 13136 20058
rect 13084 19994 13136 20000
rect 13188 19854 13216 20590
rect 13280 19854 13308 21406
rect 13556 21298 13584 21490
rect 13832 21434 13860 21966
rect 14016 21950 14228 21966
rect 14016 21894 14044 21950
rect 14004 21888 14056 21894
rect 14004 21830 14056 21836
rect 14096 21888 14148 21894
rect 14096 21830 14148 21836
rect 14108 21622 14136 21830
rect 14096 21616 14148 21622
rect 14096 21558 14148 21564
rect 14200 21486 14228 21950
rect 14188 21480 14240 21486
rect 13832 21406 14136 21434
rect 14188 21422 14240 21428
rect 13464 21270 13584 21298
rect 13464 21146 13492 21270
rect 13611 21244 13919 21253
rect 13611 21242 13617 21244
rect 13673 21242 13697 21244
rect 13753 21242 13777 21244
rect 13833 21242 13857 21244
rect 13913 21242 13919 21244
rect 13673 21190 13675 21242
rect 13855 21190 13857 21242
rect 13611 21188 13617 21190
rect 13673 21188 13697 21190
rect 13753 21188 13777 21190
rect 13833 21188 13857 21190
rect 13913 21188 13919 21190
rect 13611 21179 13919 21188
rect 13452 21140 13504 21146
rect 13452 21082 13504 21088
rect 13464 20602 13492 21082
rect 14108 21078 14136 21406
rect 14200 21146 14228 21422
rect 14188 21140 14240 21146
rect 14188 21082 14240 21088
rect 14096 21072 14148 21078
rect 14096 21014 14148 21020
rect 13820 20936 13872 20942
rect 13820 20878 13872 20884
rect 13452 20596 13504 20602
rect 13452 20538 13504 20544
rect 13832 20330 13860 20878
rect 14096 20800 14148 20806
rect 14096 20742 14148 20748
rect 13820 20324 13872 20330
rect 13820 20266 13872 20272
rect 13611 20156 13919 20165
rect 13611 20154 13617 20156
rect 13673 20154 13697 20156
rect 13753 20154 13777 20156
rect 13833 20154 13857 20156
rect 13913 20154 13919 20156
rect 13673 20102 13675 20154
rect 13855 20102 13857 20154
rect 13611 20100 13617 20102
rect 13673 20100 13697 20102
rect 13753 20100 13777 20102
rect 13833 20100 13857 20102
rect 13913 20100 13919 20102
rect 13611 20091 13919 20100
rect 13176 19848 13228 19854
rect 13176 19790 13228 19796
rect 13268 19848 13320 19854
rect 13268 19790 13320 19796
rect 12808 19712 12860 19718
rect 12808 19654 12860 19660
rect 12440 19508 12492 19514
rect 12440 19450 12492 19456
rect 11060 19372 11112 19378
rect 11060 19314 11112 19320
rect 11888 19372 11940 19378
rect 11888 19314 11940 19320
rect 12348 19372 12400 19378
rect 12348 19314 12400 19320
rect 14108 19310 14136 20742
rect 14200 20602 14228 21082
rect 14292 21010 14320 22374
rect 14372 22160 14424 22166
rect 14424 22108 14504 22114
rect 14372 22102 14504 22108
rect 14384 22086 14504 22102
rect 14476 21418 14504 22086
rect 14660 22030 14688 22442
rect 14648 22024 14700 22030
rect 14648 21966 14700 21972
rect 14740 22024 14792 22030
rect 14740 21966 14792 21972
rect 14752 21536 14780 21966
rect 14844 21894 14872 22578
rect 14936 22094 14964 23666
rect 15028 23254 15056 26454
rect 15120 25906 15148 26726
rect 15200 26240 15252 26246
rect 15200 26182 15252 26188
rect 15212 25974 15240 26182
rect 15200 25968 15252 25974
rect 15252 25928 15332 25956
rect 15200 25910 15252 25916
rect 15108 25900 15160 25906
rect 15108 25842 15160 25848
rect 15120 25294 15148 25842
rect 15200 25696 15252 25702
rect 15200 25638 15252 25644
rect 15212 25498 15240 25638
rect 15200 25492 15252 25498
rect 15200 25434 15252 25440
rect 15304 25430 15332 25928
rect 15396 25906 15424 26726
rect 15476 26240 15528 26246
rect 15476 26182 15528 26188
rect 15384 25900 15436 25906
rect 15384 25842 15436 25848
rect 15488 25786 15516 26182
rect 15580 25974 15608 26726
rect 15672 25974 15700 26930
rect 15936 26920 15988 26926
rect 15936 26862 15988 26868
rect 15752 26784 15804 26790
rect 15752 26726 15804 26732
rect 15844 26784 15896 26790
rect 15844 26726 15896 26732
rect 15568 25968 15620 25974
rect 15568 25910 15620 25916
rect 15660 25968 15712 25974
rect 15660 25910 15712 25916
rect 15764 25906 15792 26726
rect 15856 26382 15884 26726
rect 15844 26376 15896 26382
rect 15844 26318 15896 26324
rect 15752 25900 15804 25906
rect 15752 25842 15804 25848
rect 15488 25758 15608 25786
rect 15292 25424 15344 25430
rect 15292 25366 15344 25372
rect 15108 25288 15160 25294
rect 15108 25230 15160 25236
rect 15108 24880 15160 24886
rect 15108 24822 15160 24828
rect 15120 23730 15148 24822
rect 15384 24744 15436 24750
rect 15384 24686 15436 24692
rect 15396 24410 15424 24686
rect 15384 24404 15436 24410
rect 15384 24346 15436 24352
rect 15292 24200 15344 24206
rect 15292 24142 15344 24148
rect 15304 23798 15332 24142
rect 15292 23792 15344 23798
rect 15292 23734 15344 23740
rect 15108 23724 15160 23730
rect 15108 23666 15160 23672
rect 15016 23248 15068 23254
rect 15016 23190 15068 23196
rect 15304 23118 15332 23734
rect 15396 23594 15424 24346
rect 15476 24064 15528 24070
rect 15476 24006 15528 24012
rect 15384 23588 15436 23594
rect 15384 23530 15436 23536
rect 15292 23112 15344 23118
rect 15292 23054 15344 23060
rect 15488 22778 15516 24006
rect 15580 23769 15608 25758
rect 15948 25702 15976 26862
rect 16396 26376 16448 26382
rect 16396 26318 16448 26324
rect 16408 25838 16436 26318
rect 16500 26314 16528 27066
rect 17132 26920 17184 26926
rect 17132 26862 17184 26868
rect 17040 26784 17092 26790
rect 17040 26726 17092 26732
rect 16672 26444 16724 26450
rect 16672 26386 16724 26392
rect 16488 26308 16540 26314
rect 16488 26250 16540 26256
rect 16684 25906 16712 26386
rect 17052 26382 17080 26726
rect 17144 26586 17172 26862
rect 17132 26580 17184 26586
rect 17132 26522 17184 26528
rect 17040 26376 17092 26382
rect 17040 26318 17092 26324
rect 16948 26240 17000 26246
rect 16948 26182 17000 26188
rect 17132 26240 17184 26246
rect 17132 26182 17184 26188
rect 16960 25906 16988 26182
rect 16672 25900 16724 25906
rect 16592 25860 16672 25888
rect 16120 25832 16172 25838
rect 16120 25774 16172 25780
rect 16396 25832 16448 25838
rect 16396 25774 16448 25780
rect 15936 25696 15988 25702
rect 15936 25638 15988 25644
rect 15660 25288 15712 25294
rect 15660 25230 15712 25236
rect 15672 24750 15700 25230
rect 16132 25226 16160 25774
rect 16488 25696 16540 25702
rect 16488 25638 16540 25644
rect 16500 25294 16528 25638
rect 16592 25498 16620 25860
rect 16672 25842 16724 25848
rect 16948 25900 17000 25906
rect 16948 25842 17000 25848
rect 16580 25492 16632 25498
rect 16580 25434 16632 25440
rect 16488 25288 16540 25294
rect 16488 25230 16540 25236
rect 16120 25220 16172 25226
rect 16120 25162 16172 25168
rect 16120 24812 16172 24818
rect 16120 24754 16172 24760
rect 15660 24744 15712 24750
rect 15660 24686 15712 24692
rect 15844 24744 15896 24750
rect 15844 24686 15896 24692
rect 15936 24744 15988 24750
rect 15936 24686 15988 24692
rect 15660 24608 15712 24614
rect 15660 24550 15712 24556
rect 15752 24608 15804 24614
rect 15752 24550 15804 24556
rect 15672 23866 15700 24550
rect 15764 23866 15792 24550
rect 15856 23866 15884 24686
rect 15948 24070 15976 24686
rect 15936 24064 15988 24070
rect 15936 24006 15988 24012
rect 16132 23866 16160 24754
rect 17040 24676 17092 24682
rect 17040 24618 17092 24624
rect 15660 23860 15712 23866
rect 15660 23802 15712 23808
rect 15752 23860 15804 23866
rect 15752 23802 15804 23808
rect 15844 23860 15896 23866
rect 15844 23802 15896 23808
rect 16120 23860 16172 23866
rect 16120 23802 16172 23808
rect 15566 23760 15622 23769
rect 15566 23695 15568 23704
rect 15620 23695 15622 23704
rect 15568 23666 15620 23672
rect 17052 23118 17080 24618
rect 16120 23112 16172 23118
rect 16120 23054 16172 23060
rect 17040 23112 17092 23118
rect 17040 23054 17092 23060
rect 15568 22976 15620 22982
rect 15568 22918 15620 22924
rect 15580 22778 15608 22918
rect 16132 22778 16160 23054
rect 15476 22772 15528 22778
rect 15476 22714 15528 22720
rect 15568 22772 15620 22778
rect 15568 22714 15620 22720
rect 16120 22772 16172 22778
rect 16120 22714 16172 22720
rect 16488 22636 16540 22642
rect 16488 22578 16540 22584
rect 16672 22636 16724 22642
rect 16672 22578 16724 22584
rect 15108 22432 15160 22438
rect 15108 22374 15160 22380
rect 16120 22432 16172 22438
rect 16120 22374 16172 22380
rect 16396 22432 16448 22438
rect 16396 22374 16448 22380
rect 14936 22066 15056 22094
rect 14832 21888 14884 21894
rect 14832 21830 14884 21836
rect 15028 21570 15056 22066
rect 15120 22030 15148 22374
rect 16132 22234 16160 22374
rect 16120 22228 16172 22234
rect 16120 22170 16172 22176
rect 15292 22160 15344 22166
rect 15292 22102 15344 22108
rect 15108 22024 15160 22030
rect 15108 21966 15160 21972
rect 15200 22024 15252 22030
rect 15200 21966 15252 21972
rect 15120 21690 15148 21966
rect 15108 21684 15160 21690
rect 15108 21626 15160 21632
rect 15028 21554 15148 21570
rect 15212 21554 15240 21966
rect 14924 21548 14976 21554
rect 14752 21508 14872 21536
rect 14464 21412 14516 21418
rect 14464 21354 14516 21360
rect 14740 21344 14792 21350
rect 14740 21286 14792 21292
rect 14752 21146 14780 21286
rect 14844 21146 14872 21508
rect 14924 21490 14976 21496
rect 15016 21548 15148 21554
rect 15068 21542 15148 21548
rect 15016 21490 15068 21496
rect 14740 21140 14792 21146
rect 14740 21082 14792 21088
rect 14832 21140 14884 21146
rect 14832 21082 14884 21088
rect 14464 21072 14516 21078
rect 14464 21014 14516 21020
rect 14280 21004 14332 21010
rect 14280 20946 14332 20952
rect 14188 20596 14240 20602
rect 14188 20538 14240 20544
rect 14372 20392 14424 20398
rect 14372 20334 14424 20340
rect 14384 19514 14412 20334
rect 14476 19514 14504 21014
rect 14936 20602 14964 21490
rect 15120 21350 15148 21542
rect 15200 21548 15252 21554
rect 15200 21490 15252 21496
rect 15108 21344 15160 21350
rect 15108 21286 15160 21292
rect 15200 21072 15252 21078
rect 15200 21014 15252 21020
rect 15212 20602 15240 21014
rect 14924 20596 14976 20602
rect 14924 20538 14976 20544
rect 15200 20596 15252 20602
rect 15200 20538 15252 20544
rect 14556 20324 14608 20330
rect 14556 20266 14608 20272
rect 14568 20058 14596 20266
rect 14556 20052 14608 20058
rect 14556 19994 14608 20000
rect 14372 19508 14424 19514
rect 14372 19450 14424 19456
rect 14464 19508 14516 19514
rect 14464 19450 14516 19456
rect 14568 19446 14596 19994
rect 14556 19440 14608 19446
rect 14556 19382 14608 19388
rect 14936 19378 14964 20538
rect 15016 20256 15068 20262
rect 15016 20198 15068 20204
rect 15028 19854 15056 20198
rect 15304 20058 15332 22102
rect 15844 22024 15896 22030
rect 15844 21966 15896 21972
rect 15384 21888 15436 21894
rect 15384 21830 15436 21836
rect 15396 21078 15424 21830
rect 15476 21684 15528 21690
rect 15476 21626 15528 21632
rect 15488 21146 15516 21626
rect 15660 21480 15712 21486
rect 15660 21422 15712 21428
rect 15672 21146 15700 21422
rect 15752 21344 15804 21350
rect 15752 21286 15804 21292
rect 15764 21146 15792 21286
rect 15476 21140 15528 21146
rect 15476 21082 15528 21088
rect 15660 21140 15712 21146
rect 15660 21082 15712 21088
rect 15752 21140 15804 21146
rect 15752 21082 15804 21088
rect 15856 21078 15884 21966
rect 15384 21072 15436 21078
rect 15384 21014 15436 21020
rect 15844 21072 15896 21078
rect 15844 21014 15896 21020
rect 15384 20868 15436 20874
rect 15384 20810 15436 20816
rect 15660 20868 15712 20874
rect 15660 20810 15712 20816
rect 15396 20602 15424 20810
rect 15384 20596 15436 20602
rect 15384 20538 15436 20544
rect 15672 20058 15700 20810
rect 16408 20602 16436 22374
rect 16500 21690 16528 22578
rect 16488 21684 16540 21690
rect 16488 21626 16540 21632
rect 16684 21554 16712 22578
rect 17144 22574 17172 26182
rect 17328 24818 17356 28358
rect 17420 28082 17448 28358
rect 17831 28316 18139 28325
rect 17831 28314 17837 28316
rect 17893 28314 17917 28316
rect 17973 28314 17997 28316
rect 18053 28314 18077 28316
rect 18133 28314 18139 28316
rect 17893 28262 17895 28314
rect 18075 28262 18077 28314
rect 17831 28260 17837 28262
rect 17893 28260 17917 28262
rect 17973 28260 17997 28262
rect 18053 28260 18077 28262
rect 18133 28260 18139 28262
rect 17831 28251 18139 28260
rect 18248 28218 18276 28562
rect 18236 28212 18288 28218
rect 18236 28154 18288 28160
rect 17408 28076 17460 28082
rect 17408 28018 17460 28024
rect 17776 28076 17828 28082
rect 17776 28018 17828 28024
rect 17788 27470 17816 28018
rect 17776 27464 17828 27470
rect 17696 27424 17776 27452
rect 17408 27056 17460 27062
rect 17408 26998 17460 27004
rect 17420 25498 17448 26998
rect 17592 26852 17644 26858
rect 17592 26794 17644 26800
rect 17408 25492 17460 25498
rect 17408 25434 17460 25440
rect 17420 24954 17448 25434
rect 17408 24948 17460 24954
rect 17408 24890 17460 24896
rect 17604 24818 17632 26794
rect 17696 26450 17724 27424
rect 17776 27406 17828 27412
rect 17831 27228 18139 27237
rect 17831 27226 17837 27228
rect 17893 27226 17917 27228
rect 17973 27226 17997 27228
rect 18053 27226 18077 27228
rect 18133 27226 18139 27228
rect 17893 27174 17895 27226
rect 18075 27174 18077 27226
rect 17831 27172 17837 27174
rect 17893 27172 17917 27174
rect 17973 27172 17997 27174
rect 18053 27172 18077 27174
rect 18133 27172 18139 27174
rect 17831 27163 18139 27172
rect 17776 26784 17828 26790
rect 17776 26726 17828 26732
rect 17684 26444 17736 26450
rect 17684 26386 17736 26392
rect 17788 26382 17816 26726
rect 17776 26376 17828 26382
rect 17776 26318 17828 26324
rect 17831 26140 18139 26149
rect 17831 26138 17837 26140
rect 17893 26138 17917 26140
rect 17973 26138 17997 26140
rect 18053 26138 18077 26140
rect 18133 26138 18139 26140
rect 17893 26086 17895 26138
rect 18075 26086 18077 26138
rect 17831 26084 17837 26086
rect 17893 26084 17917 26086
rect 17973 26084 17997 26086
rect 18053 26084 18077 26086
rect 18133 26084 18139 26086
rect 17831 26075 18139 26084
rect 18340 25906 18368 29446
rect 18432 29306 18460 29582
rect 18420 29300 18472 29306
rect 18420 29242 18472 29248
rect 18524 29238 18552 29718
rect 18604 29640 18656 29646
rect 18708 29628 18736 30194
rect 18800 30122 18828 31690
rect 18972 31136 19024 31142
rect 18972 31078 19024 31084
rect 18984 30734 19012 31078
rect 19352 30734 19380 32710
rect 19444 32434 19472 33340
rect 19524 33322 19576 33328
rect 19616 33380 19668 33386
rect 19616 33322 19668 33328
rect 19628 33114 19656 33322
rect 19800 33312 19852 33318
rect 19800 33254 19852 33260
rect 19616 33108 19668 33114
rect 19616 33050 19668 33056
rect 19524 32904 19576 32910
rect 19522 32872 19524 32881
rect 19576 32872 19578 32881
rect 19522 32807 19578 32816
rect 19628 32434 19656 33050
rect 19812 33046 19840 33254
rect 19800 33040 19852 33046
rect 19800 32982 19852 32988
rect 19800 32768 19852 32774
rect 19800 32710 19852 32716
rect 19812 32434 19840 32710
rect 19432 32428 19484 32434
rect 19432 32370 19484 32376
rect 19616 32428 19668 32434
rect 19616 32370 19668 32376
rect 19800 32428 19852 32434
rect 19800 32370 19852 32376
rect 19444 32337 19472 32370
rect 19430 32328 19486 32337
rect 19430 32263 19486 32272
rect 19432 32224 19484 32230
rect 19432 32166 19484 32172
rect 19444 31890 19472 32166
rect 19708 32020 19760 32026
rect 19708 31962 19760 31968
rect 19432 31884 19484 31890
rect 19432 31826 19484 31832
rect 19720 31822 19748 31962
rect 19524 31816 19576 31822
rect 19708 31816 19760 31822
rect 19576 31764 19656 31770
rect 19524 31758 19656 31764
rect 19708 31758 19760 31764
rect 19536 31742 19656 31758
rect 19628 31634 19656 31742
rect 19628 31606 19748 31634
rect 19616 31476 19668 31482
rect 19616 31418 19668 31424
rect 19628 30734 19656 31418
rect 18972 30728 19024 30734
rect 18972 30670 19024 30676
rect 19340 30728 19392 30734
rect 19616 30728 19668 30734
rect 19392 30676 19472 30682
rect 19340 30670 19472 30676
rect 19616 30670 19668 30676
rect 19352 30654 19472 30670
rect 19444 30258 19472 30654
rect 19524 30660 19576 30666
rect 19524 30602 19576 30608
rect 18880 30252 18932 30258
rect 19156 30252 19208 30258
rect 18932 30212 19012 30240
rect 18880 30194 18932 30200
rect 18984 30122 19012 30212
rect 19156 30194 19208 30200
rect 19432 30252 19484 30258
rect 19432 30194 19484 30200
rect 18788 30116 18840 30122
rect 18788 30058 18840 30064
rect 18972 30116 19024 30122
rect 18972 30058 19024 30064
rect 18880 30048 18932 30054
rect 18880 29990 18932 29996
rect 18656 29600 18736 29628
rect 18604 29582 18656 29588
rect 18604 29504 18656 29510
rect 18604 29446 18656 29452
rect 18696 29504 18748 29510
rect 18696 29446 18748 29452
rect 18616 29306 18644 29446
rect 18604 29300 18656 29306
rect 18604 29242 18656 29248
rect 18512 29232 18564 29238
rect 18708 29186 18736 29446
rect 18892 29306 18920 29990
rect 19168 29850 19196 30194
rect 19536 30122 19564 30602
rect 19524 30116 19576 30122
rect 19524 30058 19576 30064
rect 19340 30048 19392 30054
rect 19340 29990 19392 29996
rect 19352 29850 19380 29990
rect 19156 29844 19208 29850
rect 19156 29786 19208 29792
rect 19340 29844 19392 29850
rect 19340 29786 19392 29792
rect 19064 29776 19116 29782
rect 19720 29730 19748 31606
rect 19800 31272 19852 31278
rect 19800 31214 19852 31220
rect 19812 30802 19840 31214
rect 19800 30796 19852 30802
rect 19800 30738 19852 30744
rect 19892 30728 19944 30734
rect 19892 30670 19944 30676
rect 19904 30326 19932 30670
rect 19996 30433 20024 36722
rect 20536 36712 20588 36718
rect 20536 36654 20588 36660
rect 20076 36576 20128 36582
rect 20076 36518 20128 36524
rect 20088 35766 20116 36518
rect 20444 36304 20496 36310
rect 20444 36246 20496 36252
rect 20168 36032 20220 36038
rect 20168 35974 20220 35980
rect 20076 35760 20128 35766
rect 20076 35702 20128 35708
rect 20180 34202 20208 35974
rect 20456 35834 20484 36246
rect 20548 35834 20576 36654
rect 20640 36242 20668 37198
rect 20732 36582 20760 37198
rect 21088 37120 21140 37126
rect 21088 37062 21140 37068
rect 21640 37120 21692 37126
rect 21640 37062 21692 37068
rect 20720 36576 20772 36582
rect 20720 36518 20772 36524
rect 20628 36236 20680 36242
rect 20628 36178 20680 36184
rect 20732 36174 20760 36518
rect 20812 36236 20864 36242
rect 20812 36178 20864 36184
rect 20720 36168 20772 36174
rect 20720 36110 20772 36116
rect 20444 35828 20496 35834
rect 20444 35770 20496 35776
rect 20536 35828 20588 35834
rect 20536 35770 20588 35776
rect 20824 35086 20852 36178
rect 20904 36032 20956 36038
rect 20904 35974 20956 35980
rect 20916 35290 20944 35974
rect 21100 35834 21128 37062
rect 21652 36922 21680 37062
rect 21928 36922 21956 37198
rect 21640 36916 21692 36922
rect 21640 36858 21692 36864
rect 21916 36916 21968 36922
rect 21916 36858 21968 36864
rect 21364 36100 21416 36106
rect 21364 36042 21416 36048
rect 21376 35834 21404 36042
rect 21824 36032 21876 36038
rect 21824 35974 21876 35980
rect 21836 35834 21864 35974
rect 21088 35828 21140 35834
rect 21088 35770 21140 35776
rect 21364 35828 21416 35834
rect 21364 35770 21416 35776
rect 21824 35828 21876 35834
rect 21824 35770 21876 35776
rect 21928 35630 21956 36858
rect 22052 36476 22360 36485
rect 22052 36474 22058 36476
rect 22114 36474 22138 36476
rect 22194 36474 22218 36476
rect 22274 36474 22298 36476
rect 22354 36474 22360 36476
rect 22114 36422 22116 36474
rect 22296 36422 22298 36474
rect 22052 36420 22058 36422
rect 22114 36420 22138 36422
rect 22194 36420 22218 36422
rect 22274 36420 22298 36422
rect 22354 36420 22360 36422
rect 22052 36411 22360 36420
rect 22192 36032 22244 36038
rect 22192 35974 22244 35980
rect 22284 36032 22336 36038
rect 22284 35974 22336 35980
rect 21916 35624 21968 35630
rect 21916 35566 21968 35572
rect 21272 35488 21324 35494
rect 21272 35430 21324 35436
rect 21824 35488 21876 35494
rect 21824 35430 21876 35436
rect 20904 35284 20956 35290
rect 20904 35226 20956 35232
rect 20812 35080 20864 35086
rect 20812 35022 20864 35028
rect 21284 35018 21312 35430
rect 21836 35086 21864 35430
rect 21928 35290 21956 35566
rect 22204 35562 22232 35974
rect 22296 35698 22324 35974
rect 22284 35692 22336 35698
rect 22284 35634 22336 35640
rect 22192 35556 22244 35562
rect 22192 35498 22244 35504
rect 22052 35388 22360 35397
rect 22052 35386 22058 35388
rect 22114 35386 22138 35388
rect 22194 35386 22218 35388
rect 22274 35386 22298 35388
rect 22354 35386 22360 35388
rect 22114 35334 22116 35386
rect 22296 35334 22298 35386
rect 22052 35332 22058 35334
rect 22114 35332 22138 35334
rect 22194 35332 22218 35334
rect 22274 35332 22298 35334
rect 22354 35332 22360 35334
rect 22052 35323 22360 35332
rect 21916 35284 21968 35290
rect 21916 35226 21968 35232
rect 22388 35154 22416 37606
rect 22468 37460 22520 37466
rect 22468 37402 22520 37408
rect 22480 35834 22508 37402
rect 22572 37262 22600 38150
rect 22664 37466 22692 38150
rect 22652 37460 22704 37466
rect 22652 37402 22704 37408
rect 22560 37256 22612 37262
rect 22560 37198 22612 37204
rect 23020 37120 23072 37126
rect 23020 37062 23072 37068
rect 23032 36854 23060 37062
rect 23020 36848 23072 36854
rect 23020 36790 23072 36796
rect 22468 35828 22520 35834
rect 22468 35770 22520 35776
rect 22468 35692 22520 35698
rect 22468 35634 22520 35640
rect 22376 35148 22428 35154
rect 22376 35090 22428 35096
rect 22480 35086 22508 35634
rect 22560 35556 22612 35562
rect 22560 35498 22612 35504
rect 22572 35290 22600 35498
rect 22652 35488 22704 35494
rect 22652 35430 22704 35436
rect 22560 35284 22612 35290
rect 22560 35226 22612 35232
rect 21824 35080 21876 35086
rect 21824 35022 21876 35028
rect 22468 35080 22520 35086
rect 22468 35022 22520 35028
rect 22560 35080 22612 35086
rect 22560 35022 22612 35028
rect 21272 35012 21324 35018
rect 21272 34954 21324 34960
rect 20628 34740 20680 34746
rect 20628 34682 20680 34688
rect 20640 34610 20668 34682
rect 22468 34672 22520 34678
rect 22468 34614 22520 34620
rect 20628 34604 20680 34610
rect 20628 34546 20680 34552
rect 20812 34400 20864 34406
rect 20812 34342 20864 34348
rect 21364 34400 21416 34406
rect 21364 34342 21416 34348
rect 20168 34196 20220 34202
rect 20168 34138 20220 34144
rect 20824 33998 20852 34342
rect 20812 33992 20864 33998
rect 20812 33934 20864 33940
rect 20720 33856 20772 33862
rect 20720 33798 20772 33804
rect 20996 33856 21048 33862
rect 20996 33798 21048 33804
rect 20168 33516 20220 33522
rect 20168 33458 20220 33464
rect 20180 33318 20208 33458
rect 20168 33312 20220 33318
rect 20168 33254 20220 33260
rect 20444 33312 20496 33318
rect 20444 33254 20496 33260
rect 20456 33114 20484 33254
rect 20444 33108 20496 33114
rect 20732 33096 20760 33798
rect 21008 33522 21036 33798
rect 21376 33590 21404 34342
rect 22052 34300 22360 34309
rect 22052 34298 22058 34300
rect 22114 34298 22138 34300
rect 22194 34298 22218 34300
rect 22274 34298 22298 34300
rect 22354 34298 22360 34300
rect 22114 34246 22116 34298
rect 22296 34246 22298 34298
rect 22052 34244 22058 34246
rect 22114 34244 22138 34246
rect 22194 34244 22218 34246
rect 22274 34244 22298 34246
rect 22354 34244 22360 34246
rect 22052 34235 22360 34244
rect 22284 33924 22336 33930
rect 22284 33866 22336 33872
rect 21364 33584 21416 33590
rect 21364 33526 21416 33532
rect 20996 33516 21048 33522
rect 20996 33458 21048 33464
rect 21088 33312 21140 33318
rect 21088 33254 21140 33260
rect 21100 33114 21128 33254
rect 20444 33050 20496 33056
rect 20640 33068 20760 33096
rect 21088 33108 21140 33114
rect 20076 33040 20128 33046
rect 20076 32982 20128 32988
rect 20088 32910 20116 32982
rect 20076 32904 20128 32910
rect 20076 32846 20128 32852
rect 20352 32904 20404 32910
rect 20352 32846 20404 32852
rect 20640 32858 20668 33068
rect 21088 33050 21140 33056
rect 20720 32972 20772 32978
rect 20772 32932 20852 32960
rect 20720 32914 20772 32920
rect 20088 32434 20116 32846
rect 20260 32768 20312 32774
rect 20260 32710 20312 32716
rect 20076 32428 20128 32434
rect 20076 32370 20128 32376
rect 20076 32292 20128 32298
rect 20076 32234 20128 32240
rect 20088 31822 20116 32234
rect 20272 32026 20300 32710
rect 20364 32570 20392 32846
rect 20640 32830 20760 32858
rect 20352 32564 20404 32570
rect 20352 32506 20404 32512
rect 20260 32020 20312 32026
rect 20260 31962 20312 31968
rect 20076 31816 20128 31822
rect 20076 31758 20128 31764
rect 20352 31136 20404 31142
rect 20352 31078 20404 31084
rect 20260 30728 20312 30734
rect 20260 30670 20312 30676
rect 19982 30424 20038 30433
rect 20272 30394 20300 30670
rect 19982 30359 20038 30368
rect 20260 30388 20312 30394
rect 20260 30330 20312 30336
rect 19892 30320 19944 30326
rect 19892 30262 19944 30268
rect 20364 30258 20392 31078
rect 20444 30728 20496 30734
rect 20444 30670 20496 30676
rect 20456 30394 20484 30670
rect 20536 30592 20588 30598
rect 20536 30534 20588 30540
rect 20548 30433 20576 30534
rect 20534 30424 20590 30433
rect 20444 30388 20496 30394
rect 20534 30359 20590 30368
rect 20444 30330 20496 30336
rect 20168 30252 20220 30258
rect 20168 30194 20220 30200
rect 20352 30252 20404 30258
rect 20352 30194 20404 30200
rect 19892 30184 19944 30190
rect 19892 30126 19944 30132
rect 19904 29850 19932 30126
rect 19892 29844 19944 29850
rect 19892 29786 19944 29792
rect 19064 29718 19116 29724
rect 19076 29646 19104 29718
rect 19168 29702 19748 29730
rect 19984 29776 20036 29782
rect 19984 29718 20036 29724
rect 18972 29640 19024 29646
rect 18972 29582 19024 29588
rect 19064 29640 19116 29646
rect 19064 29582 19116 29588
rect 18984 29306 19012 29582
rect 18880 29300 18932 29306
rect 18880 29242 18932 29248
rect 18972 29300 19024 29306
rect 18972 29242 19024 29248
rect 18564 29180 18736 29186
rect 18512 29174 18736 29180
rect 18524 29158 18736 29174
rect 18604 28960 18656 28966
rect 18604 28902 18656 28908
rect 18616 28626 18644 28902
rect 18604 28620 18656 28626
rect 18604 28562 18656 28568
rect 18420 28416 18472 28422
rect 18420 28358 18472 28364
rect 18432 28082 18460 28358
rect 18420 28076 18472 28082
rect 18420 28018 18472 28024
rect 18420 26920 18472 26926
rect 18420 26862 18472 26868
rect 18432 26382 18460 26862
rect 18420 26376 18472 26382
rect 18420 26318 18472 26324
rect 18328 25900 18380 25906
rect 18328 25842 18380 25848
rect 18432 25770 18460 26318
rect 18604 26240 18656 26246
rect 18604 26182 18656 26188
rect 18420 25764 18472 25770
rect 18420 25706 18472 25712
rect 18616 25158 18644 26182
rect 18604 25152 18656 25158
rect 18604 25094 18656 25100
rect 17831 25052 18139 25061
rect 17831 25050 17837 25052
rect 17893 25050 17917 25052
rect 17973 25050 17997 25052
rect 18053 25050 18077 25052
rect 18133 25050 18139 25052
rect 17893 24998 17895 25050
rect 18075 24998 18077 25050
rect 17831 24996 17837 24998
rect 17893 24996 17917 24998
rect 17973 24996 17997 24998
rect 18053 24996 18077 24998
rect 18133 24996 18139 24998
rect 17831 24987 18139 24996
rect 17316 24812 17368 24818
rect 17316 24754 17368 24760
rect 17592 24812 17644 24818
rect 17592 24754 17644 24760
rect 18144 24812 18196 24818
rect 18144 24754 18196 24760
rect 18236 24812 18288 24818
rect 18236 24754 18288 24760
rect 17328 23882 17356 24754
rect 18156 24410 18184 24754
rect 18144 24404 18196 24410
rect 18144 24346 18196 24352
rect 17684 24200 17736 24206
rect 17684 24142 17736 24148
rect 17500 24132 17552 24138
rect 17500 24074 17552 24080
rect 17328 23854 17448 23882
rect 17512 23866 17540 24074
rect 17316 23724 17368 23730
rect 17316 23666 17368 23672
rect 17328 23322 17356 23666
rect 17316 23316 17368 23322
rect 17316 23258 17368 23264
rect 17420 23118 17448 23854
rect 17500 23860 17552 23866
rect 17500 23802 17552 23808
rect 17696 23526 17724 24142
rect 18248 24070 18276 24754
rect 18328 24608 18380 24614
rect 18328 24550 18380 24556
rect 18236 24064 18288 24070
rect 18236 24006 18288 24012
rect 17831 23964 18139 23973
rect 17831 23962 17837 23964
rect 17893 23962 17917 23964
rect 17973 23962 17997 23964
rect 18053 23962 18077 23964
rect 18133 23962 18139 23964
rect 17893 23910 17895 23962
rect 18075 23910 18077 23962
rect 17831 23908 17837 23910
rect 17893 23908 17917 23910
rect 17973 23908 17997 23910
rect 18053 23908 18077 23910
rect 18133 23908 18139 23910
rect 17831 23899 18139 23908
rect 18248 23746 18276 24006
rect 18340 23866 18368 24550
rect 18616 24342 18644 25094
rect 18604 24336 18656 24342
rect 18604 24278 18656 24284
rect 18708 24274 18736 29158
rect 19076 27334 19104 29582
rect 19168 29510 19196 29702
rect 19340 29640 19392 29646
rect 19340 29582 19392 29588
rect 19156 29504 19208 29510
rect 19156 29446 19208 29452
rect 19156 29300 19208 29306
rect 19156 29242 19208 29248
rect 19168 29034 19196 29242
rect 19352 29209 19380 29582
rect 19708 29572 19760 29578
rect 19708 29514 19760 29520
rect 19338 29200 19394 29209
rect 19248 29164 19300 29170
rect 19720 29170 19748 29514
rect 19892 29504 19944 29510
rect 19892 29446 19944 29452
rect 19904 29170 19932 29446
rect 19338 29135 19340 29144
rect 19248 29106 19300 29112
rect 19392 29135 19394 29144
rect 19524 29164 19576 29170
rect 19340 29106 19392 29112
rect 19524 29106 19576 29112
rect 19708 29164 19760 29170
rect 19708 29106 19760 29112
rect 19892 29164 19944 29170
rect 19892 29106 19944 29112
rect 19156 29028 19208 29034
rect 19156 28970 19208 28976
rect 19260 27606 19288 29106
rect 19536 28218 19564 29106
rect 19720 28762 19748 29106
rect 19708 28756 19760 28762
rect 19708 28698 19760 28704
rect 19524 28212 19576 28218
rect 19524 28154 19576 28160
rect 19996 28098 20024 29718
rect 20180 28626 20208 30194
rect 20260 30048 20312 30054
rect 20260 29990 20312 29996
rect 20076 28620 20128 28626
rect 20076 28562 20128 28568
rect 20168 28620 20220 28626
rect 20168 28562 20220 28568
rect 20088 28218 20116 28562
rect 20272 28558 20300 29990
rect 20364 29782 20392 30194
rect 20732 30190 20760 32830
rect 20720 30184 20772 30190
rect 20720 30126 20772 30132
rect 20536 30048 20588 30054
rect 20536 29990 20588 29996
rect 20352 29776 20404 29782
rect 20352 29718 20404 29724
rect 20444 29640 20496 29646
rect 20444 29582 20496 29588
rect 20352 28960 20404 28966
rect 20352 28902 20404 28908
rect 20260 28552 20312 28558
rect 20260 28494 20312 28500
rect 20076 28212 20128 28218
rect 20076 28154 20128 28160
rect 19996 28070 20208 28098
rect 20364 28082 20392 28902
rect 20456 28762 20484 29582
rect 20548 28762 20576 29990
rect 20732 29646 20760 30126
rect 20824 29646 20852 32932
rect 21376 32910 21404 33526
rect 22296 33402 22324 33866
rect 22296 33374 22416 33402
rect 22052 33212 22360 33221
rect 22052 33210 22058 33212
rect 22114 33210 22138 33212
rect 22194 33210 22218 33212
rect 22274 33210 22298 33212
rect 22354 33210 22360 33212
rect 22114 33158 22116 33210
rect 22296 33158 22298 33210
rect 22052 33156 22058 33158
rect 22114 33156 22138 33158
rect 22194 33156 22218 33158
rect 22274 33156 22298 33158
rect 22354 33156 22360 33158
rect 22052 33147 22360 33156
rect 22388 33114 22416 33374
rect 22376 33108 22428 33114
rect 22376 33050 22428 33056
rect 22480 32910 22508 34614
rect 22572 33114 22600 35022
rect 22664 34542 22692 35430
rect 22744 34944 22796 34950
rect 22744 34886 22796 34892
rect 22652 34536 22704 34542
rect 22652 34478 22704 34484
rect 22664 33810 22692 34478
rect 22756 33930 22784 34886
rect 23020 34536 23072 34542
rect 23020 34478 23072 34484
rect 22744 33924 22796 33930
rect 22744 33866 22796 33872
rect 22664 33782 22784 33810
rect 22560 33108 22612 33114
rect 22560 33050 22612 33056
rect 21364 32904 21416 32910
rect 21364 32846 21416 32852
rect 22468 32904 22520 32910
rect 22468 32846 22520 32852
rect 22756 32842 22784 33782
rect 23032 33658 23060 34478
rect 23020 33652 23072 33658
rect 23020 33594 23072 33600
rect 22836 33312 22888 33318
rect 22836 33254 22888 33260
rect 22848 32978 22876 33254
rect 22836 32972 22888 32978
rect 22836 32914 22888 32920
rect 22744 32836 22796 32842
rect 22744 32778 22796 32784
rect 21088 32360 21140 32366
rect 21088 32302 21140 32308
rect 20996 31680 21048 31686
rect 20996 31622 21048 31628
rect 21008 31414 21036 31622
rect 21100 31482 21128 32302
rect 21456 32292 21508 32298
rect 21456 32234 21508 32240
rect 21180 32020 21232 32026
rect 21180 31962 21232 31968
rect 21192 31754 21220 31962
rect 21468 31958 21496 32234
rect 22468 32224 22520 32230
rect 22468 32166 22520 32172
rect 22052 32124 22360 32133
rect 22052 32122 22058 32124
rect 22114 32122 22138 32124
rect 22194 32122 22218 32124
rect 22274 32122 22298 32124
rect 22354 32122 22360 32124
rect 22114 32070 22116 32122
rect 22296 32070 22298 32122
rect 22052 32068 22058 32070
rect 22114 32068 22138 32070
rect 22194 32068 22218 32070
rect 22274 32068 22298 32070
rect 22354 32068 22360 32070
rect 22052 32059 22360 32068
rect 22100 32020 22152 32026
rect 22100 31962 22152 31968
rect 21456 31952 21508 31958
rect 21456 31894 21508 31900
rect 21192 31726 21312 31754
rect 21088 31476 21140 31482
rect 21088 31418 21140 31424
rect 20996 31408 21048 31414
rect 20996 31350 21048 31356
rect 21100 30734 21128 31418
rect 21088 30728 21140 30734
rect 21088 30670 21140 30676
rect 20996 30252 21048 30258
rect 20996 30194 21048 30200
rect 20628 29640 20680 29646
rect 20628 29582 20680 29588
rect 20720 29640 20772 29646
rect 20720 29582 20772 29588
rect 20812 29640 20864 29646
rect 20812 29582 20864 29588
rect 20444 28756 20496 28762
rect 20444 28698 20496 28704
rect 20536 28756 20588 28762
rect 20536 28698 20588 28704
rect 20640 28694 20668 29582
rect 21008 29306 21036 30194
rect 21284 30122 21312 31726
rect 21824 31748 21876 31754
rect 21824 31690 21876 31696
rect 21836 31346 21864 31690
rect 22112 31414 22140 31962
rect 22480 31754 22508 32166
rect 22756 31754 22784 32778
rect 22848 32434 22876 32914
rect 22836 32428 22888 32434
rect 22836 32370 22888 32376
rect 22928 32428 22980 32434
rect 22928 32370 22980 32376
rect 22940 32026 22968 32370
rect 23032 32230 23060 33594
rect 23020 32224 23072 32230
rect 23020 32166 23072 32172
rect 22928 32020 22980 32026
rect 22928 31962 22980 31968
rect 22480 31748 22612 31754
rect 22480 31726 22560 31748
rect 22756 31726 22876 31754
rect 22560 31690 22612 31696
rect 22652 31680 22704 31686
rect 22652 31622 22704 31628
rect 22100 31408 22152 31414
rect 22100 31350 22152 31356
rect 21824 31340 21876 31346
rect 21824 31282 21876 31288
rect 21836 30870 21864 31282
rect 22052 31036 22360 31045
rect 22052 31034 22058 31036
rect 22114 31034 22138 31036
rect 22194 31034 22218 31036
rect 22274 31034 22298 31036
rect 22354 31034 22360 31036
rect 22114 30982 22116 31034
rect 22296 30982 22298 31034
rect 22052 30980 22058 30982
rect 22114 30980 22138 30982
rect 22194 30980 22218 30982
rect 22274 30980 22298 30982
rect 22354 30980 22360 30982
rect 22052 30971 22360 30980
rect 22664 30938 22692 31622
rect 22652 30932 22704 30938
rect 22652 30874 22704 30880
rect 21548 30864 21600 30870
rect 21548 30806 21600 30812
rect 21824 30864 21876 30870
rect 21824 30806 21876 30812
rect 22008 30864 22060 30870
rect 22008 30806 22060 30812
rect 21272 30116 21324 30122
rect 21272 30058 21324 30064
rect 21284 29646 21312 30058
rect 21272 29640 21324 29646
rect 21272 29582 21324 29588
rect 21180 29504 21232 29510
rect 21180 29446 21232 29452
rect 20996 29300 21048 29306
rect 20996 29242 21048 29248
rect 20628 28688 20680 28694
rect 20628 28630 20680 28636
rect 21008 28626 21036 29242
rect 21192 29170 21220 29446
rect 21272 29232 21324 29238
rect 21272 29174 21324 29180
rect 21180 29164 21232 29170
rect 21180 29106 21232 29112
rect 20996 28620 21048 28626
rect 20996 28562 21048 28568
rect 19800 27872 19852 27878
rect 19800 27814 19852 27820
rect 19812 27606 19840 27814
rect 19248 27600 19300 27606
rect 19248 27542 19300 27548
rect 19800 27600 19852 27606
rect 19800 27542 19852 27548
rect 19064 27328 19116 27334
rect 19064 27270 19116 27276
rect 19798 27160 19854 27169
rect 19798 27095 19800 27104
rect 19852 27095 19854 27104
rect 19800 27066 19852 27072
rect 18788 26988 18840 26994
rect 18788 26930 18840 26936
rect 18800 25362 18828 26930
rect 19616 26920 19668 26926
rect 19616 26862 19668 26868
rect 19628 26518 19656 26862
rect 19708 26784 19760 26790
rect 19708 26726 19760 26732
rect 19720 26586 19748 26726
rect 19708 26580 19760 26586
rect 19708 26522 19760 26528
rect 19616 26512 19668 26518
rect 19616 26454 19668 26460
rect 19432 26376 19484 26382
rect 19484 26336 19564 26364
rect 19432 26318 19484 26324
rect 19340 25900 19392 25906
rect 19340 25842 19392 25848
rect 18788 25356 18840 25362
rect 18788 25298 18840 25304
rect 19156 24336 19208 24342
rect 19156 24278 19208 24284
rect 18696 24268 18748 24274
rect 18696 24210 18748 24216
rect 18328 23860 18380 23866
rect 18328 23802 18380 23808
rect 18156 23718 18276 23746
rect 17684 23520 17736 23526
rect 17684 23462 17736 23468
rect 17408 23112 17460 23118
rect 17408 23054 17460 23060
rect 17420 22642 17448 23054
rect 17408 22636 17460 22642
rect 17408 22578 17460 22584
rect 17132 22568 17184 22574
rect 17132 22510 17184 22516
rect 16764 21888 16816 21894
rect 16764 21830 16816 21836
rect 16776 21690 16804 21830
rect 16764 21684 16816 21690
rect 16764 21626 16816 21632
rect 16672 21548 16724 21554
rect 16672 21490 16724 21496
rect 16488 21344 16540 21350
rect 16488 21286 16540 21292
rect 16500 20942 16528 21286
rect 16488 20936 16540 20942
rect 16488 20878 16540 20884
rect 16684 20874 16712 21490
rect 16948 21480 17000 21486
rect 16948 21422 17000 21428
rect 16960 20942 16988 21422
rect 16948 20936 17000 20942
rect 16948 20878 17000 20884
rect 16672 20868 16724 20874
rect 16672 20810 16724 20816
rect 16396 20596 16448 20602
rect 16396 20538 16448 20544
rect 15292 20052 15344 20058
rect 15292 19994 15344 20000
rect 15660 20052 15712 20058
rect 15660 19994 15712 20000
rect 16408 19854 16436 20538
rect 17144 20466 17172 22510
rect 17500 22432 17552 22438
rect 17500 22374 17552 22380
rect 17408 22024 17460 22030
rect 17408 21966 17460 21972
rect 17316 21888 17368 21894
rect 17316 21830 17368 21836
rect 17328 21690 17356 21830
rect 17420 21690 17448 21966
rect 17316 21684 17368 21690
rect 17316 21626 17368 21632
rect 17408 21684 17460 21690
rect 17408 21626 17460 21632
rect 17512 21554 17540 22374
rect 17696 22030 17724 23462
rect 18156 23254 18184 23718
rect 18236 23520 18288 23526
rect 18236 23462 18288 23468
rect 18144 23248 18196 23254
rect 18144 23190 18196 23196
rect 18248 23186 18276 23462
rect 18236 23180 18288 23186
rect 18236 23122 18288 23128
rect 19168 23118 19196 24278
rect 19064 23112 19116 23118
rect 19064 23054 19116 23060
rect 19156 23112 19208 23118
rect 19156 23054 19208 23060
rect 18236 22976 18288 22982
rect 18236 22918 18288 22924
rect 17831 22876 18139 22885
rect 17831 22874 17837 22876
rect 17893 22874 17917 22876
rect 17973 22874 17997 22876
rect 18053 22874 18077 22876
rect 18133 22874 18139 22876
rect 17893 22822 17895 22874
rect 18075 22822 18077 22874
rect 17831 22820 17837 22822
rect 17893 22820 17917 22822
rect 17973 22820 17997 22822
rect 18053 22820 18077 22822
rect 18133 22820 18139 22822
rect 17831 22811 18139 22820
rect 18248 22642 18276 22918
rect 18236 22636 18288 22642
rect 18236 22578 18288 22584
rect 17960 22432 18012 22438
rect 17960 22374 18012 22380
rect 17972 22030 18000 22374
rect 19076 22094 19104 23054
rect 19076 22066 19288 22094
rect 17684 22024 17736 22030
rect 17684 21966 17736 21972
rect 17960 22024 18012 22030
rect 17960 21966 18012 21972
rect 18420 22024 18472 22030
rect 18420 21966 18472 21972
rect 17500 21548 17552 21554
rect 17500 21490 17552 21496
rect 17512 21078 17540 21490
rect 17500 21072 17552 21078
rect 17500 21014 17552 21020
rect 17696 20942 17724 21966
rect 17831 21788 18139 21797
rect 17831 21786 17837 21788
rect 17893 21786 17917 21788
rect 17973 21786 17997 21788
rect 18053 21786 18077 21788
rect 18133 21786 18139 21788
rect 17893 21734 17895 21786
rect 18075 21734 18077 21786
rect 17831 21732 17837 21734
rect 17893 21732 17917 21734
rect 17973 21732 17997 21734
rect 18053 21732 18077 21734
rect 18133 21732 18139 21734
rect 17831 21723 18139 21732
rect 18432 21690 18460 21966
rect 19260 21894 19288 22066
rect 18788 21888 18840 21894
rect 18788 21830 18840 21836
rect 19248 21888 19300 21894
rect 19248 21830 19300 21836
rect 18420 21684 18472 21690
rect 18420 21626 18472 21632
rect 18432 21418 18460 21626
rect 18420 21412 18472 21418
rect 18420 21354 18472 21360
rect 18696 21072 18748 21078
rect 18696 21014 18748 21020
rect 17684 20936 17736 20942
rect 17684 20878 17736 20884
rect 17696 20482 17724 20878
rect 17831 20700 18139 20709
rect 17831 20698 17837 20700
rect 17893 20698 17917 20700
rect 17973 20698 17997 20700
rect 18053 20698 18077 20700
rect 18133 20698 18139 20700
rect 17893 20646 17895 20698
rect 18075 20646 18077 20698
rect 17831 20644 17837 20646
rect 17893 20644 17917 20646
rect 17973 20644 17997 20646
rect 18053 20644 18077 20646
rect 18133 20644 18139 20646
rect 17831 20635 18139 20644
rect 17132 20460 17184 20466
rect 17696 20454 17816 20482
rect 17132 20402 17184 20408
rect 17144 19922 17172 20402
rect 17224 20392 17276 20398
rect 17224 20334 17276 20340
rect 17236 20058 17264 20334
rect 17788 20262 17816 20454
rect 17776 20256 17828 20262
rect 17776 20198 17828 20204
rect 17224 20052 17276 20058
rect 17224 19994 17276 20000
rect 17132 19916 17184 19922
rect 17132 19858 17184 19864
rect 17788 19854 17816 20198
rect 15016 19848 15068 19854
rect 15016 19790 15068 19796
rect 16396 19848 16448 19854
rect 16396 19790 16448 19796
rect 17776 19848 17828 19854
rect 17776 19790 17828 19796
rect 16408 19514 16436 19790
rect 18420 19780 18472 19786
rect 18420 19722 18472 19728
rect 17831 19612 18139 19621
rect 17831 19610 17837 19612
rect 17893 19610 17917 19612
rect 17973 19610 17997 19612
rect 18053 19610 18077 19612
rect 18133 19610 18139 19612
rect 17893 19558 17895 19610
rect 18075 19558 18077 19610
rect 17831 19556 17837 19558
rect 17893 19556 17917 19558
rect 17973 19556 17997 19558
rect 18053 19556 18077 19558
rect 18133 19556 18139 19558
rect 17831 19547 18139 19556
rect 18432 19514 18460 19722
rect 16396 19508 16448 19514
rect 16396 19450 16448 19456
rect 18420 19508 18472 19514
rect 18420 19450 18472 19456
rect 18708 19378 18736 21014
rect 18800 20874 18828 21830
rect 18788 20868 18840 20874
rect 18788 20810 18840 20816
rect 18800 19378 18828 20810
rect 18880 20800 18932 20806
rect 18880 20742 18932 20748
rect 18892 19514 18920 20742
rect 19352 20534 19380 25842
rect 19536 25770 19564 26336
rect 19524 25764 19576 25770
rect 19524 25706 19576 25712
rect 19536 25362 19564 25706
rect 19524 25356 19576 25362
rect 19524 25298 19576 25304
rect 19628 25294 19656 26454
rect 19708 26308 19760 26314
rect 19708 26250 19760 26256
rect 19720 25498 19748 26250
rect 19800 26240 19852 26246
rect 19800 26182 19852 26188
rect 19812 25906 19840 26182
rect 19984 25968 20036 25974
rect 19984 25910 20036 25916
rect 19800 25900 19852 25906
rect 19800 25842 19852 25848
rect 19708 25492 19760 25498
rect 19708 25434 19760 25440
rect 19432 25288 19484 25294
rect 19432 25230 19484 25236
rect 19616 25288 19668 25294
rect 19616 25230 19668 25236
rect 19444 24886 19472 25230
rect 19524 25220 19576 25226
rect 19524 25162 19576 25168
rect 19536 24954 19564 25162
rect 19524 24948 19576 24954
rect 19524 24890 19576 24896
rect 19432 24880 19484 24886
rect 19432 24822 19484 24828
rect 19444 24274 19472 24822
rect 19996 24818 20024 25910
rect 20076 25696 20128 25702
rect 20076 25638 20128 25644
rect 20088 25498 20116 25638
rect 20076 25492 20128 25498
rect 20076 25434 20128 25440
rect 20180 25294 20208 28070
rect 20352 28076 20404 28082
rect 20352 28018 20404 28024
rect 21088 27872 21140 27878
rect 21088 27814 21140 27820
rect 20720 27600 20772 27606
rect 20720 27542 20772 27548
rect 20732 26314 20760 27542
rect 20904 27328 20956 27334
rect 20904 27270 20956 27276
rect 20996 27328 21048 27334
rect 20996 27270 21048 27276
rect 20916 27130 20944 27270
rect 20904 27124 20956 27130
rect 20904 27066 20956 27072
rect 21008 26314 21036 27270
rect 21100 26586 21128 27814
rect 21284 27674 21312 29174
rect 21560 28994 21588 30806
rect 21732 30320 21784 30326
rect 21732 30262 21784 30268
rect 21640 30252 21692 30258
rect 21640 30194 21692 30200
rect 21652 29850 21680 30194
rect 21640 29844 21692 29850
rect 21640 29786 21692 29792
rect 21744 29782 21772 30262
rect 22020 30258 22048 30806
rect 22848 30734 22876 31726
rect 23124 30938 23152 39374
rect 26272 39196 26580 39205
rect 26272 39194 26278 39196
rect 26334 39194 26358 39196
rect 26414 39194 26438 39196
rect 26494 39194 26518 39196
rect 26574 39194 26580 39196
rect 26334 39142 26336 39194
rect 26516 39142 26518 39194
rect 26272 39140 26278 39142
rect 26334 39140 26358 39142
rect 26414 39140 26438 39142
rect 26494 39140 26518 39142
rect 26574 39140 26580 39142
rect 26272 39131 26580 39140
rect 23204 38888 23256 38894
rect 23204 38830 23256 38836
rect 23216 36786 23244 38830
rect 23940 38752 23992 38758
rect 23940 38694 23992 38700
rect 23952 38418 23980 38694
rect 23940 38412 23992 38418
rect 23940 38354 23992 38360
rect 26272 38108 26580 38117
rect 26272 38106 26278 38108
rect 26334 38106 26358 38108
rect 26414 38106 26438 38108
rect 26494 38106 26518 38108
rect 26574 38106 26580 38108
rect 26334 38054 26336 38106
rect 26516 38054 26518 38106
rect 26272 38052 26278 38054
rect 26334 38052 26358 38054
rect 26414 38052 26438 38054
rect 26494 38052 26518 38054
rect 26574 38052 26580 38054
rect 26272 38043 26580 38052
rect 23388 37800 23440 37806
rect 23388 37742 23440 37748
rect 23400 36922 23428 37742
rect 26272 37020 26580 37029
rect 26272 37018 26278 37020
rect 26334 37018 26358 37020
rect 26414 37018 26438 37020
rect 26494 37018 26518 37020
rect 26574 37018 26580 37020
rect 26334 36966 26336 37018
rect 26516 36966 26518 37018
rect 26272 36964 26278 36966
rect 26334 36964 26358 36966
rect 26414 36964 26438 36966
rect 26494 36964 26518 36966
rect 26574 36964 26580 36966
rect 26272 36955 26580 36964
rect 23388 36916 23440 36922
rect 23388 36858 23440 36864
rect 23204 36780 23256 36786
rect 23204 36722 23256 36728
rect 24492 36780 24544 36786
rect 24492 36722 24544 36728
rect 23216 36174 23244 36722
rect 23204 36168 23256 36174
rect 23204 36110 23256 36116
rect 23848 36100 23900 36106
rect 23848 36042 23900 36048
rect 23860 35834 23888 36042
rect 24504 35834 24532 36722
rect 26272 35932 26580 35941
rect 26272 35930 26278 35932
rect 26334 35930 26358 35932
rect 26414 35930 26438 35932
rect 26494 35930 26518 35932
rect 26574 35930 26580 35932
rect 26334 35878 26336 35930
rect 26516 35878 26518 35930
rect 26272 35876 26278 35878
rect 26334 35876 26358 35878
rect 26414 35876 26438 35878
rect 26494 35876 26518 35878
rect 26574 35876 26580 35878
rect 26272 35867 26580 35876
rect 23848 35828 23900 35834
rect 23848 35770 23900 35776
rect 24492 35828 24544 35834
rect 24492 35770 24544 35776
rect 24124 35692 24176 35698
rect 24124 35634 24176 35640
rect 24136 35290 24164 35634
rect 24124 35284 24176 35290
rect 24124 35226 24176 35232
rect 23572 35080 23624 35086
rect 23572 35022 23624 35028
rect 23204 34196 23256 34202
rect 23204 34138 23256 34144
rect 23216 32434 23244 34138
rect 23584 33930 23612 35022
rect 26272 34844 26580 34853
rect 26272 34842 26278 34844
rect 26334 34842 26358 34844
rect 26414 34842 26438 34844
rect 26494 34842 26518 34844
rect 26574 34842 26580 34844
rect 26334 34790 26336 34842
rect 26516 34790 26518 34842
rect 26272 34788 26278 34790
rect 26334 34788 26358 34790
rect 26414 34788 26438 34790
rect 26494 34788 26518 34790
rect 26574 34788 26580 34790
rect 26272 34779 26580 34788
rect 24124 34740 24176 34746
rect 24124 34682 24176 34688
rect 24032 33992 24084 33998
rect 24032 33934 24084 33940
rect 23572 33924 23624 33930
rect 23572 33866 23624 33872
rect 23296 33312 23348 33318
rect 23296 33254 23348 33260
rect 23308 32978 23336 33254
rect 23296 32972 23348 32978
rect 23296 32914 23348 32920
rect 23480 32768 23532 32774
rect 23480 32710 23532 32716
rect 23388 32496 23440 32502
rect 23388 32438 23440 32444
rect 23204 32428 23256 32434
rect 23204 32370 23256 32376
rect 23204 32292 23256 32298
rect 23204 32234 23256 32240
rect 23216 31822 23244 32234
rect 23296 32224 23348 32230
rect 23296 32166 23348 32172
rect 23308 31822 23336 32166
rect 23400 32026 23428 32438
rect 23388 32020 23440 32026
rect 23388 31962 23440 31968
rect 23204 31816 23256 31822
rect 23204 31758 23256 31764
rect 23296 31816 23348 31822
rect 23296 31758 23348 31764
rect 23112 30932 23164 30938
rect 23112 30874 23164 30880
rect 23216 30734 23244 31758
rect 23492 30802 23520 32710
rect 23480 30796 23532 30802
rect 23480 30738 23532 30744
rect 22836 30728 22888 30734
rect 22836 30670 22888 30676
rect 23204 30728 23256 30734
rect 23204 30670 23256 30676
rect 23216 30326 23244 30670
rect 23584 30410 23612 33866
rect 23848 33856 23900 33862
rect 23848 33798 23900 33804
rect 23940 33856 23992 33862
rect 23940 33798 23992 33804
rect 23860 32910 23888 33798
rect 23952 33658 23980 33798
rect 23940 33652 23992 33658
rect 23940 33594 23992 33600
rect 24044 33522 24072 33934
rect 24032 33516 24084 33522
rect 24032 33458 24084 33464
rect 23848 32904 23900 32910
rect 23848 32846 23900 32852
rect 23860 32570 23888 32846
rect 24044 32570 24072 33458
rect 23664 32564 23716 32570
rect 23664 32506 23716 32512
rect 23848 32564 23900 32570
rect 23848 32506 23900 32512
rect 24032 32564 24084 32570
rect 24032 32506 24084 32512
rect 23676 32026 23704 32506
rect 23940 32360 23992 32366
rect 23940 32302 23992 32308
rect 23664 32020 23716 32026
rect 23664 31962 23716 31968
rect 23676 31482 23704 31962
rect 23756 31680 23808 31686
rect 23756 31622 23808 31628
rect 23848 31680 23900 31686
rect 23848 31622 23900 31628
rect 23664 31476 23716 31482
rect 23664 31418 23716 31424
rect 23664 31340 23716 31346
rect 23664 31282 23716 31288
rect 23676 30938 23704 31282
rect 23768 31278 23796 31622
rect 23860 31482 23888 31622
rect 23952 31482 23980 32302
rect 24044 32026 24072 32506
rect 24032 32020 24084 32026
rect 24032 31962 24084 31968
rect 24136 31822 24164 34682
rect 24492 34604 24544 34610
rect 24492 34546 24544 34552
rect 24308 33856 24360 33862
rect 24308 33798 24360 33804
rect 24320 33522 24348 33798
rect 24504 33658 24532 34546
rect 24768 34536 24820 34542
rect 24768 34478 24820 34484
rect 24780 33658 24808 34478
rect 24860 34400 24912 34406
rect 24860 34342 24912 34348
rect 24872 34066 24900 34342
rect 24860 34060 24912 34066
rect 24860 34002 24912 34008
rect 26272 33756 26580 33765
rect 26272 33754 26278 33756
rect 26334 33754 26358 33756
rect 26414 33754 26438 33756
rect 26494 33754 26518 33756
rect 26574 33754 26580 33756
rect 26334 33702 26336 33754
rect 26516 33702 26518 33754
rect 26272 33700 26278 33702
rect 26334 33700 26358 33702
rect 26414 33700 26438 33702
rect 26494 33700 26518 33702
rect 26574 33700 26580 33702
rect 26272 33691 26580 33700
rect 24492 33652 24544 33658
rect 24492 33594 24544 33600
rect 24768 33652 24820 33658
rect 24768 33594 24820 33600
rect 24216 33516 24268 33522
rect 24216 33458 24268 33464
rect 24308 33516 24360 33522
rect 24308 33458 24360 33464
rect 24228 33114 24256 33458
rect 24216 33108 24268 33114
rect 24216 33050 24268 33056
rect 25320 32904 25372 32910
rect 25320 32846 25372 32852
rect 24400 32768 24452 32774
rect 24400 32710 24452 32716
rect 24412 32570 24440 32710
rect 25332 32570 25360 32846
rect 25504 32836 25556 32842
rect 25504 32778 25556 32784
rect 25516 32570 25544 32778
rect 26272 32668 26580 32677
rect 26272 32666 26278 32668
rect 26334 32666 26358 32668
rect 26414 32666 26438 32668
rect 26494 32666 26518 32668
rect 26574 32666 26580 32668
rect 26334 32614 26336 32666
rect 26516 32614 26518 32666
rect 26272 32612 26278 32614
rect 26334 32612 26358 32614
rect 26414 32612 26438 32614
rect 26494 32612 26518 32614
rect 26574 32612 26580 32614
rect 26272 32603 26580 32612
rect 24400 32564 24452 32570
rect 24400 32506 24452 32512
rect 24492 32564 24544 32570
rect 24492 32506 24544 32512
rect 25320 32564 25372 32570
rect 25320 32506 25372 32512
rect 25504 32564 25556 32570
rect 25504 32506 25556 32512
rect 24308 32020 24360 32026
rect 24308 31962 24360 31968
rect 24124 31816 24176 31822
rect 24124 31758 24176 31764
rect 24136 31482 24164 31758
rect 24320 31482 24348 31962
rect 24504 31822 24532 32506
rect 25780 32224 25832 32230
rect 25780 32166 25832 32172
rect 25792 32026 25820 32166
rect 24768 32020 24820 32026
rect 24768 31962 24820 31968
rect 25780 32020 25832 32026
rect 25780 31962 25832 31968
rect 24492 31816 24544 31822
rect 24492 31758 24544 31764
rect 24504 31482 24532 31758
rect 23848 31476 23900 31482
rect 23848 31418 23900 31424
rect 23940 31476 23992 31482
rect 23940 31418 23992 31424
rect 24124 31476 24176 31482
rect 24124 31418 24176 31424
rect 24308 31476 24360 31482
rect 24308 31418 24360 31424
rect 24492 31476 24544 31482
rect 24492 31418 24544 31424
rect 24320 31346 24348 31418
rect 24308 31340 24360 31346
rect 24308 31282 24360 31288
rect 24676 31340 24728 31346
rect 24676 31282 24728 31288
rect 23756 31272 23808 31278
rect 23756 31214 23808 31220
rect 23664 30932 23716 30938
rect 23664 30874 23716 30880
rect 23940 30592 23992 30598
rect 23940 30534 23992 30540
rect 23584 30382 23796 30410
rect 23204 30320 23256 30326
rect 23204 30262 23256 30268
rect 22008 30252 22060 30258
rect 21928 30212 22008 30240
rect 21824 30048 21876 30054
rect 21824 29990 21876 29996
rect 21732 29776 21784 29782
rect 21732 29718 21784 29724
rect 21836 29646 21864 29990
rect 21928 29646 21956 30212
rect 22008 30194 22060 30200
rect 22652 30048 22704 30054
rect 22652 29990 22704 29996
rect 23572 30048 23624 30054
rect 23572 29990 23624 29996
rect 22052 29948 22360 29957
rect 22052 29946 22058 29948
rect 22114 29946 22138 29948
rect 22194 29946 22218 29948
rect 22274 29946 22298 29948
rect 22354 29946 22360 29948
rect 22114 29894 22116 29946
rect 22296 29894 22298 29946
rect 22052 29892 22058 29894
rect 22114 29892 22138 29894
rect 22194 29892 22218 29894
rect 22274 29892 22298 29894
rect 22354 29892 22360 29894
rect 22052 29883 22360 29892
rect 21824 29640 21876 29646
rect 21824 29582 21876 29588
rect 21916 29640 21968 29646
rect 21916 29582 21968 29588
rect 21560 28966 21680 28994
rect 21364 28144 21416 28150
rect 21364 28086 21416 28092
rect 21548 28144 21600 28150
rect 21548 28086 21600 28092
rect 21272 27668 21324 27674
rect 21272 27610 21324 27616
rect 21180 27464 21232 27470
rect 21180 27406 21232 27412
rect 21192 27334 21220 27406
rect 21180 27328 21232 27334
rect 21180 27270 21232 27276
rect 21088 26580 21140 26586
rect 21088 26522 21140 26528
rect 21086 26480 21142 26489
rect 21086 26415 21142 26424
rect 20720 26308 20772 26314
rect 20720 26250 20772 26256
rect 20996 26308 21048 26314
rect 20996 26250 21048 26256
rect 20352 26240 20404 26246
rect 20352 26182 20404 26188
rect 20904 26240 20956 26246
rect 20904 26182 20956 26188
rect 20364 25906 20392 26182
rect 20352 25900 20404 25906
rect 20352 25842 20404 25848
rect 20916 25498 20944 26182
rect 20904 25492 20956 25498
rect 20904 25434 20956 25440
rect 20168 25288 20220 25294
rect 20168 25230 20220 25236
rect 20444 25220 20496 25226
rect 20444 25162 20496 25168
rect 20168 25152 20220 25158
rect 20168 25094 20220 25100
rect 19984 24812 20036 24818
rect 19984 24754 20036 24760
rect 19524 24608 19576 24614
rect 19524 24550 19576 24556
rect 19800 24608 19852 24614
rect 19800 24550 19852 24556
rect 19432 24268 19484 24274
rect 19432 24210 19484 24216
rect 19432 24064 19484 24070
rect 19432 24006 19484 24012
rect 19444 23322 19472 24006
rect 19536 23322 19564 24550
rect 19616 24268 19668 24274
rect 19616 24210 19668 24216
rect 19628 23866 19656 24210
rect 19812 23866 19840 24550
rect 19616 23860 19668 23866
rect 19616 23802 19668 23808
rect 19800 23860 19852 23866
rect 19800 23802 19852 23808
rect 20180 23730 20208 25094
rect 20260 24812 20312 24818
rect 20260 24754 20312 24760
rect 20272 24410 20300 24754
rect 20260 24404 20312 24410
rect 20260 24346 20312 24352
rect 19616 23724 19668 23730
rect 19616 23666 19668 23672
rect 20168 23724 20220 23730
rect 20168 23666 20220 23672
rect 19432 23316 19484 23322
rect 19432 23258 19484 23264
rect 19524 23316 19576 23322
rect 19524 23258 19576 23264
rect 19432 22500 19484 22506
rect 19432 22442 19484 22448
rect 19444 22030 19472 22442
rect 19432 22024 19484 22030
rect 19432 21966 19484 21972
rect 19432 21888 19484 21894
rect 19536 21842 19564 23258
rect 19628 23186 19656 23666
rect 19708 23520 19760 23526
rect 19708 23462 19760 23468
rect 19892 23520 19944 23526
rect 19892 23462 19944 23468
rect 19616 23180 19668 23186
rect 19616 23122 19668 23128
rect 19628 22642 19656 23122
rect 19720 22778 19748 23462
rect 19904 22982 19932 23462
rect 19892 22976 19944 22982
rect 19892 22918 19944 22924
rect 19708 22772 19760 22778
rect 19708 22714 19760 22720
rect 19904 22642 19932 22918
rect 19616 22636 19668 22642
rect 19616 22578 19668 22584
rect 19892 22636 19944 22642
rect 19892 22578 19944 22584
rect 20260 22636 20312 22642
rect 20260 22578 20312 22584
rect 20168 22568 20220 22574
rect 20168 22510 20220 22516
rect 19616 22432 19668 22438
rect 19616 22374 19668 22380
rect 19628 21962 19656 22374
rect 20076 22092 20128 22098
rect 20076 22034 20128 22040
rect 19616 21956 19668 21962
rect 19616 21898 19668 21904
rect 19484 21836 19564 21842
rect 19432 21830 19564 21836
rect 19892 21888 19944 21894
rect 19892 21830 19944 21836
rect 19444 21814 19564 21830
rect 19444 21690 19472 21814
rect 19432 21684 19484 21690
rect 19432 21626 19484 21632
rect 19904 21554 19932 21830
rect 20088 21554 20116 22034
rect 20180 22030 20208 22510
rect 20272 22030 20300 22578
rect 20352 22432 20404 22438
rect 20352 22374 20404 22380
rect 20364 22030 20392 22374
rect 20168 22024 20220 22030
rect 20168 21966 20220 21972
rect 20260 22024 20312 22030
rect 20260 21966 20312 21972
rect 20352 22024 20404 22030
rect 20352 21966 20404 21972
rect 20180 21690 20208 21966
rect 20168 21684 20220 21690
rect 20168 21626 20220 21632
rect 19892 21548 19944 21554
rect 19892 21490 19944 21496
rect 20076 21548 20128 21554
rect 20076 21490 20128 21496
rect 20352 21480 20404 21486
rect 20352 21422 20404 21428
rect 20168 21072 20220 21078
rect 20168 21014 20220 21020
rect 20076 20936 20128 20942
rect 20076 20878 20128 20884
rect 19340 20528 19392 20534
rect 19340 20470 19392 20476
rect 20088 20466 20116 20878
rect 20076 20460 20128 20466
rect 20076 20402 20128 20408
rect 19616 20052 19668 20058
rect 19616 19994 19668 20000
rect 18880 19508 18932 19514
rect 18880 19450 18932 19456
rect 19628 19378 19656 19994
rect 14924 19372 14976 19378
rect 14924 19314 14976 19320
rect 18696 19372 18748 19378
rect 18696 19314 18748 19320
rect 18788 19372 18840 19378
rect 18788 19314 18840 19320
rect 19616 19372 19668 19378
rect 19616 19314 19668 19320
rect 14096 19304 14148 19310
rect 14096 19246 14148 19252
rect 5170 19068 5478 19077
rect 5170 19066 5176 19068
rect 5232 19066 5256 19068
rect 5312 19066 5336 19068
rect 5392 19066 5416 19068
rect 5472 19066 5478 19068
rect 5232 19014 5234 19066
rect 5414 19014 5416 19066
rect 5170 19012 5176 19014
rect 5232 19012 5256 19014
rect 5312 19012 5336 19014
rect 5392 19012 5416 19014
rect 5472 19012 5478 19014
rect 5170 19003 5478 19012
rect 13611 19068 13919 19077
rect 13611 19066 13617 19068
rect 13673 19066 13697 19068
rect 13753 19066 13777 19068
rect 13833 19066 13857 19068
rect 13913 19066 13919 19068
rect 13673 19014 13675 19066
rect 13855 19014 13857 19066
rect 13611 19012 13617 19014
rect 13673 19012 13697 19014
rect 13753 19012 13777 19014
rect 13833 19012 13857 19014
rect 13913 19012 13919 19014
rect 13611 19003 13919 19012
rect 9390 18524 9698 18533
rect 9390 18522 9396 18524
rect 9452 18522 9476 18524
rect 9532 18522 9556 18524
rect 9612 18522 9636 18524
rect 9692 18522 9698 18524
rect 9452 18470 9454 18522
rect 9634 18470 9636 18522
rect 9390 18468 9396 18470
rect 9452 18468 9476 18470
rect 9532 18468 9556 18470
rect 9612 18468 9636 18470
rect 9692 18468 9698 18470
rect 9390 18459 9698 18468
rect 17831 18524 18139 18533
rect 17831 18522 17837 18524
rect 17893 18522 17917 18524
rect 17973 18522 17997 18524
rect 18053 18522 18077 18524
rect 18133 18522 18139 18524
rect 17893 18470 17895 18522
rect 18075 18470 18077 18522
rect 17831 18468 17837 18470
rect 17893 18468 17917 18470
rect 17973 18468 17997 18470
rect 18053 18468 18077 18470
rect 18133 18468 18139 18470
rect 17831 18459 18139 18468
rect 5170 17980 5478 17989
rect 5170 17978 5176 17980
rect 5232 17978 5256 17980
rect 5312 17978 5336 17980
rect 5392 17978 5416 17980
rect 5472 17978 5478 17980
rect 5232 17926 5234 17978
rect 5414 17926 5416 17978
rect 5170 17924 5176 17926
rect 5232 17924 5256 17926
rect 5312 17924 5336 17926
rect 5392 17924 5416 17926
rect 5472 17924 5478 17926
rect 5170 17915 5478 17924
rect 13611 17980 13919 17989
rect 13611 17978 13617 17980
rect 13673 17978 13697 17980
rect 13753 17978 13777 17980
rect 13833 17978 13857 17980
rect 13913 17978 13919 17980
rect 13673 17926 13675 17978
rect 13855 17926 13857 17978
rect 13611 17924 13617 17926
rect 13673 17924 13697 17926
rect 13753 17924 13777 17926
rect 13833 17924 13857 17926
rect 13913 17924 13919 17926
rect 13611 17915 13919 17924
rect 9390 17436 9698 17445
rect 9390 17434 9396 17436
rect 9452 17434 9476 17436
rect 9532 17434 9556 17436
rect 9612 17434 9636 17436
rect 9692 17434 9698 17436
rect 9452 17382 9454 17434
rect 9634 17382 9636 17434
rect 9390 17380 9396 17382
rect 9452 17380 9476 17382
rect 9532 17380 9556 17382
rect 9612 17380 9636 17382
rect 9692 17380 9698 17382
rect 9390 17371 9698 17380
rect 17831 17436 18139 17445
rect 17831 17434 17837 17436
rect 17893 17434 17917 17436
rect 17973 17434 17997 17436
rect 18053 17434 18077 17436
rect 18133 17434 18139 17436
rect 17893 17382 17895 17434
rect 18075 17382 18077 17434
rect 17831 17380 17837 17382
rect 17893 17380 17917 17382
rect 17973 17380 17997 17382
rect 18053 17380 18077 17382
rect 18133 17380 18139 17382
rect 17831 17371 18139 17380
rect 5170 16892 5478 16901
rect 5170 16890 5176 16892
rect 5232 16890 5256 16892
rect 5312 16890 5336 16892
rect 5392 16890 5416 16892
rect 5472 16890 5478 16892
rect 5232 16838 5234 16890
rect 5414 16838 5416 16890
rect 5170 16836 5176 16838
rect 5232 16836 5256 16838
rect 5312 16836 5336 16838
rect 5392 16836 5416 16838
rect 5472 16836 5478 16838
rect 5170 16827 5478 16836
rect 13611 16892 13919 16901
rect 13611 16890 13617 16892
rect 13673 16890 13697 16892
rect 13753 16890 13777 16892
rect 13833 16890 13857 16892
rect 13913 16890 13919 16892
rect 13673 16838 13675 16890
rect 13855 16838 13857 16890
rect 13611 16836 13617 16838
rect 13673 16836 13697 16838
rect 13753 16836 13777 16838
rect 13833 16836 13857 16838
rect 13913 16836 13919 16838
rect 13611 16827 13919 16836
rect 9390 16348 9698 16357
rect 9390 16346 9396 16348
rect 9452 16346 9476 16348
rect 9532 16346 9556 16348
rect 9612 16346 9636 16348
rect 9692 16346 9698 16348
rect 9452 16294 9454 16346
rect 9634 16294 9636 16346
rect 9390 16292 9396 16294
rect 9452 16292 9476 16294
rect 9532 16292 9556 16294
rect 9612 16292 9636 16294
rect 9692 16292 9698 16294
rect 9390 16283 9698 16292
rect 17831 16348 18139 16357
rect 17831 16346 17837 16348
rect 17893 16346 17917 16348
rect 17973 16346 17997 16348
rect 18053 16346 18077 16348
rect 18133 16346 18139 16348
rect 17893 16294 17895 16346
rect 18075 16294 18077 16346
rect 17831 16292 17837 16294
rect 17893 16292 17917 16294
rect 17973 16292 17997 16294
rect 18053 16292 18077 16294
rect 18133 16292 18139 16294
rect 17831 16283 18139 16292
rect 5170 15804 5478 15813
rect 5170 15802 5176 15804
rect 5232 15802 5256 15804
rect 5312 15802 5336 15804
rect 5392 15802 5416 15804
rect 5472 15802 5478 15804
rect 5232 15750 5234 15802
rect 5414 15750 5416 15802
rect 5170 15748 5176 15750
rect 5232 15748 5256 15750
rect 5312 15748 5336 15750
rect 5392 15748 5416 15750
rect 5472 15748 5478 15750
rect 5170 15739 5478 15748
rect 13611 15804 13919 15813
rect 13611 15802 13617 15804
rect 13673 15802 13697 15804
rect 13753 15802 13777 15804
rect 13833 15802 13857 15804
rect 13913 15802 13919 15804
rect 13673 15750 13675 15802
rect 13855 15750 13857 15802
rect 13611 15748 13617 15750
rect 13673 15748 13697 15750
rect 13753 15748 13777 15750
rect 13833 15748 13857 15750
rect 13913 15748 13919 15750
rect 13611 15739 13919 15748
rect 9390 15260 9698 15269
rect 9390 15258 9396 15260
rect 9452 15258 9476 15260
rect 9532 15258 9556 15260
rect 9612 15258 9636 15260
rect 9692 15258 9698 15260
rect 9452 15206 9454 15258
rect 9634 15206 9636 15258
rect 9390 15204 9396 15206
rect 9452 15204 9476 15206
rect 9532 15204 9556 15206
rect 9612 15204 9636 15206
rect 9692 15204 9698 15206
rect 9390 15195 9698 15204
rect 17831 15260 18139 15269
rect 17831 15258 17837 15260
rect 17893 15258 17917 15260
rect 17973 15258 17997 15260
rect 18053 15258 18077 15260
rect 18133 15258 18139 15260
rect 17893 15206 17895 15258
rect 18075 15206 18077 15258
rect 17831 15204 17837 15206
rect 17893 15204 17917 15206
rect 17973 15204 17997 15206
rect 18053 15204 18077 15206
rect 18133 15204 18139 15206
rect 17831 15195 18139 15204
rect 5170 14716 5478 14725
rect 5170 14714 5176 14716
rect 5232 14714 5256 14716
rect 5312 14714 5336 14716
rect 5392 14714 5416 14716
rect 5472 14714 5478 14716
rect 5232 14662 5234 14714
rect 5414 14662 5416 14714
rect 5170 14660 5176 14662
rect 5232 14660 5256 14662
rect 5312 14660 5336 14662
rect 5392 14660 5416 14662
rect 5472 14660 5478 14662
rect 5170 14651 5478 14660
rect 13611 14716 13919 14725
rect 13611 14714 13617 14716
rect 13673 14714 13697 14716
rect 13753 14714 13777 14716
rect 13833 14714 13857 14716
rect 13913 14714 13919 14716
rect 13673 14662 13675 14714
rect 13855 14662 13857 14714
rect 13611 14660 13617 14662
rect 13673 14660 13697 14662
rect 13753 14660 13777 14662
rect 13833 14660 13857 14662
rect 13913 14660 13919 14662
rect 13611 14651 13919 14660
rect 1584 14612 1636 14618
rect 1584 14554 1636 14560
rect 940 14408 992 14414
rect 938 14376 940 14385
rect 992 14376 994 14385
rect 938 14311 994 14320
rect 9390 14172 9698 14181
rect 9390 14170 9396 14172
rect 9452 14170 9476 14172
rect 9532 14170 9556 14172
rect 9612 14170 9636 14172
rect 9692 14170 9698 14172
rect 9452 14118 9454 14170
rect 9634 14118 9636 14170
rect 9390 14116 9396 14118
rect 9452 14116 9476 14118
rect 9532 14116 9556 14118
rect 9612 14116 9636 14118
rect 9692 14116 9698 14118
rect 9390 14107 9698 14116
rect 17831 14172 18139 14181
rect 17831 14170 17837 14172
rect 17893 14170 17917 14172
rect 17973 14170 17997 14172
rect 18053 14170 18077 14172
rect 18133 14170 18139 14172
rect 17893 14118 17895 14170
rect 18075 14118 18077 14170
rect 17831 14116 17837 14118
rect 17893 14116 17917 14118
rect 17973 14116 17997 14118
rect 18053 14116 18077 14118
rect 18133 14116 18139 14118
rect 17831 14107 18139 14116
rect 5170 13628 5478 13637
rect 5170 13626 5176 13628
rect 5232 13626 5256 13628
rect 5312 13626 5336 13628
rect 5392 13626 5416 13628
rect 5472 13626 5478 13628
rect 5232 13574 5234 13626
rect 5414 13574 5416 13626
rect 5170 13572 5176 13574
rect 5232 13572 5256 13574
rect 5312 13572 5336 13574
rect 5392 13572 5416 13574
rect 5472 13572 5478 13574
rect 5170 13563 5478 13572
rect 13611 13628 13919 13637
rect 13611 13626 13617 13628
rect 13673 13626 13697 13628
rect 13753 13626 13777 13628
rect 13833 13626 13857 13628
rect 13913 13626 13919 13628
rect 13673 13574 13675 13626
rect 13855 13574 13857 13626
rect 13611 13572 13617 13574
rect 13673 13572 13697 13574
rect 13753 13572 13777 13574
rect 13833 13572 13857 13574
rect 13913 13572 13919 13574
rect 13611 13563 13919 13572
rect 9390 13084 9698 13093
rect 9390 13082 9396 13084
rect 9452 13082 9476 13084
rect 9532 13082 9556 13084
rect 9612 13082 9636 13084
rect 9692 13082 9698 13084
rect 9452 13030 9454 13082
rect 9634 13030 9636 13082
rect 9390 13028 9396 13030
rect 9452 13028 9476 13030
rect 9532 13028 9556 13030
rect 9612 13028 9636 13030
rect 9692 13028 9698 13030
rect 9390 13019 9698 13028
rect 17831 13084 18139 13093
rect 17831 13082 17837 13084
rect 17893 13082 17917 13084
rect 17973 13082 17997 13084
rect 18053 13082 18077 13084
rect 18133 13082 18139 13084
rect 17893 13030 17895 13082
rect 18075 13030 18077 13082
rect 17831 13028 17837 13030
rect 17893 13028 17917 13030
rect 17973 13028 17997 13030
rect 18053 13028 18077 13030
rect 18133 13028 18139 13030
rect 17831 13019 18139 13028
rect 5170 12540 5478 12549
rect 5170 12538 5176 12540
rect 5232 12538 5256 12540
rect 5312 12538 5336 12540
rect 5392 12538 5416 12540
rect 5472 12538 5478 12540
rect 5232 12486 5234 12538
rect 5414 12486 5416 12538
rect 5170 12484 5176 12486
rect 5232 12484 5256 12486
rect 5312 12484 5336 12486
rect 5392 12484 5416 12486
rect 5472 12484 5478 12486
rect 5170 12475 5478 12484
rect 13611 12540 13919 12549
rect 13611 12538 13617 12540
rect 13673 12538 13697 12540
rect 13753 12538 13777 12540
rect 13833 12538 13857 12540
rect 13913 12538 13919 12540
rect 13673 12486 13675 12538
rect 13855 12486 13857 12538
rect 13611 12484 13617 12486
rect 13673 12484 13697 12486
rect 13753 12484 13777 12486
rect 13833 12484 13857 12486
rect 13913 12484 13919 12486
rect 13611 12475 13919 12484
rect 20180 12434 20208 21014
rect 20364 20942 20392 21422
rect 20456 21146 20484 25162
rect 20720 25152 20772 25158
rect 20720 25094 20772 25100
rect 20812 25152 20864 25158
rect 20812 25094 20864 25100
rect 20732 24954 20760 25094
rect 20720 24948 20772 24954
rect 20720 24890 20772 24896
rect 20534 23216 20590 23225
rect 20534 23151 20590 23160
rect 20548 23118 20576 23151
rect 20536 23112 20588 23118
rect 20536 23054 20588 23060
rect 20824 22953 20852 25094
rect 21008 24410 21036 26250
rect 21100 25906 21128 26415
rect 21088 25900 21140 25906
rect 21088 25842 21140 25848
rect 21192 25294 21220 27270
rect 21284 26994 21312 27610
rect 21376 27062 21404 28086
rect 21456 27872 21508 27878
rect 21456 27814 21508 27820
rect 21468 27130 21496 27814
rect 21456 27124 21508 27130
rect 21456 27066 21508 27072
rect 21364 27056 21416 27062
rect 21364 26998 21416 27004
rect 21272 26988 21324 26994
rect 21272 26930 21324 26936
rect 21284 26042 21312 26930
rect 21376 26246 21404 26998
rect 21468 26450 21496 27066
rect 21560 26994 21588 28086
rect 21652 27470 21680 28966
rect 22052 28860 22360 28869
rect 22052 28858 22058 28860
rect 22114 28858 22138 28860
rect 22194 28858 22218 28860
rect 22274 28858 22298 28860
rect 22354 28858 22360 28860
rect 22114 28806 22116 28858
rect 22296 28806 22298 28858
rect 22052 28804 22058 28806
rect 22114 28804 22138 28806
rect 22194 28804 22218 28806
rect 22274 28804 22298 28806
rect 22354 28804 22360 28806
rect 22052 28795 22360 28804
rect 22664 28558 22692 29990
rect 23584 29646 23612 29990
rect 23572 29640 23624 29646
rect 23572 29582 23624 29588
rect 22744 29504 22796 29510
rect 22744 29446 22796 29452
rect 23296 29504 23348 29510
rect 23296 29446 23348 29452
rect 22756 28762 22784 29446
rect 23308 29306 23336 29446
rect 23296 29300 23348 29306
rect 23296 29242 23348 29248
rect 23768 29170 23796 30382
rect 23848 30252 23900 30258
rect 23848 30194 23900 30200
rect 23860 29850 23888 30194
rect 23848 29844 23900 29850
rect 23848 29786 23900 29792
rect 23952 29646 23980 30534
rect 24688 30394 24716 31282
rect 24780 31278 24808 31962
rect 26272 31580 26580 31589
rect 26272 31578 26278 31580
rect 26334 31578 26358 31580
rect 26414 31578 26438 31580
rect 26494 31578 26518 31580
rect 26574 31578 26580 31580
rect 26334 31526 26336 31578
rect 26516 31526 26518 31578
rect 26272 31524 26278 31526
rect 26334 31524 26358 31526
rect 26414 31524 26438 31526
rect 26494 31524 26518 31526
rect 26574 31524 26580 31526
rect 26272 31515 26580 31524
rect 24768 31272 24820 31278
rect 24768 31214 24820 31220
rect 25504 31136 25556 31142
rect 25504 31078 25556 31084
rect 25516 30938 25544 31078
rect 25504 30932 25556 30938
rect 25504 30874 25556 30880
rect 26272 30492 26580 30501
rect 26272 30490 26278 30492
rect 26334 30490 26358 30492
rect 26414 30490 26438 30492
rect 26494 30490 26518 30492
rect 26574 30490 26580 30492
rect 26334 30438 26336 30490
rect 26516 30438 26518 30490
rect 26272 30436 26278 30438
rect 26334 30436 26358 30438
rect 26414 30436 26438 30438
rect 26494 30436 26518 30438
rect 26574 30436 26580 30438
rect 26272 30427 26580 30436
rect 24676 30388 24728 30394
rect 24676 30330 24728 30336
rect 29012 29646 29040 41200
rect 30493 39740 30801 39749
rect 30493 39738 30499 39740
rect 30555 39738 30579 39740
rect 30635 39738 30659 39740
rect 30715 39738 30739 39740
rect 30795 39738 30801 39740
rect 30555 39686 30557 39738
rect 30737 39686 30739 39738
rect 30493 39684 30499 39686
rect 30555 39684 30579 39686
rect 30635 39684 30659 39686
rect 30715 39684 30739 39686
rect 30795 39684 30801 39686
rect 30493 39675 30801 39684
rect 35452 39506 35480 41200
rect 35440 39500 35492 39506
rect 35440 39442 35492 39448
rect 34713 39196 35021 39205
rect 34713 39194 34719 39196
rect 34775 39194 34799 39196
rect 34855 39194 34879 39196
rect 34935 39194 34959 39196
rect 35015 39194 35021 39196
rect 34775 39142 34777 39194
rect 34957 39142 34959 39194
rect 34713 39140 34719 39142
rect 34775 39140 34799 39142
rect 34855 39140 34879 39142
rect 34935 39140 34959 39142
rect 35015 39140 35021 39142
rect 34713 39131 35021 39140
rect 30493 38652 30801 38661
rect 30493 38650 30499 38652
rect 30555 38650 30579 38652
rect 30635 38650 30659 38652
rect 30715 38650 30739 38652
rect 30795 38650 30801 38652
rect 30555 38598 30557 38650
rect 30737 38598 30739 38650
rect 30493 38596 30499 38598
rect 30555 38596 30579 38598
rect 30635 38596 30659 38598
rect 30715 38596 30739 38598
rect 30795 38596 30801 38598
rect 30493 38587 30801 38596
rect 34713 38108 35021 38117
rect 34713 38106 34719 38108
rect 34775 38106 34799 38108
rect 34855 38106 34879 38108
rect 34935 38106 34959 38108
rect 35015 38106 35021 38108
rect 34775 38054 34777 38106
rect 34957 38054 34959 38106
rect 34713 38052 34719 38054
rect 34775 38052 34799 38054
rect 34855 38052 34879 38054
rect 34935 38052 34959 38054
rect 35015 38052 35021 38054
rect 34713 38043 35021 38052
rect 30493 37564 30801 37573
rect 30493 37562 30499 37564
rect 30555 37562 30579 37564
rect 30635 37562 30659 37564
rect 30715 37562 30739 37564
rect 30795 37562 30801 37564
rect 30555 37510 30557 37562
rect 30737 37510 30739 37562
rect 30493 37508 30499 37510
rect 30555 37508 30579 37510
rect 30635 37508 30659 37510
rect 30715 37508 30739 37510
rect 30795 37508 30801 37510
rect 30493 37499 30801 37508
rect 34713 37020 35021 37029
rect 34713 37018 34719 37020
rect 34775 37018 34799 37020
rect 34855 37018 34879 37020
rect 34935 37018 34959 37020
rect 35015 37018 35021 37020
rect 34775 36966 34777 37018
rect 34957 36966 34959 37018
rect 34713 36964 34719 36966
rect 34775 36964 34799 36966
rect 34855 36964 34879 36966
rect 34935 36964 34959 36966
rect 35015 36964 35021 36966
rect 34713 36955 35021 36964
rect 30493 36476 30801 36485
rect 30493 36474 30499 36476
rect 30555 36474 30579 36476
rect 30635 36474 30659 36476
rect 30715 36474 30739 36476
rect 30795 36474 30801 36476
rect 30555 36422 30557 36474
rect 30737 36422 30739 36474
rect 30493 36420 30499 36422
rect 30555 36420 30579 36422
rect 30635 36420 30659 36422
rect 30715 36420 30739 36422
rect 30795 36420 30801 36422
rect 30493 36411 30801 36420
rect 34713 35932 35021 35941
rect 34713 35930 34719 35932
rect 34775 35930 34799 35932
rect 34855 35930 34879 35932
rect 34935 35930 34959 35932
rect 35015 35930 35021 35932
rect 34775 35878 34777 35930
rect 34957 35878 34959 35930
rect 34713 35876 34719 35878
rect 34775 35876 34799 35878
rect 34855 35876 34879 35878
rect 34935 35876 34959 35878
rect 35015 35876 35021 35878
rect 34713 35867 35021 35876
rect 30493 35388 30801 35397
rect 30493 35386 30499 35388
rect 30555 35386 30579 35388
rect 30635 35386 30659 35388
rect 30715 35386 30739 35388
rect 30795 35386 30801 35388
rect 30555 35334 30557 35386
rect 30737 35334 30739 35386
rect 30493 35332 30499 35334
rect 30555 35332 30579 35334
rect 30635 35332 30659 35334
rect 30715 35332 30739 35334
rect 30795 35332 30801 35334
rect 30493 35323 30801 35332
rect 35164 34944 35216 34950
rect 35164 34886 35216 34892
rect 34713 34844 35021 34853
rect 34713 34842 34719 34844
rect 34775 34842 34799 34844
rect 34855 34842 34879 34844
rect 34935 34842 34959 34844
rect 35015 34842 35021 34844
rect 34775 34790 34777 34842
rect 34957 34790 34959 34842
rect 34713 34788 34719 34790
rect 34775 34788 34799 34790
rect 34855 34788 34879 34790
rect 34935 34788 34959 34790
rect 35015 34788 35021 34790
rect 34713 34779 35021 34788
rect 35176 34785 35204 34886
rect 35162 34776 35218 34785
rect 35162 34711 35218 34720
rect 30493 34300 30801 34309
rect 30493 34298 30499 34300
rect 30555 34298 30579 34300
rect 30635 34298 30659 34300
rect 30715 34298 30739 34300
rect 30795 34298 30801 34300
rect 30555 34246 30557 34298
rect 30737 34246 30739 34298
rect 30493 34244 30499 34246
rect 30555 34244 30579 34246
rect 30635 34244 30659 34246
rect 30715 34244 30739 34246
rect 30795 34244 30801 34246
rect 30493 34235 30801 34244
rect 34713 33756 35021 33765
rect 34713 33754 34719 33756
rect 34775 33754 34799 33756
rect 34855 33754 34879 33756
rect 34935 33754 34959 33756
rect 35015 33754 35021 33756
rect 34775 33702 34777 33754
rect 34957 33702 34959 33754
rect 34713 33700 34719 33702
rect 34775 33700 34799 33702
rect 34855 33700 34879 33702
rect 34935 33700 34959 33702
rect 35015 33700 35021 33702
rect 34713 33691 35021 33700
rect 30493 33212 30801 33221
rect 30493 33210 30499 33212
rect 30555 33210 30579 33212
rect 30635 33210 30659 33212
rect 30715 33210 30739 33212
rect 30795 33210 30801 33212
rect 30555 33158 30557 33210
rect 30737 33158 30739 33210
rect 30493 33156 30499 33158
rect 30555 33156 30579 33158
rect 30635 33156 30659 33158
rect 30715 33156 30739 33158
rect 30795 33156 30801 33158
rect 30493 33147 30801 33156
rect 34713 32668 35021 32677
rect 34713 32666 34719 32668
rect 34775 32666 34799 32668
rect 34855 32666 34879 32668
rect 34935 32666 34959 32668
rect 35015 32666 35021 32668
rect 34775 32614 34777 32666
rect 34957 32614 34959 32666
rect 34713 32612 34719 32614
rect 34775 32612 34799 32614
rect 34855 32612 34879 32614
rect 34935 32612 34959 32614
rect 35015 32612 35021 32614
rect 34713 32603 35021 32612
rect 30493 32124 30801 32133
rect 30493 32122 30499 32124
rect 30555 32122 30579 32124
rect 30635 32122 30659 32124
rect 30715 32122 30739 32124
rect 30795 32122 30801 32124
rect 30555 32070 30557 32122
rect 30737 32070 30739 32122
rect 30493 32068 30499 32070
rect 30555 32068 30579 32070
rect 30635 32068 30659 32070
rect 30715 32068 30739 32070
rect 30795 32068 30801 32070
rect 30493 32059 30801 32068
rect 34713 31580 35021 31589
rect 34713 31578 34719 31580
rect 34775 31578 34799 31580
rect 34855 31578 34879 31580
rect 34935 31578 34959 31580
rect 35015 31578 35021 31580
rect 34775 31526 34777 31578
rect 34957 31526 34959 31578
rect 34713 31524 34719 31526
rect 34775 31524 34799 31526
rect 34855 31524 34879 31526
rect 34935 31524 34959 31526
rect 35015 31524 35021 31526
rect 34713 31515 35021 31524
rect 30493 31036 30801 31045
rect 30493 31034 30499 31036
rect 30555 31034 30579 31036
rect 30635 31034 30659 31036
rect 30715 31034 30739 31036
rect 30795 31034 30801 31036
rect 30555 30982 30557 31034
rect 30737 30982 30739 31034
rect 30493 30980 30499 30982
rect 30555 30980 30579 30982
rect 30635 30980 30659 30982
rect 30715 30980 30739 30982
rect 30795 30980 30801 30982
rect 30493 30971 30801 30980
rect 34713 30492 35021 30501
rect 34713 30490 34719 30492
rect 34775 30490 34799 30492
rect 34855 30490 34879 30492
rect 34935 30490 34959 30492
rect 35015 30490 35021 30492
rect 34775 30438 34777 30490
rect 34957 30438 34959 30490
rect 34713 30436 34719 30438
rect 34775 30436 34799 30438
rect 34855 30436 34879 30438
rect 34935 30436 34959 30438
rect 35015 30436 35021 30438
rect 34713 30427 35021 30436
rect 30493 29948 30801 29957
rect 30493 29946 30499 29948
rect 30555 29946 30579 29948
rect 30635 29946 30659 29948
rect 30715 29946 30739 29948
rect 30795 29946 30801 29948
rect 30555 29894 30557 29946
rect 30737 29894 30739 29946
rect 30493 29892 30499 29894
rect 30555 29892 30579 29894
rect 30635 29892 30659 29894
rect 30715 29892 30739 29894
rect 30795 29892 30801 29894
rect 30493 29883 30801 29892
rect 23940 29640 23992 29646
rect 23940 29582 23992 29588
rect 24032 29640 24084 29646
rect 24032 29582 24084 29588
rect 29000 29640 29052 29646
rect 29000 29582 29052 29588
rect 24044 29306 24072 29582
rect 26272 29404 26580 29413
rect 26272 29402 26278 29404
rect 26334 29402 26358 29404
rect 26414 29402 26438 29404
rect 26494 29402 26518 29404
rect 26574 29402 26580 29404
rect 26334 29350 26336 29402
rect 26516 29350 26518 29402
rect 26272 29348 26278 29350
rect 26334 29348 26358 29350
rect 26414 29348 26438 29350
rect 26494 29348 26518 29350
rect 26574 29348 26580 29350
rect 26272 29339 26580 29348
rect 34713 29404 35021 29413
rect 34713 29402 34719 29404
rect 34775 29402 34799 29404
rect 34855 29402 34879 29404
rect 34935 29402 34959 29404
rect 35015 29402 35021 29404
rect 34775 29350 34777 29402
rect 34957 29350 34959 29402
rect 34713 29348 34719 29350
rect 34775 29348 34799 29350
rect 34855 29348 34879 29350
rect 34935 29348 34959 29350
rect 35015 29348 35021 29350
rect 34713 29339 35021 29348
rect 24032 29300 24084 29306
rect 24032 29242 24084 29248
rect 23756 29164 23808 29170
rect 23756 29106 23808 29112
rect 23940 29164 23992 29170
rect 23940 29106 23992 29112
rect 23296 28960 23348 28966
rect 23296 28902 23348 28908
rect 23308 28762 23336 28902
rect 22744 28756 22796 28762
rect 22744 28698 22796 28704
rect 23296 28756 23348 28762
rect 23296 28698 23348 28704
rect 22756 28626 22784 28698
rect 22744 28620 22796 28626
rect 22744 28562 22796 28568
rect 22652 28552 22704 28558
rect 22652 28494 22704 28500
rect 22284 28416 22336 28422
rect 22284 28358 22336 28364
rect 22560 28416 22612 28422
rect 22560 28358 22612 28364
rect 21916 28076 21968 28082
rect 21916 28018 21968 28024
rect 21732 27532 21784 27538
rect 21732 27474 21784 27480
rect 21640 27464 21692 27470
rect 21640 27406 21692 27412
rect 21652 27130 21680 27406
rect 21744 27169 21772 27474
rect 21928 27334 21956 28018
rect 22296 27878 22324 28358
rect 22572 28150 22600 28358
rect 22560 28144 22612 28150
rect 22560 28086 22612 28092
rect 22284 27872 22336 27878
rect 22284 27814 22336 27820
rect 22052 27772 22360 27781
rect 22052 27770 22058 27772
rect 22114 27770 22138 27772
rect 22194 27770 22218 27772
rect 22274 27770 22298 27772
rect 22354 27770 22360 27772
rect 22114 27718 22116 27770
rect 22296 27718 22298 27770
rect 22052 27716 22058 27718
rect 22114 27716 22138 27718
rect 22194 27716 22218 27718
rect 22274 27716 22298 27718
rect 22354 27716 22360 27718
rect 22052 27707 22360 27716
rect 21916 27328 21968 27334
rect 21916 27270 21968 27276
rect 21730 27160 21786 27169
rect 21640 27124 21692 27130
rect 21730 27095 21786 27104
rect 21640 27066 21692 27072
rect 22572 27010 22600 28086
rect 23848 27872 23900 27878
rect 23848 27814 23900 27820
rect 23020 27668 23072 27674
rect 23020 27610 23072 27616
rect 22744 27464 22796 27470
rect 22744 27406 22796 27412
rect 22652 27396 22704 27402
rect 22652 27338 22704 27344
rect 22664 27130 22692 27338
rect 22652 27124 22704 27130
rect 22652 27066 22704 27072
rect 21548 26988 21600 26994
rect 21548 26930 21600 26936
rect 21744 26982 22600 27010
rect 22756 26994 22784 27406
rect 22928 27328 22980 27334
rect 22928 27270 22980 27276
rect 22940 27130 22968 27270
rect 22928 27124 22980 27130
rect 22928 27066 22980 27072
rect 22744 26988 22796 26994
rect 21456 26444 21508 26450
rect 21456 26386 21508 26392
rect 21560 26382 21588 26930
rect 21640 26784 21692 26790
rect 21640 26726 21692 26732
rect 21652 26586 21680 26726
rect 21640 26580 21692 26586
rect 21640 26522 21692 26528
rect 21744 26382 21772 26982
rect 22744 26930 22796 26936
rect 22284 26852 22336 26858
rect 22336 26812 22416 26840
rect 22284 26794 22336 26800
rect 21824 26784 21876 26790
rect 21824 26726 21876 26732
rect 21548 26376 21600 26382
rect 21548 26318 21600 26324
rect 21732 26376 21784 26382
rect 21732 26318 21784 26324
rect 21364 26240 21416 26246
rect 21560 26234 21588 26318
rect 21364 26182 21416 26188
rect 21468 26206 21588 26234
rect 21272 26036 21324 26042
rect 21272 25978 21324 25984
rect 21364 26036 21416 26042
rect 21364 25978 21416 25984
rect 21376 25838 21404 25978
rect 21468 25974 21496 26206
rect 21456 25968 21508 25974
rect 21456 25910 21508 25916
rect 21364 25832 21416 25838
rect 21364 25774 21416 25780
rect 21272 25424 21324 25430
rect 21272 25366 21324 25372
rect 21180 25288 21232 25294
rect 21180 25230 21232 25236
rect 20996 24404 21048 24410
rect 20996 24346 21048 24352
rect 21284 24206 21312 25366
rect 21272 24200 21324 24206
rect 21272 24142 21324 24148
rect 21376 23118 21404 25774
rect 21468 24750 21496 25910
rect 21640 25900 21692 25906
rect 21640 25842 21692 25848
rect 21652 25294 21680 25842
rect 21744 25362 21772 26318
rect 21836 26314 21864 26726
rect 22052 26684 22360 26693
rect 22052 26682 22058 26684
rect 22114 26682 22138 26684
rect 22194 26682 22218 26684
rect 22274 26682 22298 26684
rect 22354 26682 22360 26684
rect 22114 26630 22116 26682
rect 22296 26630 22298 26682
rect 22052 26628 22058 26630
rect 22114 26628 22138 26630
rect 22194 26628 22218 26630
rect 22274 26628 22298 26630
rect 22354 26628 22360 26630
rect 22052 26619 22360 26628
rect 22388 26586 22416 26812
rect 22468 26784 22520 26790
rect 22468 26726 22520 26732
rect 22376 26580 22428 26586
rect 22296 26540 22376 26568
rect 22100 26444 22152 26450
rect 22100 26386 22152 26392
rect 21824 26308 21876 26314
rect 21824 26250 21876 26256
rect 21836 25974 21864 26250
rect 21916 26240 21968 26246
rect 21916 26182 21968 26188
rect 21928 26042 21956 26182
rect 21916 26036 21968 26042
rect 21916 25978 21968 25984
rect 21824 25968 21876 25974
rect 21824 25910 21876 25916
rect 21928 25362 21956 25978
rect 22112 25702 22140 26386
rect 22296 25906 22324 26540
rect 22376 26522 22428 26528
rect 22284 25900 22336 25906
rect 22284 25842 22336 25848
rect 22100 25696 22152 25702
rect 22100 25638 22152 25644
rect 22376 25696 22428 25702
rect 22376 25638 22428 25644
rect 22052 25596 22360 25605
rect 22052 25594 22058 25596
rect 22114 25594 22138 25596
rect 22194 25594 22218 25596
rect 22274 25594 22298 25596
rect 22354 25594 22360 25596
rect 22114 25542 22116 25594
rect 22296 25542 22298 25594
rect 22052 25540 22058 25542
rect 22114 25540 22138 25542
rect 22194 25540 22218 25542
rect 22274 25540 22298 25542
rect 22354 25540 22360 25542
rect 22052 25531 22360 25540
rect 22388 25498 22416 25638
rect 22376 25492 22428 25498
rect 22376 25434 22428 25440
rect 21732 25356 21784 25362
rect 21732 25298 21784 25304
rect 21916 25356 21968 25362
rect 21916 25298 21968 25304
rect 21640 25288 21692 25294
rect 21640 25230 21692 25236
rect 21824 25220 21876 25226
rect 21824 25162 21876 25168
rect 21548 24948 21600 24954
rect 21548 24890 21600 24896
rect 21456 24744 21508 24750
rect 21456 24686 21508 24692
rect 21560 24274 21588 24890
rect 21732 24336 21784 24342
rect 21732 24278 21784 24284
rect 21548 24268 21600 24274
rect 21548 24210 21600 24216
rect 21640 23656 21692 23662
rect 21640 23598 21692 23604
rect 21652 23254 21680 23598
rect 21640 23248 21692 23254
rect 21640 23190 21692 23196
rect 21364 23112 21416 23118
rect 21364 23054 21416 23060
rect 21548 23112 21600 23118
rect 21548 23054 21600 23060
rect 20810 22944 20866 22953
rect 20810 22879 20866 22888
rect 20824 22234 20852 22879
rect 21376 22642 21404 23054
rect 21560 22642 21588 23054
rect 21640 22976 21692 22982
rect 21640 22918 21692 22924
rect 21364 22636 21416 22642
rect 21364 22578 21416 22584
rect 21548 22636 21600 22642
rect 21548 22578 21600 22584
rect 21376 22234 21404 22578
rect 20812 22228 20864 22234
rect 20812 22170 20864 22176
rect 21364 22228 21416 22234
rect 21364 22170 21416 22176
rect 20824 21690 20852 22170
rect 21560 22166 21588 22578
rect 21548 22160 21600 22166
rect 21548 22102 21600 22108
rect 20904 22024 20956 22030
rect 20904 21966 20956 21972
rect 20996 22024 21048 22030
rect 20996 21966 21048 21972
rect 20812 21684 20864 21690
rect 20812 21626 20864 21632
rect 20720 21480 20772 21486
rect 20720 21422 20772 21428
rect 20628 21344 20680 21350
rect 20628 21286 20680 21292
rect 20640 21146 20668 21286
rect 20444 21140 20496 21146
rect 20444 21082 20496 21088
rect 20628 21140 20680 21146
rect 20628 21082 20680 21088
rect 20732 20942 20760 21422
rect 20916 21350 20944 21966
rect 20812 21344 20864 21350
rect 20812 21286 20864 21292
rect 20904 21344 20956 21350
rect 20904 21286 20956 21292
rect 20352 20936 20404 20942
rect 20352 20878 20404 20884
rect 20720 20936 20772 20942
rect 20720 20878 20772 20884
rect 20260 20256 20312 20262
rect 20260 20198 20312 20204
rect 20272 19786 20300 20198
rect 20364 20058 20392 20878
rect 20720 20596 20772 20602
rect 20720 20538 20772 20544
rect 20536 20256 20588 20262
rect 20536 20198 20588 20204
rect 20548 20058 20576 20198
rect 20352 20052 20404 20058
rect 20352 19994 20404 20000
rect 20536 20052 20588 20058
rect 20536 19994 20588 20000
rect 20260 19780 20312 19786
rect 20260 19722 20312 19728
rect 20732 19514 20760 20538
rect 20824 20534 20852 21286
rect 20812 20528 20864 20534
rect 20812 20470 20864 20476
rect 20812 20324 20864 20330
rect 20812 20266 20864 20272
rect 20824 20058 20852 20266
rect 20812 20052 20864 20058
rect 20812 19994 20864 20000
rect 20720 19508 20772 19514
rect 20720 19450 20772 19456
rect 20916 19310 20944 21286
rect 21008 20058 21036 21966
rect 21272 21888 21324 21894
rect 21272 21830 21324 21836
rect 21088 21616 21140 21622
rect 21088 21558 21140 21564
rect 20996 20052 21048 20058
rect 20996 19994 21048 20000
rect 21100 19854 21128 21558
rect 21284 21554 21312 21830
rect 21548 21616 21600 21622
rect 21652 21604 21680 22918
rect 21744 22642 21772 24278
rect 21836 24206 21864 25162
rect 22480 24818 22508 26726
rect 22652 26376 22704 26382
rect 22652 26318 22704 26324
rect 22664 25974 22692 26318
rect 22652 25968 22704 25974
rect 22652 25910 22704 25916
rect 22560 25696 22612 25702
rect 22560 25638 22612 25644
rect 22652 25696 22704 25702
rect 22652 25638 22704 25644
rect 22572 25226 22600 25638
rect 22560 25220 22612 25226
rect 22560 25162 22612 25168
rect 22664 24954 22692 25638
rect 22652 24948 22704 24954
rect 22652 24890 22704 24896
rect 22468 24812 22520 24818
rect 22468 24754 22520 24760
rect 22052 24508 22360 24517
rect 22052 24506 22058 24508
rect 22114 24506 22138 24508
rect 22194 24506 22218 24508
rect 22274 24506 22298 24508
rect 22354 24506 22360 24508
rect 22114 24454 22116 24506
rect 22296 24454 22298 24506
rect 22052 24452 22058 24454
rect 22114 24452 22138 24454
rect 22194 24452 22218 24454
rect 22274 24452 22298 24454
rect 22354 24452 22360 24454
rect 22052 24443 22360 24452
rect 21824 24200 21876 24206
rect 21824 24142 21876 24148
rect 21836 23118 21864 24142
rect 22284 24064 22336 24070
rect 22284 24006 22336 24012
rect 22296 23633 22324 24006
rect 22480 23866 22508 24754
rect 22756 24698 22784 26930
rect 23032 26926 23060 27610
rect 23296 27464 23348 27470
rect 23296 27406 23348 27412
rect 23308 27130 23336 27406
rect 23296 27124 23348 27130
rect 23296 27066 23348 27072
rect 23204 27056 23256 27062
rect 23204 26998 23256 27004
rect 23020 26920 23072 26926
rect 22848 26880 23020 26908
rect 22848 25362 22876 26880
rect 23020 26862 23072 26868
rect 23216 26518 23244 26998
rect 23204 26512 23256 26518
rect 23204 26454 23256 26460
rect 23216 26382 23244 26454
rect 23204 26376 23256 26382
rect 23204 26318 23256 26324
rect 23112 26240 23164 26246
rect 23112 26182 23164 26188
rect 23124 25906 23152 26182
rect 23112 25900 23164 25906
rect 23112 25842 23164 25848
rect 23860 25838 23888 27814
rect 23952 27418 23980 29106
rect 24216 28960 24268 28966
rect 24216 28902 24268 28908
rect 24228 28558 24256 28902
rect 30493 28860 30801 28869
rect 30493 28858 30499 28860
rect 30555 28858 30579 28860
rect 30635 28858 30659 28860
rect 30715 28858 30739 28860
rect 30795 28858 30801 28860
rect 30555 28806 30557 28858
rect 30737 28806 30739 28858
rect 30493 28804 30499 28806
rect 30555 28804 30579 28806
rect 30635 28804 30659 28806
rect 30715 28804 30739 28806
rect 30795 28804 30801 28806
rect 30493 28795 30801 28804
rect 24216 28552 24268 28558
rect 24216 28494 24268 28500
rect 26272 28316 26580 28325
rect 26272 28314 26278 28316
rect 26334 28314 26358 28316
rect 26414 28314 26438 28316
rect 26494 28314 26518 28316
rect 26574 28314 26580 28316
rect 26334 28262 26336 28314
rect 26516 28262 26518 28314
rect 26272 28260 26278 28262
rect 26334 28260 26358 28262
rect 26414 28260 26438 28262
rect 26494 28260 26518 28262
rect 26574 28260 26580 28262
rect 26272 28251 26580 28260
rect 34713 28316 35021 28325
rect 34713 28314 34719 28316
rect 34775 28314 34799 28316
rect 34855 28314 34879 28316
rect 34935 28314 34959 28316
rect 35015 28314 35021 28316
rect 34775 28262 34777 28314
rect 34957 28262 34959 28314
rect 34713 28260 34719 28262
rect 34775 28260 34799 28262
rect 34855 28260 34879 28262
rect 34935 28260 34959 28262
rect 35015 28260 35021 28262
rect 34713 28251 35021 28260
rect 30493 27772 30801 27781
rect 30493 27770 30499 27772
rect 30555 27770 30579 27772
rect 30635 27770 30659 27772
rect 30715 27770 30739 27772
rect 30795 27770 30801 27772
rect 30555 27718 30557 27770
rect 30737 27718 30739 27770
rect 30493 27716 30499 27718
rect 30555 27716 30579 27718
rect 30635 27716 30659 27718
rect 30715 27716 30739 27718
rect 30795 27716 30801 27718
rect 30493 27707 30801 27716
rect 34520 27464 34572 27470
rect 34518 27432 34520 27441
rect 34572 27432 34574 27441
rect 23952 27390 24072 27418
rect 23940 27328 23992 27334
rect 23940 27270 23992 27276
rect 23952 27130 23980 27270
rect 23940 27124 23992 27130
rect 23940 27066 23992 27072
rect 23756 25832 23808 25838
rect 23756 25774 23808 25780
rect 23848 25832 23900 25838
rect 23848 25774 23900 25780
rect 23112 25696 23164 25702
rect 23112 25638 23164 25644
rect 22836 25356 22888 25362
rect 22836 25298 22888 25304
rect 23124 25294 23152 25638
rect 23112 25288 23164 25294
rect 23112 25230 23164 25236
rect 23020 25220 23072 25226
rect 23020 25162 23072 25168
rect 23032 24818 23060 25162
rect 23020 24812 23072 24818
rect 23020 24754 23072 24760
rect 23768 24750 23796 25774
rect 23860 25158 23888 25774
rect 23848 25152 23900 25158
rect 23848 25094 23900 25100
rect 22664 24682 22784 24698
rect 23756 24744 23808 24750
rect 23756 24686 23808 24692
rect 22652 24676 22784 24682
rect 22704 24670 22784 24676
rect 22652 24618 22704 24624
rect 22664 24410 22692 24618
rect 22652 24404 22704 24410
rect 22652 24346 22704 24352
rect 22560 24336 22612 24342
rect 22560 24278 22612 24284
rect 22376 23860 22428 23866
rect 22376 23802 22428 23808
rect 22468 23860 22520 23866
rect 22468 23802 22520 23808
rect 22282 23624 22338 23633
rect 21928 23582 22282 23610
rect 21928 23186 21956 23582
rect 22282 23559 22338 23568
rect 22052 23420 22360 23429
rect 22052 23418 22058 23420
rect 22114 23418 22138 23420
rect 22194 23418 22218 23420
rect 22274 23418 22298 23420
rect 22354 23418 22360 23420
rect 22114 23366 22116 23418
rect 22296 23366 22298 23418
rect 22052 23364 22058 23366
rect 22114 23364 22138 23366
rect 22194 23364 22218 23366
rect 22274 23364 22298 23366
rect 22354 23364 22360 23366
rect 22052 23355 22360 23364
rect 22192 23316 22244 23322
rect 22192 23258 22244 23264
rect 21916 23180 21968 23186
rect 22204 23168 22232 23258
rect 21916 23122 21968 23128
rect 22112 23140 22232 23168
rect 21824 23112 21876 23118
rect 21824 23054 21876 23060
rect 22008 23112 22060 23118
rect 22112 23100 22140 23140
rect 22060 23072 22140 23100
rect 22008 23054 22060 23060
rect 21916 23044 21968 23050
rect 21916 22986 21968 22992
rect 21732 22636 21784 22642
rect 21732 22578 21784 22584
rect 21600 21576 21680 21604
rect 21548 21558 21600 21564
rect 21272 21548 21324 21554
rect 21744 21536 21772 22578
rect 21928 22234 21956 22986
rect 22006 22808 22062 22817
rect 22006 22743 22008 22752
rect 22060 22743 22062 22752
rect 22008 22714 22060 22720
rect 22112 22506 22140 23072
rect 22388 23066 22416 23802
rect 22468 23656 22520 23662
rect 22468 23598 22520 23604
rect 22480 23322 22508 23598
rect 22572 23526 22600 24278
rect 22664 23730 22692 24346
rect 23204 24200 23256 24206
rect 23204 24142 23256 24148
rect 22928 24064 22980 24070
rect 22928 24006 22980 24012
rect 22940 23866 22968 24006
rect 23216 23866 23244 24142
rect 23848 24064 23900 24070
rect 23848 24006 23900 24012
rect 23860 23866 23888 24006
rect 22928 23860 22980 23866
rect 22928 23802 22980 23808
rect 23204 23860 23256 23866
rect 23204 23802 23256 23808
rect 23848 23860 23900 23866
rect 23848 23802 23900 23808
rect 22652 23724 22704 23730
rect 22652 23666 22704 23672
rect 23664 23724 23716 23730
rect 23664 23666 23716 23672
rect 22560 23520 22612 23526
rect 22560 23462 22612 23468
rect 22572 23322 22600 23462
rect 22468 23316 22520 23322
rect 22468 23258 22520 23264
rect 22560 23316 22612 23322
rect 22560 23258 22612 23264
rect 22204 23038 22416 23066
rect 22468 23112 22520 23118
rect 22468 23054 22520 23060
rect 22204 22778 22232 23038
rect 22284 22976 22336 22982
rect 22284 22918 22336 22924
rect 22374 22944 22430 22953
rect 22192 22772 22244 22778
rect 22192 22714 22244 22720
rect 22296 22692 22324 22918
rect 22480 22930 22508 23054
rect 22430 22902 22508 22930
rect 22560 22976 22612 22982
rect 22560 22918 22612 22924
rect 22374 22879 22430 22888
rect 22572 22778 22600 22918
rect 22560 22772 22612 22778
rect 22560 22714 22612 22720
rect 22468 22704 22520 22710
rect 22296 22664 22468 22692
rect 22468 22646 22520 22652
rect 22376 22568 22428 22574
rect 22664 22556 22692 23666
rect 22836 23656 22888 23662
rect 22836 23598 22888 23604
rect 23018 23624 23074 23633
rect 22848 22574 22876 23598
rect 23018 23559 23074 23568
rect 23032 23186 23060 23559
rect 23020 23180 23072 23186
rect 23020 23122 23072 23128
rect 22928 23112 22980 23118
rect 22928 23054 22980 23060
rect 22940 22778 22968 23054
rect 23296 22976 23348 22982
rect 23296 22918 23348 22924
rect 22928 22772 22980 22778
rect 22928 22714 22980 22720
rect 23308 22710 23336 22918
rect 23296 22704 23348 22710
rect 23296 22646 23348 22652
rect 23572 22636 23624 22642
rect 23572 22578 23624 22584
rect 22428 22528 22692 22556
rect 22836 22568 22888 22574
rect 22376 22510 22428 22516
rect 22836 22510 22888 22516
rect 22100 22500 22152 22506
rect 22100 22442 22152 22448
rect 22052 22332 22360 22341
rect 22052 22330 22058 22332
rect 22114 22330 22138 22332
rect 22194 22330 22218 22332
rect 22274 22330 22298 22332
rect 22354 22330 22360 22332
rect 22114 22278 22116 22330
rect 22296 22278 22298 22330
rect 22052 22276 22058 22278
rect 22114 22276 22138 22278
rect 22194 22276 22218 22278
rect 22274 22276 22298 22278
rect 22354 22276 22360 22278
rect 22052 22267 22360 22276
rect 21916 22228 21968 22234
rect 21916 22170 21968 22176
rect 21916 22092 21968 22098
rect 21916 22034 21968 22040
rect 21824 21684 21876 21690
rect 21824 21626 21876 21632
rect 21836 21554 21864 21626
rect 21272 21490 21324 21496
rect 21652 21508 21772 21536
rect 21824 21548 21876 21554
rect 21548 20936 21600 20942
rect 21652 20924 21680 21508
rect 21824 21490 21876 21496
rect 21732 21344 21784 21350
rect 21732 21286 21784 21292
rect 21744 21078 21772 21286
rect 21732 21072 21784 21078
rect 21732 21014 21784 21020
rect 21600 20896 21680 20924
rect 21732 20936 21784 20942
rect 21548 20878 21600 20884
rect 21732 20878 21784 20884
rect 21180 20596 21232 20602
rect 21180 20538 21232 20544
rect 21088 19848 21140 19854
rect 21088 19790 21140 19796
rect 21192 19718 21220 20538
rect 21548 20324 21600 20330
rect 21548 20266 21600 20272
rect 21180 19712 21232 19718
rect 21180 19654 21232 19660
rect 21560 19514 21588 20266
rect 21744 20058 21772 20878
rect 21836 20466 21864 21490
rect 21824 20460 21876 20466
rect 21824 20402 21876 20408
rect 21732 20052 21784 20058
rect 21732 19994 21784 20000
rect 21836 19854 21864 20402
rect 21928 20398 21956 22034
rect 22388 21350 22416 22510
rect 22468 22024 22520 22030
rect 22468 21966 22520 21972
rect 22480 21690 22508 21966
rect 22468 21684 22520 21690
rect 22468 21626 22520 21632
rect 22376 21344 22428 21350
rect 22376 21286 22428 21292
rect 22052 21244 22360 21253
rect 22052 21242 22058 21244
rect 22114 21242 22138 21244
rect 22194 21242 22218 21244
rect 22274 21242 22298 21244
rect 22354 21242 22360 21244
rect 22114 21190 22116 21242
rect 22296 21190 22298 21242
rect 22052 21188 22058 21190
rect 22114 21188 22138 21190
rect 22194 21188 22218 21190
rect 22274 21188 22298 21190
rect 22354 21188 22360 21190
rect 22052 21179 22360 21188
rect 22284 21140 22336 21146
rect 22284 21082 22336 21088
rect 22296 20942 22324 21082
rect 22284 20936 22336 20942
rect 22204 20896 22284 20924
rect 22204 20466 22232 20896
rect 22284 20878 22336 20884
rect 22376 20936 22428 20942
rect 22376 20878 22428 20884
rect 22284 20800 22336 20806
rect 22284 20742 22336 20748
rect 22296 20466 22324 20742
rect 22192 20460 22244 20466
rect 22192 20402 22244 20408
rect 22284 20460 22336 20466
rect 22284 20402 22336 20408
rect 21916 20392 21968 20398
rect 21916 20334 21968 20340
rect 21916 20256 21968 20262
rect 21916 20198 21968 20204
rect 21928 19854 21956 20198
rect 22052 20156 22360 20165
rect 22052 20154 22058 20156
rect 22114 20154 22138 20156
rect 22194 20154 22218 20156
rect 22274 20154 22298 20156
rect 22354 20154 22360 20156
rect 22114 20102 22116 20154
rect 22296 20102 22298 20154
rect 22052 20100 22058 20102
rect 22114 20100 22138 20102
rect 22194 20100 22218 20102
rect 22274 20100 22298 20102
rect 22354 20100 22360 20102
rect 22052 20091 22360 20100
rect 22388 19922 22416 20878
rect 22480 20262 22508 21626
rect 22652 21548 22704 21554
rect 22652 21490 22704 21496
rect 22560 21344 22612 21350
rect 22560 21286 22612 21292
rect 22572 21146 22600 21286
rect 22560 21140 22612 21146
rect 22560 21082 22612 21088
rect 22468 20256 22520 20262
rect 22468 20198 22520 20204
rect 22480 20058 22508 20198
rect 22664 20058 22692 21490
rect 22848 20874 22876 22510
rect 23584 22030 23612 22578
rect 23676 22234 23704 23666
rect 23848 23044 23900 23050
rect 23848 22986 23900 22992
rect 23860 22817 23888 22986
rect 23846 22808 23902 22817
rect 23846 22743 23902 22752
rect 23664 22228 23716 22234
rect 23664 22170 23716 22176
rect 23572 22024 23624 22030
rect 23572 21966 23624 21972
rect 23480 21480 23532 21486
rect 23480 21422 23532 21428
rect 23492 21146 23520 21422
rect 23480 21140 23532 21146
rect 23480 21082 23532 21088
rect 22744 20868 22796 20874
rect 22744 20810 22796 20816
rect 22836 20868 22888 20874
rect 22836 20810 22888 20816
rect 22756 20534 22784 20810
rect 23572 20800 23624 20806
rect 23572 20742 23624 20748
rect 23584 20534 23612 20742
rect 22744 20528 22796 20534
rect 22744 20470 22796 20476
rect 23572 20528 23624 20534
rect 23572 20470 23624 20476
rect 23204 20460 23256 20466
rect 23204 20402 23256 20408
rect 23216 20058 23244 20402
rect 22468 20052 22520 20058
rect 22468 19994 22520 20000
rect 22652 20052 22704 20058
rect 22652 19994 22704 20000
rect 23204 20052 23256 20058
rect 23204 19994 23256 20000
rect 22376 19916 22428 19922
rect 22376 19858 22428 19864
rect 21824 19848 21876 19854
rect 21824 19790 21876 19796
rect 21916 19848 21968 19854
rect 21916 19790 21968 19796
rect 22284 19780 22336 19786
rect 22284 19722 22336 19728
rect 22296 19514 22324 19722
rect 22664 19718 22692 19994
rect 22652 19712 22704 19718
rect 22652 19654 22704 19660
rect 21548 19508 21600 19514
rect 21548 19450 21600 19456
rect 22284 19508 22336 19514
rect 22284 19450 22336 19456
rect 20904 19304 20956 19310
rect 20904 19246 20956 19252
rect 22052 19068 22360 19077
rect 22052 19066 22058 19068
rect 22114 19066 22138 19068
rect 22194 19066 22218 19068
rect 22274 19066 22298 19068
rect 22354 19066 22360 19068
rect 22114 19014 22116 19066
rect 22296 19014 22298 19066
rect 22052 19012 22058 19014
rect 22114 19012 22138 19014
rect 22194 19012 22218 19014
rect 22274 19012 22298 19014
rect 22354 19012 22360 19014
rect 22052 19003 22360 19012
rect 22052 17980 22360 17989
rect 22052 17978 22058 17980
rect 22114 17978 22138 17980
rect 22194 17978 22218 17980
rect 22274 17978 22298 17980
rect 22354 17978 22360 17980
rect 22114 17926 22116 17978
rect 22296 17926 22298 17978
rect 22052 17924 22058 17926
rect 22114 17924 22138 17926
rect 22194 17924 22218 17926
rect 22274 17924 22298 17926
rect 22354 17924 22360 17926
rect 22052 17915 22360 17924
rect 22052 16892 22360 16901
rect 22052 16890 22058 16892
rect 22114 16890 22138 16892
rect 22194 16890 22218 16892
rect 22274 16890 22298 16892
rect 22354 16890 22360 16892
rect 22114 16838 22116 16890
rect 22296 16838 22298 16890
rect 22052 16836 22058 16838
rect 22114 16836 22138 16838
rect 22194 16836 22218 16838
rect 22274 16836 22298 16838
rect 22354 16836 22360 16838
rect 22052 16827 22360 16836
rect 22052 15804 22360 15813
rect 22052 15802 22058 15804
rect 22114 15802 22138 15804
rect 22194 15802 22218 15804
rect 22274 15802 22298 15804
rect 22354 15802 22360 15804
rect 22114 15750 22116 15802
rect 22296 15750 22298 15802
rect 22052 15748 22058 15750
rect 22114 15748 22138 15750
rect 22194 15748 22218 15750
rect 22274 15748 22298 15750
rect 22354 15748 22360 15750
rect 22052 15739 22360 15748
rect 22052 14716 22360 14725
rect 22052 14714 22058 14716
rect 22114 14714 22138 14716
rect 22194 14714 22218 14716
rect 22274 14714 22298 14716
rect 22354 14714 22360 14716
rect 22114 14662 22116 14714
rect 22296 14662 22298 14714
rect 22052 14660 22058 14662
rect 22114 14660 22138 14662
rect 22194 14660 22218 14662
rect 22274 14660 22298 14662
rect 22354 14660 22360 14662
rect 22052 14651 22360 14660
rect 22052 13628 22360 13637
rect 22052 13626 22058 13628
rect 22114 13626 22138 13628
rect 22194 13626 22218 13628
rect 22274 13626 22298 13628
rect 22354 13626 22360 13628
rect 22114 13574 22116 13626
rect 22296 13574 22298 13626
rect 22052 13572 22058 13574
rect 22114 13572 22138 13574
rect 22194 13572 22218 13574
rect 22274 13572 22298 13574
rect 22354 13572 22360 13574
rect 22052 13563 22360 13572
rect 24044 13190 24072 27390
rect 34518 27367 34574 27376
rect 24584 27328 24636 27334
rect 24584 27270 24636 27276
rect 24860 27328 24912 27334
rect 24860 27270 24912 27276
rect 24596 26790 24624 27270
rect 24872 26994 24900 27270
rect 26272 27228 26580 27237
rect 26272 27226 26278 27228
rect 26334 27226 26358 27228
rect 26414 27226 26438 27228
rect 26494 27226 26518 27228
rect 26574 27226 26580 27228
rect 26334 27174 26336 27226
rect 26516 27174 26518 27226
rect 26272 27172 26278 27174
rect 26334 27172 26358 27174
rect 26414 27172 26438 27174
rect 26494 27172 26518 27174
rect 26574 27172 26580 27174
rect 26272 27163 26580 27172
rect 34713 27228 35021 27237
rect 34713 27226 34719 27228
rect 34775 27226 34799 27228
rect 34855 27226 34879 27228
rect 34935 27226 34959 27228
rect 35015 27226 35021 27228
rect 34775 27174 34777 27226
rect 34957 27174 34959 27226
rect 34713 27172 34719 27174
rect 34775 27172 34799 27174
rect 34855 27172 34879 27174
rect 34935 27172 34959 27174
rect 35015 27172 35021 27174
rect 34713 27163 35021 27172
rect 24860 26988 24912 26994
rect 24860 26930 24912 26936
rect 24584 26784 24636 26790
rect 24584 26726 24636 26732
rect 24596 26489 24624 26726
rect 30493 26684 30801 26693
rect 30493 26682 30499 26684
rect 30555 26682 30579 26684
rect 30635 26682 30659 26684
rect 30715 26682 30739 26684
rect 30795 26682 30801 26684
rect 30555 26630 30557 26682
rect 30737 26630 30739 26682
rect 30493 26628 30499 26630
rect 30555 26628 30579 26630
rect 30635 26628 30659 26630
rect 30715 26628 30739 26630
rect 30795 26628 30801 26630
rect 30493 26619 30801 26628
rect 24582 26480 24638 26489
rect 24582 26415 24638 26424
rect 26272 26140 26580 26149
rect 26272 26138 26278 26140
rect 26334 26138 26358 26140
rect 26414 26138 26438 26140
rect 26494 26138 26518 26140
rect 26574 26138 26580 26140
rect 26334 26086 26336 26138
rect 26516 26086 26518 26138
rect 26272 26084 26278 26086
rect 26334 26084 26358 26086
rect 26414 26084 26438 26086
rect 26494 26084 26518 26086
rect 26574 26084 26580 26086
rect 26272 26075 26580 26084
rect 34713 26140 35021 26149
rect 34713 26138 34719 26140
rect 34775 26138 34799 26140
rect 34855 26138 34879 26140
rect 34935 26138 34959 26140
rect 35015 26138 35021 26140
rect 34775 26086 34777 26138
rect 34957 26086 34959 26138
rect 34713 26084 34719 26086
rect 34775 26084 34799 26086
rect 34855 26084 34879 26086
rect 34935 26084 34959 26086
rect 35015 26084 35021 26086
rect 34713 26075 35021 26084
rect 30493 25596 30801 25605
rect 30493 25594 30499 25596
rect 30555 25594 30579 25596
rect 30635 25594 30659 25596
rect 30715 25594 30739 25596
rect 30795 25594 30801 25596
rect 30555 25542 30557 25594
rect 30737 25542 30739 25594
rect 30493 25540 30499 25542
rect 30555 25540 30579 25542
rect 30635 25540 30659 25542
rect 30715 25540 30739 25542
rect 30795 25540 30801 25542
rect 30493 25531 30801 25540
rect 24216 25288 24268 25294
rect 24216 25230 24268 25236
rect 24228 25158 24256 25230
rect 24216 25152 24268 25158
rect 24216 25094 24268 25100
rect 24860 25152 24912 25158
rect 24860 25094 24912 25100
rect 24228 24614 24256 25094
rect 24872 24818 24900 25094
rect 26272 25052 26580 25061
rect 26272 25050 26278 25052
rect 26334 25050 26358 25052
rect 26414 25050 26438 25052
rect 26494 25050 26518 25052
rect 26574 25050 26580 25052
rect 26334 24998 26336 25050
rect 26516 24998 26518 25050
rect 26272 24996 26278 24998
rect 26334 24996 26358 24998
rect 26414 24996 26438 24998
rect 26494 24996 26518 24998
rect 26574 24996 26580 24998
rect 26272 24987 26580 24996
rect 34713 25052 35021 25061
rect 34713 25050 34719 25052
rect 34775 25050 34799 25052
rect 34855 25050 34879 25052
rect 34935 25050 34959 25052
rect 35015 25050 35021 25052
rect 34775 24998 34777 25050
rect 34957 24998 34959 25050
rect 34713 24996 34719 24998
rect 34775 24996 34799 24998
rect 34855 24996 34879 24998
rect 34935 24996 34959 24998
rect 35015 24996 35021 24998
rect 34713 24987 35021 24996
rect 24860 24812 24912 24818
rect 24860 24754 24912 24760
rect 24216 24608 24268 24614
rect 24216 24550 24268 24556
rect 30493 24508 30801 24517
rect 30493 24506 30499 24508
rect 30555 24506 30579 24508
rect 30635 24506 30659 24508
rect 30715 24506 30739 24508
rect 30795 24506 30801 24508
rect 30555 24454 30557 24506
rect 30737 24454 30739 24506
rect 30493 24452 30499 24454
rect 30555 24452 30579 24454
rect 30635 24452 30659 24454
rect 30715 24452 30739 24454
rect 30795 24452 30801 24454
rect 30493 24443 30801 24452
rect 24492 24064 24544 24070
rect 24492 24006 24544 24012
rect 24584 24064 24636 24070
rect 24584 24006 24636 24012
rect 24504 23526 24532 24006
rect 24596 23730 24624 24006
rect 26272 23964 26580 23973
rect 26272 23962 26278 23964
rect 26334 23962 26358 23964
rect 26414 23962 26438 23964
rect 26494 23962 26518 23964
rect 26574 23962 26580 23964
rect 26334 23910 26336 23962
rect 26516 23910 26518 23962
rect 26272 23908 26278 23910
rect 26334 23908 26358 23910
rect 26414 23908 26438 23910
rect 26494 23908 26518 23910
rect 26574 23908 26580 23910
rect 26272 23899 26580 23908
rect 34713 23964 35021 23973
rect 34713 23962 34719 23964
rect 34775 23962 34799 23964
rect 34855 23962 34879 23964
rect 34935 23962 34959 23964
rect 35015 23962 35021 23964
rect 34775 23910 34777 23962
rect 34957 23910 34959 23962
rect 34713 23908 34719 23910
rect 34775 23908 34799 23910
rect 34855 23908 34879 23910
rect 34935 23908 34959 23910
rect 35015 23908 35021 23910
rect 34713 23899 35021 23908
rect 24584 23724 24636 23730
rect 24584 23666 24636 23672
rect 24492 23520 24544 23526
rect 24492 23462 24544 23468
rect 24504 23225 24532 23462
rect 30493 23420 30801 23429
rect 30493 23418 30499 23420
rect 30555 23418 30579 23420
rect 30635 23418 30659 23420
rect 30715 23418 30739 23420
rect 30795 23418 30801 23420
rect 30555 23366 30557 23418
rect 30737 23366 30739 23418
rect 30493 23364 30499 23366
rect 30555 23364 30579 23366
rect 30635 23364 30659 23366
rect 30715 23364 30739 23366
rect 30795 23364 30801 23366
rect 30493 23355 30801 23364
rect 24490 23216 24546 23225
rect 24400 23180 24452 23186
rect 24490 23151 24546 23160
rect 24400 23122 24452 23128
rect 24124 22976 24176 22982
rect 24124 22918 24176 22924
rect 24216 22976 24268 22982
rect 24216 22918 24268 22924
rect 24308 22976 24360 22982
rect 24308 22918 24360 22924
rect 24136 22642 24164 22918
rect 24124 22636 24176 22642
rect 24124 22578 24176 22584
rect 24228 22438 24256 22918
rect 24216 22432 24268 22438
rect 24216 22374 24268 22380
rect 24320 22098 24348 22918
rect 24412 22778 24440 23122
rect 26272 22876 26580 22885
rect 26272 22874 26278 22876
rect 26334 22874 26358 22876
rect 26414 22874 26438 22876
rect 26494 22874 26518 22876
rect 26574 22874 26580 22876
rect 26334 22822 26336 22874
rect 26516 22822 26518 22874
rect 26272 22820 26278 22822
rect 26334 22820 26358 22822
rect 26414 22820 26438 22822
rect 26494 22820 26518 22822
rect 26574 22820 26580 22822
rect 26272 22811 26580 22820
rect 34713 22876 35021 22885
rect 34713 22874 34719 22876
rect 34775 22874 34799 22876
rect 34855 22874 34879 22876
rect 34935 22874 34959 22876
rect 35015 22874 35021 22876
rect 34775 22822 34777 22874
rect 34957 22822 34959 22874
rect 34713 22820 34719 22822
rect 34775 22820 34799 22822
rect 34855 22820 34879 22822
rect 34935 22820 34959 22822
rect 35015 22820 35021 22822
rect 34713 22811 35021 22820
rect 24400 22772 24452 22778
rect 24400 22714 24452 22720
rect 30493 22332 30801 22341
rect 30493 22330 30499 22332
rect 30555 22330 30579 22332
rect 30635 22330 30659 22332
rect 30715 22330 30739 22332
rect 30795 22330 30801 22332
rect 30555 22278 30557 22330
rect 30737 22278 30739 22330
rect 30493 22276 30499 22278
rect 30555 22276 30579 22278
rect 30635 22276 30659 22278
rect 30715 22276 30739 22278
rect 30795 22276 30801 22278
rect 30493 22267 30801 22276
rect 24308 22092 24360 22098
rect 24308 22034 24360 22040
rect 26272 21788 26580 21797
rect 26272 21786 26278 21788
rect 26334 21786 26358 21788
rect 26414 21786 26438 21788
rect 26494 21786 26518 21788
rect 26574 21786 26580 21788
rect 26334 21734 26336 21786
rect 26516 21734 26518 21786
rect 26272 21732 26278 21734
rect 26334 21732 26358 21734
rect 26414 21732 26438 21734
rect 26494 21732 26518 21734
rect 26574 21732 26580 21734
rect 26272 21723 26580 21732
rect 34713 21788 35021 21797
rect 34713 21786 34719 21788
rect 34775 21786 34799 21788
rect 34855 21786 34879 21788
rect 34935 21786 34959 21788
rect 35015 21786 35021 21788
rect 34775 21734 34777 21786
rect 34957 21734 34959 21786
rect 34713 21732 34719 21734
rect 34775 21732 34799 21734
rect 34855 21732 34879 21734
rect 34935 21732 34959 21734
rect 35015 21732 35021 21734
rect 34713 21723 35021 21732
rect 30493 21244 30801 21253
rect 30493 21242 30499 21244
rect 30555 21242 30579 21244
rect 30635 21242 30659 21244
rect 30715 21242 30739 21244
rect 30795 21242 30801 21244
rect 30555 21190 30557 21242
rect 30737 21190 30739 21242
rect 30493 21188 30499 21190
rect 30555 21188 30579 21190
rect 30635 21188 30659 21190
rect 30715 21188 30739 21190
rect 30795 21188 30801 21190
rect 30493 21179 30801 21188
rect 26272 20700 26580 20709
rect 26272 20698 26278 20700
rect 26334 20698 26358 20700
rect 26414 20698 26438 20700
rect 26494 20698 26518 20700
rect 26574 20698 26580 20700
rect 26334 20646 26336 20698
rect 26516 20646 26518 20698
rect 26272 20644 26278 20646
rect 26334 20644 26358 20646
rect 26414 20644 26438 20646
rect 26494 20644 26518 20646
rect 26574 20644 26580 20646
rect 26272 20635 26580 20644
rect 34713 20700 35021 20709
rect 34713 20698 34719 20700
rect 34775 20698 34799 20700
rect 34855 20698 34879 20700
rect 34935 20698 34959 20700
rect 35015 20698 35021 20700
rect 34775 20646 34777 20698
rect 34957 20646 34959 20698
rect 34713 20644 34719 20646
rect 34775 20644 34799 20646
rect 34855 20644 34879 20646
rect 34935 20644 34959 20646
rect 35015 20644 35021 20646
rect 34713 20635 35021 20644
rect 33140 20256 33192 20262
rect 33140 20198 33192 20204
rect 30493 20156 30801 20165
rect 30493 20154 30499 20156
rect 30555 20154 30579 20156
rect 30635 20154 30659 20156
rect 30715 20154 30739 20156
rect 30795 20154 30801 20156
rect 30555 20102 30557 20154
rect 30737 20102 30739 20154
rect 30493 20100 30499 20102
rect 30555 20100 30579 20102
rect 30635 20100 30659 20102
rect 30715 20100 30739 20102
rect 30795 20100 30801 20102
rect 30493 20091 30801 20100
rect 33152 19854 33180 20198
rect 33140 19848 33192 19854
rect 33140 19790 33192 19796
rect 34610 19816 34666 19825
rect 34610 19751 34612 19760
rect 34664 19751 34666 19760
rect 34612 19722 34664 19728
rect 26272 19612 26580 19621
rect 26272 19610 26278 19612
rect 26334 19610 26358 19612
rect 26414 19610 26438 19612
rect 26494 19610 26518 19612
rect 26574 19610 26580 19612
rect 26334 19558 26336 19610
rect 26516 19558 26518 19610
rect 26272 19556 26278 19558
rect 26334 19556 26358 19558
rect 26414 19556 26438 19558
rect 26494 19556 26518 19558
rect 26574 19556 26580 19558
rect 26272 19547 26580 19556
rect 34713 19612 35021 19621
rect 34713 19610 34719 19612
rect 34775 19610 34799 19612
rect 34855 19610 34879 19612
rect 34935 19610 34959 19612
rect 35015 19610 35021 19612
rect 34775 19558 34777 19610
rect 34957 19558 34959 19610
rect 34713 19556 34719 19558
rect 34775 19556 34799 19558
rect 34855 19556 34879 19558
rect 34935 19556 34959 19558
rect 35015 19556 35021 19558
rect 34713 19547 35021 19556
rect 30493 19068 30801 19077
rect 30493 19066 30499 19068
rect 30555 19066 30579 19068
rect 30635 19066 30659 19068
rect 30715 19066 30739 19068
rect 30795 19066 30801 19068
rect 30555 19014 30557 19066
rect 30737 19014 30739 19066
rect 30493 19012 30499 19014
rect 30555 19012 30579 19014
rect 30635 19012 30659 19014
rect 30715 19012 30739 19014
rect 30795 19012 30801 19014
rect 30493 19003 30801 19012
rect 26272 18524 26580 18533
rect 26272 18522 26278 18524
rect 26334 18522 26358 18524
rect 26414 18522 26438 18524
rect 26494 18522 26518 18524
rect 26574 18522 26580 18524
rect 26334 18470 26336 18522
rect 26516 18470 26518 18522
rect 26272 18468 26278 18470
rect 26334 18468 26358 18470
rect 26414 18468 26438 18470
rect 26494 18468 26518 18470
rect 26574 18468 26580 18470
rect 26272 18459 26580 18468
rect 34713 18524 35021 18533
rect 34713 18522 34719 18524
rect 34775 18522 34799 18524
rect 34855 18522 34879 18524
rect 34935 18522 34959 18524
rect 35015 18522 35021 18524
rect 34775 18470 34777 18522
rect 34957 18470 34959 18522
rect 34713 18468 34719 18470
rect 34775 18468 34799 18470
rect 34855 18468 34879 18470
rect 34935 18468 34959 18470
rect 35015 18468 35021 18470
rect 34713 18459 35021 18468
rect 30493 17980 30801 17989
rect 30493 17978 30499 17980
rect 30555 17978 30579 17980
rect 30635 17978 30659 17980
rect 30715 17978 30739 17980
rect 30795 17978 30801 17980
rect 30555 17926 30557 17978
rect 30737 17926 30739 17978
rect 30493 17924 30499 17926
rect 30555 17924 30579 17926
rect 30635 17924 30659 17926
rect 30715 17924 30739 17926
rect 30795 17924 30801 17926
rect 30493 17915 30801 17924
rect 26272 17436 26580 17445
rect 26272 17434 26278 17436
rect 26334 17434 26358 17436
rect 26414 17434 26438 17436
rect 26494 17434 26518 17436
rect 26574 17434 26580 17436
rect 26334 17382 26336 17434
rect 26516 17382 26518 17434
rect 26272 17380 26278 17382
rect 26334 17380 26358 17382
rect 26414 17380 26438 17382
rect 26494 17380 26518 17382
rect 26574 17380 26580 17382
rect 26272 17371 26580 17380
rect 34713 17436 35021 17445
rect 34713 17434 34719 17436
rect 34775 17434 34799 17436
rect 34855 17434 34879 17436
rect 34935 17434 34959 17436
rect 35015 17434 35021 17436
rect 34775 17382 34777 17434
rect 34957 17382 34959 17434
rect 34713 17380 34719 17382
rect 34775 17380 34799 17382
rect 34855 17380 34879 17382
rect 34935 17380 34959 17382
rect 35015 17380 35021 17382
rect 34713 17371 35021 17380
rect 30493 16892 30801 16901
rect 30493 16890 30499 16892
rect 30555 16890 30579 16892
rect 30635 16890 30659 16892
rect 30715 16890 30739 16892
rect 30795 16890 30801 16892
rect 30555 16838 30557 16890
rect 30737 16838 30739 16890
rect 30493 16836 30499 16838
rect 30555 16836 30579 16838
rect 30635 16836 30659 16838
rect 30715 16836 30739 16838
rect 30795 16836 30801 16838
rect 30493 16827 30801 16836
rect 26272 16348 26580 16357
rect 26272 16346 26278 16348
rect 26334 16346 26358 16348
rect 26414 16346 26438 16348
rect 26494 16346 26518 16348
rect 26574 16346 26580 16348
rect 26334 16294 26336 16346
rect 26516 16294 26518 16346
rect 26272 16292 26278 16294
rect 26334 16292 26358 16294
rect 26414 16292 26438 16294
rect 26494 16292 26518 16294
rect 26574 16292 26580 16294
rect 26272 16283 26580 16292
rect 34713 16348 35021 16357
rect 34713 16346 34719 16348
rect 34775 16346 34799 16348
rect 34855 16346 34879 16348
rect 34935 16346 34959 16348
rect 35015 16346 35021 16348
rect 34775 16294 34777 16346
rect 34957 16294 34959 16346
rect 34713 16292 34719 16294
rect 34775 16292 34799 16294
rect 34855 16292 34879 16294
rect 34935 16292 34959 16294
rect 35015 16292 35021 16294
rect 34713 16283 35021 16292
rect 30493 15804 30801 15813
rect 30493 15802 30499 15804
rect 30555 15802 30579 15804
rect 30635 15802 30659 15804
rect 30715 15802 30739 15804
rect 30795 15802 30801 15804
rect 30555 15750 30557 15802
rect 30737 15750 30739 15802
rect 30493 15748 30499 15750
rect 30555 15748 30579 15750
rect 30635 15748 30659 15750
rect 30715 15748 30739 15750
rect 30795 15748 30801 15750
rect 30493 15739 30801 15748
rect 26272 15260 26580 15269
rect 26272 15258 26278 15260
rect 26334 15258 26358 15260
rect 26414 15258 26438 15260
rect 26494 15258 26518 15260
rect 26574 15258 26580 15260
rect 26334 15206 26336 15258
rect 26516 15206 26518 15258
rect 26272 15204 26278 15206
rect 26334 15204 26358 15206
rect 26414 15204 26438 15206
rect 26494 15204 26518 15206
rect 26574 15204 26580 15206
rect 26272 15195 26580 15204
rect 34713 15260 35021 15269
rect 34713 15258 34719 15260
rect 34775 15258 34799 15260
rect 34855 15258 34879 15260
rect 34935 15258 34959 15260
rect 35015 15258 35021 15260
rect 34775 15206 34777 15258
rect 34957 15206 34959 15258
rect 34713 15204 34719 15206
rect 34775 15204 34799 15206
rect 34855 15204 34879 15206
rect 34935 15204 34959 15206
rect 35015 15204 35021 15206
rect 34713 15195 35021 15204
rect 30493 14716 30801 14725
rect 30493 14714 30499 14716
rect 30555 14714 30579 14716
rect 30635 14714 30659 14716
rect 30715 14714 30739 14716
rect 30795 14714 30801 14716
rect 30555 14662 30557 14714
rect 30737 14662 30739 14714
rect 30493 14660 30499 14662
rect 30555 14660 30579 14662
rect 30635 14660 30659 14662
rect 30715 14660 30739 14662
rect 30795 14660 30801 14662
rect 30493 14651 30801 14660
rect 26272 14172 26580 14181
rect 26272 14170 26278 14172
rect 26334 14170 26358 14172
rect 26414 14170 26438 14172
rect 26494 14170 26518 14172
rect 26574 14170 26580 14172
rect 26334 14118 26336 14170
rect 26516 14118 26518 14170
rect 26272 14116 26278 14118
rect 26334 14116 26358 14118
rect 26414 14116 26438 14118
rect 26494 14116 26518 14118
rect 26574 14116 26580 14118
rect 26272 14107 26580 14116
rect 34713 14172 35021 14181
rect 34713 14170 34719 14172
rect 34775 14170 34799 14172
rect 34855 14170 34879 14172
rect 34935 14170 34959 14172
rect 35015 14170 35021 14172
rect 34775 14118 34777 14170
rect 34957 14118 34959 14170
rect 34713 14116 34719 14118
rect 34775 14116 34799 14118
rect 34855 14116 34879 14118
rect 34935 14116 34959 14118
rect 35015 14116 35021 14118
rect 34713 14107 35021 14116
rect 30493 13628 30801 13637
rect 30493 13626 30499 13628
rect 30555 13626 30579 13628
rect 30635 13626 30659 13628
rect 30715 13626 30739 13628
rect 30795 13626 30801 13628
rect 30555 13574 30557 13626
rect 30737 13574 30739 13626
rect 30493 13572 30499 13574
rect 30555 13572 30579 13574
rect 30635 13572 30659 13574
rect 30715 13572 30739 13574
rect 30795 13572 30801 13574
rect 30493 13563 30801 13572
rect 24032 13184 24084 13190
rect 24032 13126 24084 13132
rect 35164 13184 35216 13190
rect 35164 13126 35216 13132
rect 26272 13084 26580 13093
rect 26272 13082 26278 13084
rect 26334 13082 26358 13084
rect 26414 13082 26438 13084
rect 26494 13082 26518 13084
rect 26574 13082 26580 13084
rect 26334 13030 26336 13082
rect 26516 13030 26518 13082
rect 26272 13028 26278 13030
rect 26334 13028 26358 13030
rect 26414 13028 26438 13030
rect 26494 13028 26518 13030
rect 26574 13028 26580 13030
rect 26272 13019 26580 13028
rect 34713 13084 35021 13093
rect 34713 13082 34719 13084
rect 34775 13082 34799 13084
rect 34855 13082 34879 13084
rect 34935 13082 34959 13084
rect 35015 13082 35021 13084
rect 34775 13030 34777 13082
rect 34957 13030 34959 13082
rect 34713 13028 34719 13030
rect 34775 13028 34799 13030
rect 34855 13028 34879 13030
rect 34935 13028 34959 13030
rect 35015 13028 35021 13030
rect 34713 13019 35021 13028
rect 35176 13025 35204 13126
rect 35162 13016 35218 13025
rect 35162 12951 35218 12960
rect 22052 12540 22360 12549
rect 22052 12538 22058 12540
rect 22114 12538 22138 12540
rect 22194 12538 22218 12540
rect 22274 12538 22298 12540
rect 22354 12538 22360 12540
rect 22114 12486 22116 12538
rect 22296 12486 22298 12538
rect 22052 12484 22058 12486
rect 22114 12484 22138 12486
rect 22194 12484 22218 12486
rect 22274 12484 22298 12486
rect 22354 12484 22360 12486
rect 22052 12475 22360 12484
rect 30493 12540 30801 12549
rect 30493 12538 30499 12540
rect 30555 12538 30579 12540
rect 30635 12538 30659 12540
rect 30715 12538 30739 12540
rect 30795 12538 30801 12540
rect 30555 12486 30557 12538
rect 30737 12486 30739 12538
rect 30493 12484 30499 12486
rect 30555 12484 30579 12486
rect 30635 12484 30659 12486
rect 30715 12484 30739 12486
rect 30795 12484 30801 12486
rect 30493 12475 30801 12484
rect 20180 12406 20300 12434
rect 9390 11996 9698 12005
rect 9390 11994 9396 11996
rect 9452 11994 9476 11996
rect 9532 11994 9556 11996
rect 9612 11994 9636 11996
rect 9692 11994 9698 11996
rect 9452 11942 9454 11994
rect 9634 11942 9636 11994
rect 9390 11940 9396 11942
rect 9452 11940 9476 11942
rect 9532 11940 9556 11942
rect 9612 11940 9636 11942
rect 9692 11940 9698 11942
rect 9390 11931 9698 11940
rect 17831 11996 18139 12005
rect 17831 11994 17837 11996
rect 17893 11994 17917 11996
rect 17973 11994 17997 11996
rect 18053 11994 18077 11996
rect 18133 11994 18139 11996
rect 17893 11942 17895 11994
rect 18075 11942 18077 11994
rect 17831 11940 17837 11942
rect 17893 11940 17917 11942
rect 17973 11940 17997 11942
rect 18053 11940 18077 11942
rect 18133 11940 18139 11942
rect 17831 11931 18139 11940
rect 5170 11452 5478 11461
rect 5170 11450 5176 11452
rect 5232 11450 5256 11452
rect 5312 11450 5336 11452
rect 5392 11450 5416 11452
rect 5472 11450 5478 11452
rect 5232 11398 5234 11450
rect 5414 11398 5416 11450
rect 5170 11396 5176 11398
rect 5232 11396 5256 11398
rect 5312 11396 5336 11398
rect 5392 11396 5416 11398
rect 5472 11396 5478 11398
rect 5170 11387 5478 11396
rect 13611 11452 13919 11461
rect 13611 11450 13617 11452
rect 13673 11450 13697 11452
rect 13753 11450 13777 11452
rect 13833 11450 13857 11452
rect 13913 11450 13919 11452
rect 13673 11398 13675 11450
rect 13855 11398 13857 11450
rect 13611 11396 13617 11398
rect 13673 11396 13697 11398
rect 13753 11396 13777 11398
rect 13833 11396 13857 11398
rect 13913 11396 13919 11398
rect 13611 11387 13919 11396
rect 9390 10908 9698 10917
rect 9390 10906 9396 10908
rect 9452 10906 9476 10908
rect 9532 10906 9556 10908
rect 9612 10906 9636 10908
rect 9692 10906 9698 10908
rect 9452 10854 9454 10906
rect 9634 10854 9636 10906
rect 9390 10852 9396 10854
rect 9452 10852 9476 10854
rect 9532 10852 9556 10854
rect 9612 10852 9636 10854
rect 9692 10852 9698 10854
rect 9390 10843 9698 10852
rect 17831 10908 18139 10917
rect 17831 10906 17837 10908
rect 17893 10906 17917 10908
rect 17973 10906 17997 10908
rect 18053 10906 18077 10908
rect 18133 10906 18139 10908
rect 17893 10854 17895 10906
rect 18075 10854 18077 10906
rect 17831 10852 17837 10854
rect 17893 10852 17917 10854
rect 17973 10852 17997 10854
rect 18053 10852 18077 10854
rect 18133 10852 18139 10854
rect 17831 10843 18139 10852
rect 5170 10364 5478 10373
rect 5170 10362 5176 10364
rect 5232 10362 5256 10364
rect 5312 10362 5336 10364
rect 5392 10362 5416 10364
rect 5472 10362 5478 10364
rect 5232 10310 5234 10362
rect 5414 10310 5416 10362
rect 5170 10308 5176 10310
rect 5232 10308 5256 10310
rect 5312 10308 5336 10310
rect 5392 10308 5416 10310
rect 5472 10308 5478 10310
rect 5170 10299 5478 10308
rect 13611 10364 13919 10373
rect 13611 10362 13617 10364
rect 13673 10362 13697 10364
rect 13753 10362 13777 10364
rect 13833 10362 13857 10364
rect 13913 10362 13919 10364
rect 13673 10310 13675 10362
rect 13855 10310 13857 10362
rect 13611 10308 13617 10310
rect 13673 10308 13697 10310
rect 13753 10308 13777 10310
rect 13833 10308 13857 10310
rect 13913 10308 13919 10310
rect 13611 10299 13919 10308
rect 9390 9820 9698 9829
rect 9390 9818 9396 9820
rect 9452 9818 9476 9820
rect 9532 9818 9556 9820
rect 9612 9818 9636 9820
rect 9692 9818 9698 9820
rect 9452 9766 9454 9818
rect 9634 9766 9636 9818
rect 9390 9764 9396 9766
rect 9452 9764 9476 9766
rect 9532 9764 9556 9766
rect 9612 9764 9636 9766
rect 9692 9764 9698 9766
rect 9390 9755 9698 9764
rect 17831 9820 18139 9829
rect 17831 9818 17837 9820
rect 17893 9818 17917 9820
rect 17973 9818 17997 9820
rect 18053 9818 18077 9820
rect 18133 9818 18139 9820
rect 17893 9766 17895 9818
rect 18075 9766 18077 9818
rect 17831 9764 17837 9766
rect 17893 9764 17917 9766
rect 17973 9764 17997 9766
rect 18053 9764 18077 9766
rect 18133 9764 18139 9766
rect 17831 9755 18139 9764
rect 5170 9276 5478 9285
rect 5170 9274 5176 9276
rect 5232 9274 5256 9276
rect 5312 9274 5336 9276
rect 5392 9274 5416 9276
rect 5472 9274 5478 9276
rect 5232 9222 5234 9274
rect 5414 9222 5416 9274
rect 5170 9220 5176 9222
rect 5232 9220 5256 9222
rect 5312 9220 5336 9222
rect 5392 9220 5416 9222
rect 5472 9220 5478 9222
rect 5170 9211 5478 9220
rect 13611 9276 13919 9285
rect 13611 9274 13617 9276
rect 13673 9274 13697 9276
rect 13753 9274 13777 9276
rect 13833 9274 13857 9276
rect 13913 9274 13919 9276
rect 13673 9222 13675 9274
rect 13855 9222 13857 9274
rect 13611 9220 13617 9222
rect 13673 9220 13697 9222
rect 13753 9220 13777 9222
rect 13833 9220 13857 9222
rect 13913 9220 13919 9222
rect 13611 9211 13919 9220
rect 9390 8732 9698 8741
rect 9390 8730 9396 8732
rect 9452 8730 9476 8732
rect 9532 8730 9556 8732
rect 9612 8730 9636 8732
rect 9692 8730 9698 8732
rect 9452 8678 9454 8730
rect 9634 8678 9636 8730
rect 9390 8676 9396 8678
rect 9452 8676 9476 8678
rect 9532 8676 9556 8678
rect 9612 8676 9636 8678
rect 9692 8676 9698 8678
rect 9390 8667 9698 8676
rect 17831 8732 18139 8741
rect 17831 8730 17837 8732
rect 17893 8730 17917 8732
rect 17973 8730 17997 8732
rect 18053 8730 18077 8732
rect 18133 8730 18139 8732
rect 17893 8678 17895 8730
rect 18075 8678 18077 8730
rect 17831 8676 17837 8678
rect 17893 8676 17917 8678
rect 17973 8676 17997 8678
rect 18053 8676 18077 8678
rect 18133 8676 18139 8678
rect 17831 8667 18139 8676
rect 5170 8188 5478 8197
rect 5170 8186 5176 8188
rect 5232 8186 5256 8188
rect 5312 8186 5336 8188
rect 5392 8186 5416 8188
rect 5472 8186 5478 8188
rect 5232 8134 5234 8186
rect 5414 8134 5416 8186
rect 5170 8132 5176 8134
rect 5232 8132 5256 8134
rect 5312 8132 5336 8134
rect 5392 8132 5416 8134
rect 5472 8132 5478 8134
rect 5170 8123 5478 8132
rect 13611 8188 13919 8197
rect 13611 8186 13617 8188
rect 13673 8186 13697 8188
rect 13753 8186 13777 8188
rect 13833 8186 13857 8188
rect 13913 8186 13919 8188
rect 13673 8134 13675 8186
rect 13855 8134 13857 8186
rect 13611 8132 13617 8134
rect 13673 8132 13697 8134
rect 13753 8132 13777 8134
rect 13833 8132 13857 8134
rect 13913 8132 13919 8134
rect 13611 8123 13919 8132
rect 9390 7644 9698 7653
rect 9390 7642 9396 7644
rect 9452 7642 9476 7644
rect 9532 7642 9556 7644
rect 9612 7642 9636 7644
rect 9692 7642 9698 7644
rect 9452 7590 9454 7642
rect 9634 7590 9636 7642
rect 9390 7588 9396 7590
rect 9452 7588 9476 7590
rect 9532 7588 9556 7590
rect 9612 7588 9636 7590
rect 9692 7588 9698 7590
rect 9390 7579 9698 7588
rect 17831 7644 18139 7653
rect 17831 7642 17837 7644
rect 17893 7642 17917 7644
rect 17973 7642 17997 7644
rect 18053 7642 18077 7644
rect 18133 7642 18139 7644
rect 17893 7590 17895 7642
rect 18075 7590 18077 7642
rect 17831 7588 17837 7590
rect 17893 7588 17917 7590
rect 17973 7588 17997 7590
rect 18053 7588 18077 7590
rect 18133 7588 18139 7590
rect 17831 7579 18139 7588
rect 1400 7200 1452 7206
rect 1400 7142 1452 7148
rect 1412 6905 1440 7142
rect 5170 7100 5478 7109
rect 5170 7098 5176 7100
rect 5232 7098 5256 7100
rect 5312 7098 5336 7100
rect 5392 7098 5416 7100
rect 5472 7098 5478 7100
rect 5232 7046 5234 7098
rect 5414 7046 5416 7098
rect 5170 7044 5176 7046
rect 5232 7044 5256 7046
rect 5312 7044 5336 7046
rect 5392 7044 5416 7046
rect 5472 7044 5478 7046
rect 5170 7035 5478 7044
rect 13611 7100 13919 7109
rect 13611 7098 13617 7100
rect 13673 7098 13697 7100
rect 13753 7098 13777 7100
rect 13833 7098 13857 7100
rect 13913 7098 13919 7100
rect 13673 7046 13675 7098
rect 13855 7046 13857 7098
rect 13611 7044 13617 7046
rect 13673 7044 13697 7046
rect 13753 7044 13777 7046
rect 13833 7044 13857 7046
rect 13913 7044 13919 7046
rect 13611 7035 13919 7044
rect 1398 6896 1454 6905
rect 1398 6831 1454 6840
rect 9390 6556 9698 6565
rect 9390 6554 9396 6556
rect 9452 6554 9476 6556
rect 9532 6554 9556 6556
rect 9612 6554 9636 6556
rect 9692 6554 9698 6556
rect 9452 6502 9454 6554
rect 9634 6502 9636 6554
rect 9390 6500 9396 6502
rect 9452 6500 9476 6502
rect 9532 6500 9556 6502
rect 9612 6500 9636 6502
rect 9692 6500 9698 6502
rect 9390 6491 9698 6500
rect 17831 6556 18139 6565
rect 17831 6554 17837 6556
rect 17893 6554 17917 6556
rect 17973 6554 17997 6556
rect 18053 6554 18077 6556
rect 18133 6554 18139 6556
rect 17893 6502 17895 6554
rect 18075 6502 18077 6554
rect 17831 6500 17837 6502
rect 17893 6500 17917 6502
rect 17973 6500 17997 6502
rect 18053 6500 18077 6502
rect 18133 6500 18139 6502
rect 17831 6491 18139 6500
rect 5170 6012 5478 6021
rect 5170 6010 5176 6012
rect 5232 6010 5256 6012
rect 5312 6010 5336 6012
rect 5392 6010 5416 6012
rect 5472 6010 5478 6012
rect 5232 5958 5234 6010
rect 5414 5958 5416 6010
rect 5170 5956 5176 5958
rect 5232 5956 5256 5958
rect 5312 5956 5336 5958
rect 5392 5956 5416 5958
rect 5472 5956 5478 5958
rect 5170 5947 5478 5956
rect 13611 6012 13919 6021
rect 13611 6010 13617 6012
rect 13673 6010 13697 6012
rect 13753 6010 13777 6012
rect 13833 6010 13857 6012
rect 13913 6010 13919 6012
rect 13673 5958 13675 6010
rect 13855 5958 13857 6010
rect 13611 5956 13617 5958
rect 13673 5956 13697 5958
rect 13753 5956 13777 5958
rect 13833 5956 13857 5958
rect 13913 5956 13919 5958
rect 13611 5947 13919 5956
rect 9390 5468 9698 5477
rect 9390 5466 9396 5468
rect 9452 5466 9476 5468
rect 9532 5466 9556 5468
rect 9612 5466 9636 5468
rect 9692 5466 9698 5468
rect 9452 5414 9454 5466
rect 9634 5414 9636 5466
rect 9390 5412 9396 5414
rect 9452 5412 9476 5414
rect 9532 5412 9556 5414
rect 9612 5412 9636 5414
rect 9692 5412 9698 5414
rect 9390 5403 9698 5412
rect 17831 5468 18139 5477
rect 17831 5466 17837 5468
rect 17893 5466 17917 5468
rect 17973 5466 17997 5468
rect 18053 5466 18077 5468
rect 18133 5466 18139 5468
rect 17893 5414 17895 5466
rect 18075 5414 18077 5466
rect 17831 5412 17837 5414
rect 17893 5412 17917 5414
rect 17973 5412 17997 5414
rect 18053 5412 18077 5414
rect 18133 5412 18139 5414
rect 17831 5403 18139 5412
rect 5170 4924 5478 4933
rect 5170 4922 5176 4924
rect 5232 4922 5256 4924
rect 5312 4922 5336 4924
rect 5392 4922 5416 4924
rect 5472 4922 5478 4924
rect 5232 4870 5234 4922
rect 5414 4870 5416 4922
rect 5170 4868 5176 4870
rect 5232 4868 5256 4870
rect 5312 4868 5336 4870
rect 5392 4868 5416 4870
rect 5472 4868 5478 4870
rect 5170 4859 5478 4868
rect 13611 4924 13919 4933
rect 13611 4922 13617 4924
rect 13673 4922 13697 4924
rect 13753 4922 13777 4924
rect 13833 4922 13857 4924
rect 13913 4922 13919 4924
rect 13673 4870 13675 4922
rect 13855 4870 13857 4922
rect 13611 4868 13617 4870
rect 13673 4868 13697 4870
rect 13753 4868 13777 4870
rect 13833 4868 13857 4870
rect 13913 4868 13919 4870
rect 13611 4859 13919 4868
rect 9390 4380 9698 4389
rect 9390 4378 9396 4380
rect 9452 4378 9476 4380
rect 9532 4378 9556 4380
rect 9612 4378 9636 4380
rect 9692 4378 9698 4380
rect 9452 4326 9454 4378
rect 9634 4326 9636 4378
rect 9390 4324 9396 4326
rect 9452 4324 9476 4326
rect 9532 4324 9556 4326
rect 9612 4324 9636 4326
rect 9692 4324 9698 4326
rect 9390 4315 9698 4324
rect 17831 4380 18139 4389
rect 17831 4378 17837 4380
rect 17893 4378 17917 4380
rect 17973 4378 17997 4380
rect 18053 4378 18077 4380
rect 18133 4378 18139 4380
rect 17893 4326 17895 4378
rect 18075 4326 18077 4378
rect 17831 4324 17837 4326
rect 17893 4324 17917 4326
rect 17973 4324 17997 4326
rect 18053 4324 18077 4326
rect 18133 4324 18139 4326
rect 17831 4315 18139 4324
rect 5170 3836 5478 3845
rect 5170 3834 5176 3836
rect 5232 3834 5256 3836
rect 5312 3834 5336 3836
rect 5392 3834 5416 3836
rect 5472 3834 5478 3836
rect 5232 3782 5234 3834
rect 5414 3782 5416 3834
rect 5170 3780 5176 3782
rect 5232 3780 5256 3782
rect 5312 3780 5336 3782
rect 5392 3780 5416 3782
rect 5472 3780 5478 3782
rect 5170 3771 5478 3780
rect 13611 3836 13919 3845
rect 13611 3834 13617 3836
rect 13673 3834 13697 3836
rect 13753 3834 13777 3836
rect 13833 3834 13857 3836
rect 13913 3834 13919 3836
rect 13673 3782 13675 3834
rect 13855 3782 13857 3834
rect 13611 3780 13617 3782
rect 13673 3780 13697 3782
rect 13753 3780 13777 3782
rect 13833 3780 13857 3782
rect 13913 3780 13919 3782
rect 13611 3771 13919 3780
rect 9390 3292 9698 3301
rect 9390 3290 9396 3292
rect 9452 3290 9476 3292
rect 9532 3290 9556 3292
rect 9612 3290 9636 3292
rect 9692 3290 9698 3292
rect 9452 3238 9454 3290
rect 9634 3238 9636 3290
rect 9390 3236 9396 3238
rect 9452 3236 9476 3238
rect 9532 3236 9556 3238
rect 9612 3236 9636 3238
rect 9692 3236 9698 3238
rect 9390 3227 9698 3236
rect 17831 3292 18139 3301
rect 17831 3290 17837 3292
rect 17893 3290 17917 3292
rect 17973 3290 17997 3292
rect 18053 3290 18077 3292
rect 18133 3290 18139 3292
rect 17893 3238 17895 3290
rect 18075 3238 18077 3290
rect 17831 3236 17837 3238
rect 17893 3236 17917 3238
rect 17973 3236 17997 3238
rect 18053 3236 18077 3238
rect 18133 3236 18139 3238
rect 17831 3227 18139 3236
rect 5170 2748 5478 2757
rect 5170 2746 5176 2748
rect 5232 2746 5256 2748
rect 5312 2746 5336 2748
rect 5392 2746 5416 2748
rect 5472 2746 5478 2748
rect 5232 2694 5234 2746
rect 5414 2694 5416 2746
rect 5170 2692 5176 2694
rect 5232 2692 5256 2694
rect 5312 2692 5336 2694
rect 5392 2692 5416 2694
rect 5472 2692 5478 2694
rect 5170 2683 5478 2692
rect 13611 2748 13919 2757
rect 13611 2746 13617 2748
rect 13673 2746 13697 2748
rect 13753 2746 13777 2748
rect 13833 2746 13857 2748
rect 13913 2746 13919 2748
rect 13673 2694 13675 2746
rect 13855 2694 13857 2746
rect 13611 2692 13617 2694
rect 13673 2692 13697 2694
rect 13753 2692 13777 2694
rect 13833 2692 13857 2694
rect 13913 2692 13919 2694
rect 13611 2683 13919 2692
rect 20272 2446 20300 12406
rect 26272 11996 26580 12005
rect 26272 11994 26278 11996
rect 26334 11994 26358 11996
rect 26414 11994 26438 11996
rect 26494 11994 26518 11996
rect 26574 11994 26580 11996
rect 26334 11942 26336 11994
rect 26516 11942 26518 11994
rect 26272 11940 26278 11942
rect 26334 11940 26358 11942
rect 26414 11940 26438 11942
rect 26494 11940 26518 11942
rect 26574 11940 26580 11942
rect 26272 11931 26580 11940
rect 34713 11996 35021 12005
rect 34713 11994 34719 11996
rect 34775 11994 34799 11996
rect 34855 11994 34879 11996
rect 34935 11994 34959 11996
rect 35015 11994 35021 11996
rect 34775 11942 34777 11994
rect 34957 11942 34959 11994
rect 34713 11940 34719 11942
rect 34775 11940 34799 11942
rect 34855 11940 34879 11942
rect 34935 11940 34959 11942
rect 35015 11940 35021 11942
rect 34713 11931 35021 11940
rect 22052 11452 22360 11461
rect 22052 11450 22058 11452
rect 22114 11450 22138 11452
rect 22194 11450 22218 11452
rect 22274 11450 22298 11452
rect 22354 11450 22360 11452
rect 22114 11398 22116 11450
rect 22296 11398 22298 11450
rect 22052 11396 22058 11398
rect 22114 11396 22138 11398
rect 22194 11396 22218 11398
rect 22274 11396 22298 11398
rect 22354 11396 22360 11398
rect 22052 11387 22360 11396
rect 30493 11452 30801 11461
rect 30493 11450 30499 11452
rect 30555 11450 30579 11452
rect 30635 11450 30659 11452
rect 30715 11450 30739 11452
rect 30795 11450 30801 11452
rect 30555 11398 30557 11450
rect 30737 11398 30739 11450
rect 30493 11396 30499 11398
rect 30555 11396 30579 11398
rect 30635 11396 30659 11398
rect 30715 11396 30739 11398
rect 30795 11396 30801 11398
rect 30493 11387 30801 11396
rect 26272 10908 26580 10917
rect 26272 10906 26278 10908
rect 26334 10906 26358 10908
rect 26414 10906 26438 10908
rect 26494 10906 26518 10908
rect 26574 10906 26580 10908
rect 26334 10854 26336 10906
rect 26516 10854 26518 10906
rect 26272 10852 26278 10854
rect 26334 10852 26358 10854
rect 26414 10852 26438 10854
rect 26494 10852 26518 10854
rect 26574 10852 26580 10854
rect 26272 10843 26580 10852
rect 34713 10908 35021 10917
rect 34713 10906 34719 10908
rect 34775 10906 34799 10908
rect 34855 10906 34879 10908
rect 34935 10906 34959 10908
rect 35015 10906 35021 10908
rect 34775 10854 34777 10906
rect 34957 10854 34959 10906
rect 34713 10852 34719 10854
rect 34775 10852 34799 10854
rect 34855 10852 34879 10854
rect 34935 10852 34959 10854
rect 35015 10852 35021 10854
rect 34713 10843 35021 10852
rect 22052 10364 22360 10373
rect 22052 10362 22058 10364
rect 22114 10362 22138 10364
rect 22194 10362 22218 10364
rect 22274 10362 22298 10364
rect 22354 10362 22360 10364
rect 22114 10310 22116 10362
rect 22296 10310 22298 10362
rect 22052 10308 22058 10310
rect 22114 10308 22138 10310
rect 22194 10308 22218 10310
rect 22274 10308 22298 10310
rect 22354 10308 22360 10310
rect 22052 10299 22360 10308
rect 30493 10364 30801 10373
rect 30493 10362 30499 10364
rect 30555 10362 30579 10364
rect 30635 10362 30659 10364
rect 30715 10362 30739 10364
rect 30795 10362 30801 10364
rect 30555 10310 30557 10362
rect 30737 10310 30739 10362
rect 30493 10308 30499 10310
rect 30555 10308 30579 10310
rect 30635 10308 30659 10310
rect 30715 10308 30739 10310
rect 30795 10308 30801 10310
rect 30493 10299 30801 10308
rect 26272 9820 26580 9829
rect 26272 9818 26278 9820
rect 26334 9818 26358 9820
rect 26414 9818 26438 9820
rect 26494 9818 26518 9820
rect 26574 9818 26580 9820
rect 26334 9766 26336 9818
rect 26516 9766 26518 9818
rect 26272 9764 26278 9766
rect 26334 9764 26358 9766
rect 26414 9764 26438 9766
rect 26494 9764 26518 9766
rect 26574 9764 26580 9766
rect 26272 9755 26580 9764
rect 34713 9820 35021 9829
rect 34713 9818 34719 9820
rect 34775 9818 34799 9820
rect 34855 9818 34879 9820
rect 34935 9818 34959 9820
rect 35015 9818 35021 9820
rect 34775 9766 34777 9818
rect 34957 9766 34959 9818
rect 34713 9764 34719 9766
rect 34775 9764 34799 9766
rect 34855 9764 34879 9766
rect 34935 9764 34959 9766
rect 35015 9764 35021 9766
rect 34713 9755 35021 9764
rect 22052 9276 22360 9285
rect 22052 9274 22058 9276
rect 22114 9274 22138 9276
rect 22194 9274 22218 9276
rect 22274 9274 22298 9276
rect 22354 9274 22360 9276
rect 22114 9222 22116 9274
rect 22296 9222 22298 9274
rect 22052 9220 22058 9222
rect 22114 9220 22138 9222
rect 22194 9220 22218 9222
rect 22274 9220 22298 9222
rect 22354 9220 22360 9222
rect 22052 9211 22360 9220
rect 30493 9276 30801 9285
rect 30493 9274 30499 9276
rect 30555 9274 30579 9276
rect 30635 9274 30659 9276
rect 30715 9274 30739 9276
rect 30795 9274 30801 9276
rect 30555 9222 30557 9274
rect 30737 9222 30739 9274
rect 30493 9220 30499 9222
rect 30555 9220 30579 9222
rect 30635 9220 30659 9222
rect 30715 9220 30739 9222
rect 30795 9220 30801 9222
rect 30493 9211 30801 9220
rect 26272 8732 26580 8741
rect 26272 8730 26278 8732
rect 26334 8730 26358 8732
rect 26414 8730 26438 8732
rect 26494 8730 26518 8732
rect 26574 8730 26580 8732
rect 26334 8678 26336 8730
rect 26516 8678 26518 8730
rect 26272 8676 26278 8678
rect 26334 8676 26358 8678
rect 26414 8676 26438 8678
rect 26494 8676 26518 8678
rect 26574 8676 26580 8678
rect 26272 8667 26580 8676
rect 34713 8732 35021 8741
rect 34713 8730 34719 8732
rect 34775 8730 34799 8732
rect 34855 8730 34879 8732
rect 34935 8730 34959 8732
rect 35015 8730 35021 8732
rect 34775 8678 34777 8730
rect 34957 8678 34959 8730
rect 34713 8676 34719 8678
rect 34775 8676 34799 8678
rect 34855 8676 34879 8678
rect 34935 8676 34959 8678
rect 35015 8676 35021 8678
rect 34713 8667 35021 8676
rect 22052 8188 22360 8197
rect 22052 8186 22058 8188
rect 22114 8186 22138 8188
rect 22194 8186 22218 8188
rect 22274 8186 22298 8188
rect 22354 8186 22360 8188
rect 22114 8134 22116 8186
rect 22296 8134 22298 8186
rect 22052 8132 22058 8134
rect 22114 8132 22138 8134
rect 22194 8132 22218 8134
rect 22274 8132 22298 8134
rect 22354 8132 22360 8134
rect 22052 8123 22360 8132
rect 30493 8188 30801 8197
rect 30493 8186 30499 8188
rect 30555 8186 30579 8188
rect 30635 8186 30659 8188
rect 30715 8186 30739 8188
rect 30795 8186 30801 8188
rect 30555 8134 30557 8186
rect 30737 8134 30739 8186
rect 30493 8132 30499 8134
rect 30555 8132 30579 8134
rect 30635 8132 30659 8134
rect 30715 8132 30739 8134
rect 30795 8132 30801 8134
rect 30493 8123 30801 8132
rect 26272 7644 26580 7653
rect 26272 7642 26278 7644
rect 26334 7642 26358 7644
rect 26414 7642 26438 7644
rect 26494 7642 26518 7644
rect 26574 7642 26580 7644
rect 26334 7590 26336 7642
rect 26516 7590 26518 7642
rect 26272 7588 26278 7590
rect 26334 7588 26358 7590
rect 26414 7588 26438 7590
rect 26494 7588 26518 7590
rect 26574 7588 26580 7590
rect 26272 7579 26580 7588
rect 34713 7644 35021 7653
rect 34713 7642 34719 7644
rect 34775 7642 34799 7644
rect 34855 7642 34879 7644
rect 34935 7642 34959 7644
rect 35015 7642 35021 7644
rect 34775 7590 34777 7642
rect 34957 7590 34959 7642
rect 34713 7588 34719 7590
rect 34775 7588 34799 7590
rect 34855 7588 34879 7590
rect 34935 7588 34959 7590
rect 35015 7588 35021 7590
rect 34713 7579 35021 7588
rect 22052 7100 22360 7109
rect 22052 7098 22058 7100
rect 22114 7098 22138 7100
rect 22194 7098 22218 7100
rect 22274 7098 22298 7100
rect 22354 7098 22360 7100
rect 22114 7046 22116 7098
rect 22296 7046 22298 7098
rect 22052 7044 22058 7046
rect 22114 7044 22138 7046
rect 22194 7044 22218 7046
rect 22274 7044 22298 7046
rect 22354 7044 22360 7046
rect 22052 7035 22360 7044
rect 30493 7100 30801 7109
rect 30493 7098 30499 7100
rect 30555 7098 30579 7100
rect 30635 7098 30659 7100
rect 30715 7098 30739 7100
rect 30795 7098 30801 7100
rect 30555 7046 30557 7098
rect 30737 7046 30739 7098
rect 30493 7044 30499 7046
rect 30555 7044 30579 7046
rect 30635 7044 30659 7046
rect 30715 7044 30739 7046
rect 30795 7044 30801 7046
rect 30493 7035 30801 7044
rect 26272 6556 26580 6565
rect 26272 6554 26278 6556
rect 26334 6554 26358 6556
rect 26414 6554 26438 6556
rect 26494 6554 26518 6556
rect 26574 6554 26580 6556
rect 26334 6502 26336 6554
rect 26516 6502 26518 6554
rect 26272 6500 26278 6502
rect 26334 6500 26358 6502
rect 26414 6500 26438 6502
rect 26494 6500 26518 6502
rect 26574 6500 26580 6502
rect 26272 6491 26580 6500
rect 34713 6556 35021 6565
rect 34713 6554 34719 6556
rect 34775 6554 34799 6556
rect 34855 6554 34879 6556
rect 34935 6554 34959 6556
rect 35015 6554 35021 6556
rect 34775 6502 34777 6554
rect 34957 6502 34959 6554
rect 34713 6500 34719 6502
rect 34775 6500 34799 6502
rect 34855 6500 34879 6502
rect 34935 6500 34959 6502
rect 35015 6500 35021 6502
rect 34713 6491 35021 6500
rect 22052 6012 22360 6021
rect 22052 6010 22058 6012
rect 22114 6010 22138 6012
rect 22194 6010 22218 6012
rect 22274 6010 22298 6012
rect 22354 6010 22360 6012
rect 22114 5958 22116 6010
rect 22296 5958 22298 6010
rect 22052 5956 22058 5958
rect 22114 5956 22138 5958
rect 22194 5956 22218 5958
rect 22274 5956 22298 5958
rect 22354 5956 22360 5958
rect 22052 5947 22360 5956
rect 30493 6012 30801 6021
rect 30493 6010 30499 6012
rect 30555 6010 30579 6012
rect 30635 6010 30659 6012
rect 30715 6010 30739 6012
rect 30795 6010 30801 6012
rect 30555 5958 30557 6010
rect 30737 5958 30739 6010
rect 30493 5956 30499 5958
rect 30555 5956 30579 5958
rect 30635 5956 30659 5958
rect 30715 5956 30739 5958
rect 30795 5956 30801 5958
rect 30493 5947 30801 5956
rect 34518 5672 34574 5681
rect 34518 5607 34520 5616
rect 34572 5607 34574 5616
rect 34520 5578 34572 5584
rect 26272 5468 26580 5477
rect 26272 5466 26278 5468
rect 26334 5466 26358 5468
rect 26414 5466 26438 5468
rect 26494 5466 26518 5468
rect 26574 5466 26580 5468
rect 26334 5414 26336 5466
rect 26516 5414 26518 5466
rect 26272 5412 26278 5414
rect 26334 5412 26358 5414
rect 26414 5412 26438 5414
rect 26494 5412 26518 5414
rect 26574 5412 26580 5414
rect 26272 5403 26580 5412
rect 34713 5468 35021 5477
rect 34713 5466 34719 5468
rect 34775 5466 34799 5468
rect 34855 5466 34879 5468
rect 34935 5466 34959 5468
rect 35015 5466 35021 5468
rect 34775 5414 34777 5466
rect 34957 5414 34959 5466
rect 34713 5412 34719 5414
rect 34775 5412 34799 5414
rect 34855 5412 34879 5414
rect 34935 5412 34959 5414
rect 35015 5412 35021 5414
rect 34713 5403 35021 5412
rect 22052 4924 22360 4933
rect 22052 4922 22058 4924
rect 22114 4922 22138 4924
rect 22194 4922 22218 4924
rect 22274 4922 22298 4924
rect 22354 4922 22360 4924
rect 22114 4870 22116 4922
rect 22296 4870 22298 4922
rect 22052 4868 22058 4870
rect 22114 4868 22138 4870
rect 22194 4868 22218 4870
rect 22274 4868 22298 4870
rect 22354 4868 22360 4870
rect 22052 4859 22360 4868
rect 30493 4924 30801 4933
rect 30493 4922 30499 4924
rect 30555 4922 30579 4924
rect 30635 4922 30659 4924
rect 30715 4922 30739 4924
rect 30795 4922 30801 4924
rect 30555 4870 30557 4922
rect 30737 4870 30739 4922
rect 30493 4868 30499 4870
rect 30555 4868 30579 4870
rect 30635 4868 30659 4870
rect 30715 4868 30739 4870
rect 30795 4868 30801 4870
rect 30493 4859 30801 4868
rect 26272 4380 26580 4389
rect 26272 4378 26278 4380
rect 26334 4378 26358 4380
rect 26414 4378 26438 4380
rect 26494 4378 26518 4380
rect 26574 4378 26580 4380
rect 26334 4326 26336 4378
rect 26516 4326 26518 4378
rect 26272 4324 26278 4326
rect 26334 4324 26358 4326
rect 26414 4324 26438 4326
rect 26494 4324 26518 4326
rect 26574 4324 26580 4326
rect 26272 4315 26580 4324
rect 34713 4380 35021 4389
rect 34713 4378 34719 4380
rect 34775 4378 34799 4380
rect 34855 4378 34879 4380
rect 34935 4378 34959 4380
rect 35015 4378 35021 4380
rect 34775 4326 34777 4378
rect 34957 4326 34959 4378
rect 34713 4324 34719 4326
rect 34775 4324 34799 4326
rect 34855 4324 34879 4326
rect 34935 4324 34959 4326
rect 35015 4324 35021 4326
rect 34713 4315 35021 4324
rect 22052 3836 22360 3845
rect 22052 3834 22058 3836
rect 22114 3834 22138 3836
rect 22194 3834 22218 3836
rect 22274 3834 22298 3836
rect 22354 3834 22360 3836
rect 22114 3782 22116 3834
rect 22296 3782 22298 3834
rect 22052 3780 22058 3782
rect 22114 3780 22138 3782
rect 22194 3780 22218 3782
rect 22274 3780 22298 3782
rect 22354 3780 22360 3782
rect 22052 3771 22360 3780
rect 30493 3836 30801 3845
rect 30493 3834 30499 3836
rect 30555 3834 30579 3836
rect 30635 3834 30659 3836
rect 30715 3834 30739 3836
rect 30795 3834 30801 3836
rect 30555 3782 30557 3834
rect 30737 3782 30739 3834
rect 30493 3780 30499 3782
rect 30555 3780 30579 3782
rect 30635 3780 30659 3782
rect 30715 3780 30739 3782
rect 30795 3780 30801 3782
rect 30493 3771 30801 3780
rect 26272 3292 26580 3301
rect 26272 3290 26278 3292
rect 26334 3290 26358 3292
rect 26414 3290 26438 3292
rect 26494 3290 26518 3292
rect 26574 3290 26580 3292
rect 26334 3238 26336 3290
rect 26516 3238 26518 3290
rect 26272 3236 26278 3238
rect 26334 3236 26358 3238
rect 26414 3236 26438 3238
rect 26494 3236 26518 3238
rect 26574 3236 26580 3238
rect 26272 3227 26580 3236
rect 34713 3292 35021 3301
rect 34713 3290 34719 3292
rect 34775 3290 34799 3292
rect 34855 3290 34879 3292
rect 34935 3290 34959 3292
rect 35015 3290 35021 3292
rect 34775 3238 34777 3290
rect 34957 3238 34959 3290
rect 34713 3236 34719 3238
rect 34775 3236 34799 3238
rect 34855 3236 34879 3238
rect 34935 3236 34959 3238
rect 35015 3236 35021 3238
rect 34713 3227 35021 3236
rect 22052 2748 22360 2757
rect 22052 2746 22058 2748
rect 22114 2746 22138 2748
rect 22194 2746 22218 2748
rect 22274 2746 22298 2748
rect 22354 2746 22360 2748
rect 22114 2694 22116 2746
rect 22296 2694 22298 2746
rect 22052 2692 22058 2694
rect 22114 2692 22138 2694
rect 22194 2692 22218 2694
rect 22274 2692 22298 2694
rect 22354 2692 22360 2694
rect 22052 2683 22360 2692
rect 30493 2748 30801 2757
rect 30493 2746 30499 2748
rect 30555 2746 30579 2748
rect 30635 2746 30659 2748
rect 30715 2746 30739 2748
rect 30795 2746 30801 2748
rect 30555 2694 30557 2746
rect 30737 2694 30739 2746
rect 30493 2692 30499 2694
rect 30555 2692 30579 2694
rect 30635 2692 30659 2694
rect 30715 2692 30739 2694
rect 30795 2692 30801 2694
rect 30493 2683 30801 2692
rect 20720 2508 20772 2514
rect 20720 2450 20772 2456
rect 13636 2440 13688 2446
rect 13636 2382 13688 2388
rect 20260 2440 20312 2446
rect 20260 2382 20312 2388
rect 20 2304 72 2310
rect 20 2246 72 2252
rect 6552 2304 6604 2310
rect 6552 2246 6604 2252
rect 32 800 60 2246
rect 6564 1170 6592 2246
rect 9390 2204 9698 2213
rect 9390 2202 9396 2204
rect 9452 2202 9476 2204
rect 9532 2202 9556 2204
rect 9612 2202 9636 2204
rect 9692 2202 9698 2204
rect 9452 2150 9454 2202
rect 9634 2150 9636 2202
rect 9390 2148 9396 2150
rect 9452 2148 9476 2150
rect 9532 2148 9556 2150
rect 9612 2148 9636 2150
rect 9692 2148 9698 2150
rect 9390 2139 9698 2148
rect 13648 1306 13676 2382
rect 17831 2204 18139 2213
rect 17831 2202 17837 2204
rect 17893 2202 17917 2204
rect 17973 2202 17997 2204
rect 18053 2202 18077 2204
rect 18133 2202 18139 2204
rect 17893 2150 17895 2202
rect 18075 2150 18077 2202
rect 17831 2148 17837 2150
rect 17893 2148 17917 2150
rect 17973 2148 17997 2150
rect 18053 2148 18077 2150
rect 18133 2148 18139 2150
rect 17831 2139 18139 2148
rect 20732 1442 20760 2450
rect 27160 2304 27212 2310
rect 27160 2246 27212 2252
rect 34244 2304 34296 2310
rect 34244 2246 34296 2252
rect 26272 2204 26580 2213
rect 26272 2202 26278 2204
rect 26334 2202 26358 2204
rect 26414 2202 26438 2204
rect 26494 2202 26518 2204
rect 26574 2202 26580 2204
rect 26334 2150 26336 2202
rect 26516 2150 26518 2202
rect 26272 2148 26278 2150
rect 26334 2148 26358 2150
rect 26414 2148 26438 2150
rect 26494 2148 26518 2150
rect 26574 2148 26580 2150
rect 26272 2139 26580 2148
rect 6472 1142 6592 1170
rect 13556 1278 13676 1306
rect 20640 1414 20760 1442
rect 6472 800 6500 1142
rect 13556 800 13584 1278
rect 20640 800 20668 1414
rect 27172 1170 27200 2246
rect 34256 1170 34284 2246
rect 34713 2204 35021 2213
rect 34713 2202 34719 2204
rect 34775 2202 34799 2204
rect 34855 2202 34879 2204
rect 34935 2202 34959 2204
rect 35015 2202 35021 2204
rect 34775 2150 34777 2202
rect 34957 2150 34959 2202
rect 34713 2148 34719 2150
rect 34775 2148 34799 2150
rect 34855 2148 34879 2150
rect 34935 2148 34959 2150
rect 35015 2148 35021 2150
rect 34713 2139 35021 2148
rect 27080 1142 27200 1170
rect 34164 1142 34284 1170
rect 27080 800 27108 1142
rect 34164 800 34192 1142
rect -10 0 102 800
rect 6430 0 6542 800
rect 13514 0 13626 800
rect 20598 0 20710 800
rect 27038 0 27150 800
rect 34122 0 34234 800
<< via2 >>
rect 5176 39738 5232 39740
rect 5256 39738 5312 39740
rect 5336 39738 5392 39740
rect 5416 39738 5472 39740
rect 5176 39686 5222 39738
rect 5222 39686 5232 39738
rect 5256 39686 5286 39738
rect 5286 39686 5298 39738
rect 5298 39686 5312 39738
rect 5336 39686 5350 39738
rect 5350 39686 5362 39738
rect 5362 39686 5392 39738
rect 5416 39686 5426 39738
rect 5426 39686 5472 39738
rect 5176 39684 5232 39686
rect 5256 39684 5312 39686
rect 5336 39684 5392 39686
rect 5416 39684 5472 39686
rect 13617 39738 13673 39740
rect 13697 39738 13753 39740
rect 13777 39738 13833 39740
rect 13857 39738 13913 39740
rect 13617 39686 13663 39738
rect 13663 39686 13673 39738
rect 13697 39686 13727 39738
rect 13727 39686 13739 39738
rect 13739 39686 13753 39738
rect 13777 39686 13791 39738
rect 13791 39686 13803 39738
rect 13803 39686 13833 39738
rect 13857 39686 13867 39738
rect 13867 39686 13913 39738
rect 13617 39684 13673 39686
rect 13697 39684 13753 39686
rect 13777 39684 13833 39686
rect 13857 39684 13913 39686
rect 5176 38650 5232 38652
rect 5256 38650 5312 38652
rect 5336 38650 5392 38652
rect 5416 38650 5472 38652
rect 5176 38598 5222 38650
rect 5222 38598 5232 38650
rect 5256 38598 5286 38650
rect 5286 38598 5298 38650
rect 5298 38598 5312 38650
rect 5336 38598 5350 38650
rect 5350 38598 5362 38650
rect 5362 38598 5392 38650
rect 5416 38598 5426 38650
rect 5426 38598 5472 38650
rect 5176 38596 5232 38598
rect 5256 38596 5312 38598
rect 5336 38596 5392 38598
rect 5416 38596 5472 38598
rect 9396 39194 9452 39196
rect 9476 39194 9532 39196
rect 9556 39194 9612 39196
rect 9636 39194 9692 39196
rect 9396 39142 9442 39194
rect 9442 39142 9452 39194
rect 9476 39142 9506 39194
rect 9506 39142 9518 39194
rect 9518 39142 9532 39194
rect 9556 39142 9570 39194
rect 9570 39142 9582 39194
rect 9582 39142 9612 39194
rect 9636 39142 9646 39194
rect 9646 39142 9692 39194
rect 9396 39140 9452 39142
rect 9476 39140 9532 39142
rect 9556 39140 9612 39142
rect 9636 39140 9692 39142
rect 13617 38650 13673 38652
rect 13697 38650 13753 38652
rect 13777 38650 13833 38652
rect 13857 38650 13913 38652
rect 13617 38598 13663 38650
rect 13663 38598 13673 38650
rect 13697 38598 13727 38650
rect 13727 38598 13739 38650
rect 13739 38598 13753 38650
rect 13777 38598 13791 38650
rect 13791 38598 13803 38650
rect 13803 38598 13833 38650
rect 13857 38598 13867 38650
rect 13867 38598 13913 38650
rect 13617 38596 13673 38598
rect 13697 38596 13753 38598
rect 13777 38596 13833 38598
rect 13857 38596 13913 38598
rect 5176 37562 5232 37564
rect 5256 37562 5312 37564
rect 5336 37562 5392 37564
rect 5416 37562 5472 37564
rect 5176 37510 5222 37562
rect 5222 37510 5232 37562
rect 5256 37510 5286 37562
rect 5286 37510 5298 37562
rect 5298 37510 5312 37562
rect 5336 37510 5350 37562
rect 5350 37510 5362 37562
rect 5362 37510 5392 37562
rect 5416 37510 5426 37562
rect 5426 37510 5472 37562
rect 5176 37508 5232 37510
rect 5256 37508 5312 37510
rect 5336 37508 5392 37510
rect 5416 37508 5472 37510
rect 5176 36474 5232 36476
rect 5256 36474 5312 36476
rect 5336 36474 5392 36476
rect 5416 36474 5472 36476
rect 5176 36422 5222 36474
rect 5222 36422 5232 36474
rect 5256 36422 5286 36474
rect 5286 36422 5298 36474
rect 5298 36422 5312 36474
rect 5336 36422 5350 36474
rect 5350 36422 5362 36474
rect 5362 36422 5392 36474
rect 5416 36422 5426 36474
rect 5426 36422 5472 36474
rect 5176 36420 5232 36422
rect 5256 36420 5312 36422
rect 5336 36420 5392 36422
rect 5416 36420 5472 36422
rect 938 36116 940 36136
rect 940 36116 992 36136
rect 992 36116 994 36136
rect 938 36080 994 36116
rect 5176 35386 5232 35388
rect 5256 35386 5312 35388
rect 5336 35386 5392 35388
rect 5416 35386 5472 35388
rect 5176 35334 5222 35386
rect 5222 35334 5232 35386
rect 5256 35334 5286 35386
rect 5286 35334 5298 35386
rect 5298 35334 5312 35386
rect 5336 35334 5350 35386
rect 5350 35334 5362 35386
rect 5362 35334 5392 35386
rect 5416 35334 5426 35386
rect 5426 35334 5472 35386
rect 5176 35332 5232 35334
rect 5256 35332 5312 35334
rect 5336 35332 5392 35334
rect 5416 35332 5472 35334
rect 5176 34298 5232 34300
rect 5256 34298 5312 34300
rect 5336 34298 5392 34300
rect 5416 34298 5472 34300
rect 5176 34246 5222 34298
rect 5222 34246 5232 34298
rect 5256 34246 5286 34298
rect 5286 34246 5298 34298
rect 5298 34246 5312 34298
rect 5336 34246 5350 34298
rect 5350 34246 5362 34298
rect 5362 34246 5392 34298
rect 5416 34246 5426 34298
rect 5426 34246 5472 34298
rect 5176 34244 5232 34246
rect 5256 34244 5312 34246
rect 5336 34244 5392 34246
rect 5416 34244 5472 34246
rect 5176 33210 5232 33212
rect 5256 33210 5312 33212
rect 5336 33210 5392 33212
rect 5416 33210 5472 33212
rect 5176 33158 5222 33210
rect 5222 33158 5232 33210
rect 5256 33158 5286 33210
rect 5286 33158 5298 33210
rect 5298 33158 5312 33210
rect 5336 33158 5350 33210
rect 5350 33158 5362 33210
rect 5362 33158 5392 33210
rect 5416 33158 5426 33210
rect 5426 33158 5472 33210
rect 5176 33156 5232 33158
rect 5256 33156 5312 33158
rect 5336 33156 5392 33158
rect 5416 33156 5472 33158
rect 5176 32122 5232 32124
rect 5256 32122 5312 32124
rect 5336 32122 5392 32124
rect 5416 32122 5472 32124
rect 5176 32070 5222 32122
rect 5222 32070 5232 32122
rect 5256 32070 5286 32122
rect 5286 32070 5298 32122
rect 5298 32070 5312 32122
rect 5336 32070 5350 32122
rect 5350 32070 5362 32122
rect 5362 32070 5392 32122
rect 5416 32070 5426 32122
rect 5426 32070 5472 32122
rect 5176 32068 5232 32070
rect 5256 32068 5312 32070
rect 5336 32068 5392 32070
rect 5416 32068 5472 32070
rect 5176 31034 5232 31036
rect 5256 31034 5312 31036
rect 5336 31034 5392 31036
rect 5416 31034 5472 31036
rect 5176 30982 5222 31034
rect 5222 30982 5232 31034
rect 5256 30982 5286 31034
rect 5286 30982 5298 31034
rect 5298 30982 5312 31034
rect 5336 30982 5350 31034
rect 5350 30982 5362 31034
rect 5362 30982 5392 31034
rect 5416 30982 5426 31034
rect 5426 30982 5472 31034
rect 5176 30980 5232 30982
rect 5256 30980 5312 30982
rect 5336 30980 5392 30982
rect 5416 30980 5472 30982
rect 5176 29946 5232 29948
rect 5256 29946 5312 29948
rect 5336 29946 5392 29948
rect 5416 29946 5472 29948
rect 5176 29894 5222 29946
rect 5222 29894 5232 29946
rect 5256 29894 5286 29946
rect 5286 29894 5298 29946
rect 5298 29894 5312 29946
rect 5336 29894 5350 29946
rect 5350 29894 5362 29946
rect 5362 29894 5392 29946
rect 5416 29894 5426 29946
rect 5426 29894 5472 29946
rect 5176 29892 5232 29894
rect 5256 29892 5312 29894
rect 5336 29892 5392 29894
rect 5416 29892 5472 29894
rect 9396 38106 9452 38108
rect 9476 38106 9532 38108
rect 9556 38106 9612 38108
rect 9636 38106 9692 38108
rect 9396 38054 9442 38106
rect 9442 38054 9452 38106
rect 9476 38054 9506 38106
rect 9506 38054 9518 38106
rect 9518 38054 9532 38106
rect 9556 38054 9570 38106
rect 9570 38054 9582 38106
rect 9582 38054 9612 38106
rect 9636 38054 9646 38106
rect 9646 38054 9692 38106
rect 9396 38052 9452 38054
rect 9476 38052 9532 38054
rect 9556 38052 9612 38054
rect 9636 38052 9692 38054
rect 1398 28872 1454 28928
rect 938 21800 994 21856
rect 5176 28858 5232 28860
rect 5256 28858 5312 28860
rect 5336 28858 5392 28860
rect 5416 28858 5472 28860
rect 5176 28806 5222 28858
rect 5222 28806 5232 28858
rect 5256 28806 5286 28858
rect 5286 28806 5298 28858
rect 5298 28806 5312 28858
rect 5336 28806 5350 28858
rect 5350 28806 5362 28858
rect 5362 28806 5392 28858
rect 5416 28806 5426 28858
rect 5426 28806 5472 28858
rect 5176 28804 5232 28806
rect 5256 28804 5312 28806
rect 5336 28804 5392 28806
rect 5416 28804 5472 28806
rect 5176 27770 5232 27772
rect 5256 27770 5312 27772
rect 5336 27770 5392 27772
rect 5416 27770 5472 27772
rect 5176 27718 5222 27770
rect 5222 27718 5232 27770
rect 5256 27718 5286 27770
rect 5286 27718 5298 27770
rect 5298 27718 5312 27770
rect 5336 27718 5350 27770
rect 5350 27718 5362 27770
rect 5362 27718 5392 27770
rect 5416 27718 5426 27770
rect 5426 27718 5472 27770
rect 5176 27716 5232 27718
rect 5256 27716 5312 27718
rect 5336 27716 5392 27718
rect 5416 27716 5472 27718
rect 5176 26682 5232 26684
rect 5256 26682 5312 26684
rect 5336 26682 5392 26684
rect 5416 26682 5472 26684
rect 5176 26630 5222 26682
rect 5222 26630 5232 26682
rect 5256 26630 5286 26682
rect 5286 26630 5298 26682
rect 5298 26630 5312 26682
rect 5336 26630 5350 26682
rect 5350 26630 5362 26682
rect 5362 26630 5392 26682
rect 5416 26630 5426 26682
rect 5426 26630 5472 26682
rect 5176 26628 5232 26630
rect 5256 26628 5312 26630
rect 5336 26628 5392 26630
rect 5416 26628 5472 26630
rect 5176 25594 5232 25596
rect 5256 25594 5312 25596
rect 5336 25594 5392 25596
rect 5416 25594 5472 25596
rect 5176 25542 5222 25594
rect 5222 25542 5232 25594
rect 5256 25542 5286 25594
rect 5286 25542 5298 25594
rect 5298 25542 5312 25594
rect 5336 25542 5350 25594
rect 5350 25542 5362 25594
rect 5362 25542 5392 25594
rect 5416 25542 5426 25594
rect 5426 25542 5472 25594
rect 5176 25540 5232 25542
rect 5256 25540 5312 25542
rect 5336 25540 5392 25542
rect 5416 25540 5472 25542
rect 5176 24506 5232 24508
rect 5256 24506 5312 24508
rect 5336 24506 5392 24508
rect 5416 24506 5472 24508
rect 5176 24454 5222 24506
rect 5222 24454 5232 24506
rect 5256 24454 5286 24506
rect 5286 24454 5298 24506
rect 5298 24454 5312 24506
rect 5336 24454 5350 24506
rect 5350 24454 5362 24506
rect 5362 24454 5392 24506
rect 5416 24454 5426 24506
rect 5426 24454 5472 24506
rect 5176 24452 5232 24454
rect 5256 24452 5312 24454
rect 5336 24452 5392 24454
rect 5416 24452 5472 24454
rect 5176 23418 5232 23420
rect 5256 23418 5312 23420
rect 5336 23418 5392 23420
rect 5416 23418 5472 23420
rect 5176 23366 5222 23418
rect 5222 23366 5232 23418
rect 5256 23366 5286 23418
rect 5286 23366 5298 23418
rect 5298 23366 5312 23418
rect 5336 23366 5350 23418
rect 5350 23366 5362 23418
rect 5362 23366 5392 23418
rect 5416 23366 5426 23418
rect 5426 23366 5472 23418
rect 5176 23364 5232 23366
rect 5256 23364 5312 23366
rect 5336 23364 5392 23366
rect 5416 23364 5472 23366
rect 5176 22330 5232 22332
rect 5256 22330 5312 22332
rect 5336 22330 5392 22332
rect 5416 22330 5472 22332
rect 5176 22278 5222 22330
rect 5222 22278 5232 22330
rect 5256 22278 5286 22330
rect 5286 22278 5298 22330
rect 5298 22278 5312 22330
rect 5336 22278 5350 22330
rect 5350 22278 5362 22330
rect 5362 22278 5392 22330
rect 5416 22278 5426 22330
rect 5426 22278 5472 22330
rect 5176 22276 5232 22278
rect 5256 22276 5312 22278
rect 5336 22276 5392 22278
rect 5416 22276 5472 22278
rect 5176 21242 5232 21244
rect 5256 21242 5312 21244
rect 5336 21242 5392 21244
rect 5416 21242 5472 21244
rect 5176 21190 5222 21242
rect 5222 21190 5232 21242
rect 5256 21190 5286 21242
rect 5286 21190 5298 21242
rect 5298 21190 5312 21242
rect 5336 21190 5350 21242
rect 5350 21190 5362 21242
rect 5362 21190 5392 21242
rect 5416 21190 5426 21242
rect 5426 21190 5472 21242
rect 5176 21188 5232 21190
rect 5256 21188 5312 21190
rect 5336 21188 5392 21190
rect 5416 21188 5472 21190
rect 5176 20154 5232 20156
rect 5256 20154 5312 20156
rect 5336 20154 5392 20156
rect 5416 20154 5472 20156
rect 5176 20102 5222 20154
rect 5222 20102 5232 20154
rect 5256 20102 5286 20154
rect 5286 20102 5298 20154
rect 5298 20102 5312 20154
rect 5336 20102 5350 20154
rect 5350 20102 5362 20154
rect 5362 20102 5392 20154
rect 5416 20102 5426 20154
rect 5426 20102 5472 20154
rect 5176 20100 5232 20102
rect 5256 20100 5312 20102
rect 5336 20100 5392 20102
rect 5416 20100 5472 20102
rect 9396 37018 9452 37020
rect 9476 37018 9532 37020
rect 9556 37018 9612 37020
rect 9636 37018 9692 37020
rect 9396 36966 9442 37018
rect 9442 36966 9452 37018
rect 9476 36966 9506 37018
rect 9506 36966 9518 37018
rect 9518 36966 9532 37018
rect 9556 36966 9570 37018
rect 9570 36966 9582 37018
rect 9582 36966 9612 37018
rect 9636 36966 9646 37018
rect 9646 36966 9692 37018
rect 9396 36964 9452 36966
rect 9476 36964 9532 36966
rect 9556 36964 9612 36966
rect 9636 36964 9692 36966
rect 9396 35930 9452 35932
rect 9476 35930 9532 35932
rect 9556 35930 9612 35932
rect 9636 35930 9692 35932
rect 9396 35878 9442 35930
rect 9442 35878 9452 35930
rect 9476 35878 9506 35930
rect 9506 35878 9518 35930
rect 9518 35878 9532 35930
rect 9556 35878 9570 35930
rect 9570 35878 9582 35930
rect 9582 35878 9612 35930
rect 9636 35878 9646 35930
rect 9646 35878 9692 35930
rect 9396 35876 9452 35878
rect 9476 35876 9532 35878
rect 9556 35876 9612 35878
rect 9636 35876 9692 35878
rect 9396 34842 9452 34844
rect 9476 34842 9532 34844
rect 9556 34842 9612 34844
rect 9636 34842 9692 34844
rect 9396 34790 9442 34842
rect 9442 34790 9452 34842
rect 9476 34790 9506 34842
rect 9506 34790 9518 34842
rect 9518 34790 9532 34842
rect 9556 34790 9570 34842
rect 9570 34790 9582 34842
rect 9582 34790 9612 34842
rect 9636 34790 9646 34842
rect 9646 34790 9692 34842
rect 9396 34788 9452 34790
rect 9476 34788 9532 34790
rect 9556 34788 9612 34790
rect 9636 34788 9692 34790
rect 9396 33754 9452 33756
rect 9476 33754 9532 33756
rect 9556 33754 9612 33756
rect 9636 33754 9692 33756
rect 9396 33702 9442 33754
rect 9442 33702 9452 33754
rect 9476 33702 9506 33754
rect 9506 33702 9518 33754
rect 9518 33702 9532 33754
rect 9556 33702 9570 33754
rect 9570 33702 9582 33754
rect 9582 33702 9612 33754
rect 9636 33702 9646 33754
rect 9646 33702 9692 33754
rect 9396 33700 9452 33702
rect 9476 33700 9532 33702
rect 9556 33700 9612 33702
rect 9636 33700 9692 33702
rect 11518 35028 11520 35048
rect 11520 35028 11572 35048
rect 11572 35028 11574 35048
rect 11518 34992 11574 35028
rect 9396 32666 9452 32668
rect 9476 32666 9532 32668
rect 9556 32666 9612 32668
rect 9636 32666 9692 32668
rect 9396 32614 9442 32666
rect 9442 32614 9452 32666
rect 9476 32614 9506 32666
rect 9506 32614 9518 32666
rect 9518 32614 9532 32666
rect 9556 32614 9570 32666
rect 9570 32614 9582 32666
rect 9582 32614 9612 32666
rect 9636 32614 9646 32666
rect 9646 32614 9692 32666
rect 9396 32612 9452 32614
rect 9476 32612 9532 32614
rect 9556 32612 9612 32614
rect 9636 32612 9692 32614
rect 9954 32428 10010 32464
rect 10230 32564 10286 32600
rect 10230 32544 10232 32564
rect 10232 32544 10284 32564
rect 10284 32544 10286 32564
rect 9954 32408 9956 32428
rect 9956 32408 10008 32428
rect 10008 32408 10010 32428
rect 9396 31578 9452 31580
rect 9476 31578 9532 31580
rect 9556 31578 9612 31580
rect 9636 31578 9692 31580
rect 9396 31526 9442 31578
rect 9442 31526 9452 31578
rect 9476 31526 9506 31578
rect 9506 31526 9518 31578
rect 9518 31526 9532 31578
rect 9556 31526 9570 31578
rect 9570 31526 9582 31578
rect 9582 31526 9612 31578
rect 9636 31526 9646 31578
rect 9646 31526 9692 31578
rect 9396 31524 9452 31526
rect 9476 31524 9532 31526
rect 9556 31524 9612 31526
rect 9636 31524 9692 31526
rect 9396 30490 9452 30492
rect 9476 30490 9532 30492
rect 9556 30490 9612 30492
rect 9636 30490 9692 30492
rect 9396 30438 9442 30490
rect 9442 30438 9452 30490
rect 9476 30438 9506 30490
rect 9506 30438 9518 30490
rect 9518 30438 9532 30490
rect 9556 30438 9570 30490
rect 9570 30438 9582 30490
rect 9582 30438 9612 30490
rect 9636 30438 9646 30490
rect 9646 30438 9692 30490
rect 9396 30436 9452 30438
rect 9476 30436 9532 30438
rect 9556 30436 9612 30438
rect 9636 30436 9692 30438
rect 10506 32544 10562 32600
rect 10690 32444 10692 32464
rect 10692 32444 10744 32464
rect 10744 32444 10746 32464
rect 10690 32408 10746 32444
rect 13617 37562 13673 37564
rect 13697 37562 13753 37564
rect 13777 37562 13833 37564
rect 13857 37562 13913 37564
rect 13617 37510 13663 37562
rect 13663 37510 13673 37562
rect 13697 37510 13727 37562
rect 13727 37510 13739 37562
rect 13739 37510 13753 37562
rect 13777 37510 13791 37562
rect 13791 37510 13803 37562
rect 13803 37510 13833 37562
rect 13857 37510 13867 37562
rect 13867 37510 13913 37562
rect 13617 37508 13673 37510
rect 13697 37508 13753 37510
rect 13777 37508 13833 37510
rect 13857 37508 13913 37510
rect 11886 34584 11942 34640
rect 9396 29402 9452 29404
rect 9476 29402 9532 29404
rect 9556 29402 9612 29404
rect 9636 29402 9692 29404
rect 9396 29350 9442 29402
rect 9442 29350 9452 29402
rect 9476 29350 9506 29402
rect 9506 29350 9518 29402
rect 9518 29350 9532 29402
rect 9556 29350 9570 29402
rect 9570 29350 9582 29402
rect 9582 29350 9612 29402
rect 9636 29350 9646 29402
rect 9646 29350 9692 29402
rect 9396 29348 9452 29350
rect 9476 29348 9532 29350
rect 9556 29348 9612 29350
rect 9636 29348 9692 29350
rect 9396 28314 9452 28316
rect 9476 28314 9532 28316
rect 9556 28314 9612 28316
rect 9636 28314 9692 28316
rect 9396 28262 9442 28314
rect 9442 28262 9452 28314
rect 9476 28262 9506 28314
rect 9506 28262 9518 28314
rect 9518 28262 9532 28314
rect 9556 28262 9570 28314
rect 9570 28262 9582 28314
rect 9582 28262 9612 28314
rect 9636 28262 9646 28314
rect 9646 28262 9692 28314
rect 9396 28260 9452 28262
rect 9476 28260 9532 28262
rect 9556 28260 9612 28262
rect 9636 28260 9692 28262
rect 9396 27226 9452 27228
rect 9476 27226 9532 27228
rect 9556 27226 9612 27228
rect 9636 27226 9692 27228
rect 9396 27174 9442 27226
rect 9442 27174 9452 27226
rect 9476 27174 9506 27226
rect 9506 27174 9518 27226
rect 9518 27174 9532 27226
rect 9556 27174 9570 27226
rect 9570 27174 9582 27226
rect 9582 27174 9612 27226
rect 9636 27174 9646 27226
rect 9646 27174 9692 27226
rect 9396 27172 9452 27174
rect 9476 27172 9532 27174
rect 9556 27172 9612 27174
rect 9636 27172 9692 27174
rect 9396 26138 9452 26140
rect 9476 26138 9532 26140
rect 9556 26138 9612 26140
rect 9636 26138 9692 26140
rect 9396 26086 9442 26138
rect 9442 26086 9452 26138
rect 9476 26086 9506 26138
rect 9506 26086 9518 26138
rect 9518 26086 9532 26138
rect 9556 26086 9570 26138
rect 9570 26086 9582 26138
rect 9582 26086 9612 26138
rect 9636 26086 9646 26138
rect 9646 26086 9692 26138
rect 9396 26084 9452 26086
rect 9476 26084 9532 26086
rect 9556 26084 9612 26086
rect 9636 26084 9692 26086
rect 13617 36474 13673 36476
rect 13697 36474 13753 36476
rect 13777 36474 13833 36476
rect 13857 36474 13913 36476
rect 13617 36422 13663 36474
rect 13663 36422 13673 36474
rect 13697 36422 13727 36474
rect 13727 36422 13739 36474
rect 13739 36422 13753 36474
rect 13777 36422 13791 36474
rect 13791 36422 13803 36474
rect 13803 36422 13833 36474
rect 13857 36422 13867 36474
rect 13867 36422 13913 36474
rect 13617 36420 13673 36422
rect 13697 36420 13753 36422
rect 13777 36420 13833 36422
rect 13857 36420 13913 36422
rect 13617 35386 13673 35388
rect 13697 35386 13753 35388
rect 13777 35386 13833 35388
rect 13857 35386 13913 35388
rect 13617 35334 13663 35386
rect 13663 35334 13673 35386
rect 13697 35334 13727 35386
rect 13727 35334 13739 35386
rect 13739 35334 13753 35386
rect 13777 35334 13791 35386
rect 13791 35334 13803 35386
rect 13803 35334 13833 35386
rect 13857 35334 13867 35386
rect 13867 35334 13913 35386
rect 13617 35332 13673 35334
rect 13697 35332 13753 35334
rect 13777 35332 13833 35334
rect 13857 35332 13913 35334
rect 13617 34298 13673 34300
rect 13697 34298 13753 34300
rect 13777 34298 13833 34300
rect 13857 34298 13913 34300
rect 13617 34246 13663 34298
rect 13663 34246 13673 34298
rect 13697 34246 13727 34298
rect 13727 34246 13739 34298
rect 13739 34246 13753 34298
rect 13777 34246 13791 34298
rect 13791 34246 13803 34298
rect 13803 34246 13833 34298
rect 13857 34246 13867 34298
rect 13867 34246 13913 34298
rect 13617 34244 13673 34246
rect 13697 34244 13753 34246
rect 13777 34244 13833 34246
rect 13857 34244 13913 34246
rect 15198 34584 15254 34640
rect 13617 33210 13673 33212
rect 13697 33210 13753 33212
rect 13777 33210 13833 33212
rect 13857 33210 13913 33212
rect 13617 33158 13663 33210
rect 13663 33158 13673 33210
rect 13697 33158 13727 33210
rect 13727 33158 13739 33210
rect 13739 33158 13753 33210
rect 13777 33158 13791 33210
rect 13791 33158 13803 33210
rect 13803 33158 13833 33210
rect 13857 33158 13867 33210
rect 13867 33158 13913 33210
rect 13617 33156 13673 33158
rect 13697 33156 13753 33158
rect 13777 33156 13833 33158
rect 13857 33156 13913 33158
rect 14002 32272 14058 32328
rect 13617 32122 13673 32124
rect 13697 32122 13753 32124
rect 13777 32122 13833 32124
rect 13857 32122 13913 32124
rect 13617 32070 13663 32122
rect 13663 32070 13673 32122
rect 13697 32070 13727 32122
rect 13727 32070 13739 32122
rect 13739 32070 13753 32122
rect 13777 32070 13791 32122
rect 13791 32070 13803 32122
rect 13803 32070 13833 32122
rect 13857 32070 13867 32122
rect 13867 32070 13913 32122
rect 13617 32068 13673 32070
rect 13697 32068 13753 32070
rect 13777 32068 13833 32070
rect 13857 32068 13913 32070
rect 14830 32952 14886 33008
rect 14738 32408 14794 32464
rect 13617 31034 13673 31036
rect 13697 31034 13753 31036
rect 13777 31034 13833 31036
rect 13857 31034 13913 31036
rect 13617 30982 13663 31034
rect 13663 30982 13673 31034
rect 13697 30982 13727 31034
rect 13727 30982 13739 31034
rect 13739 30982 13753 31034
rect 13777 30982 13791 31034
rect 13791 30982 13803 31034
rect 13803 30982 13833 31034
rect 13857 30982 13867 31034
rect 13867 30982 13913 31034
rect 13617 30980 13673 30982
rect 13697 30980 13753 30982
rect 13777 30980 13833 30982
rect 13857 30980 13913 30982
rect 13617 29946 13673 29948
rect 13697 29946 13753 29948
rect 13777 29946 13833 29948
rect 13857 29946 13913 29948
rect 13617 29894 13663 29946
rect 13663 29894 13673 29946
rect 13697 29894 13727 29946
rect 13727 29894 13739 29946
rect 13739 29894 13753 29946
rect 13777 29894 13791 29946
rect 13791 29894 13803 29946
rect 13803 29894 13833 29946
rect 13857 29894 13867 29946
rect 13867 29894 13913 29946
rect 13617 29892 13673 29894
rect 13697 29892 13753 29894
rect 13777 29892 13833 29894
rect 13857 29892 13913 29894
rect 13617 28858 13673 28860
rect 13697 28858 13753 28860
rect 13777 28858 13833 28860
rect 13857 28858 13913 28860
rect 13617 28806 13663 28858
rect 13663 28806 13673 28858
rect 13697 28806 13727 28858
rect 13727 28806 13739 28858
rect 13739 28806 13753 28858
rect 13777 28806 13791 28858
rect 13791 28806 13803 28858
rect 13803 28806 13833 28858
rect 13857 28806 13867 28858
rect 13867 28806 13913 28858
rect 13617 28804 13673 28806
rect 13697 28804 13753 28806
rect 13777 28804 13833 28806
rect 13857 28804 13913 28806
rect 9396 25050 9452 25052
rect 9476 25050 9532 25052
rect 9556 25050 9612 25052
rect 9636 25050 9692 25052
rect 9396 24998 9442 25050
rect 9442 24998 9452 25050
rect 9476 24998 9506 25050
rect 9506 24998 9518 25050
rect 9518 24998 9532 25050
rect 9556 24998 9570 25050
rect 9570 24998 9582 25050
rect 9582 24998 9612 25050
rect 9636 24998 9646 25050
rect 9646 24998 9692 25050
rect 9396 24996 9452 24998
rect 9476 24996 9532 24998
rect 9556 24996 9612 24998
rect 9636 24996 9692 24998
rect 9396 23962 9452 23964
rect 9476 23962 9532 23964
rect 9556 23962 9612 23964
rect 9636 23962 9692 23964
rect 9396 23910 9442 23962
rect 9442 23910 9452 23962
rect 9476 23910 9506 23962
rect 9506 23910 9518 23962
rect 9518 23910 9532 23962
rect 9556 23910 9570 23962
rect 9570 23910 9582 23962
rect 9582 23910 9612 23962
rect 9636 23910 9646 23962
rect 9646 23910 9692 23962
rect 9396 23908 9452 23910
rect 9476 23908 9532 23910
rect 9556 23908 9612 23910
rect 9636 23908 9692 23910
rect 9396 22874 9452 22876
rect 9476 22874 9532 22876
rect 9556 22874 9612 22876
rect 9636 22874 9692 22876
rect 9396 22822 9442 22874
rect 9442 22822 9452 22874
rect 9476 22822 9506 22874
rect 9506 22822 9518 22874
rect 9518 22822 9532 22874
rect 9556 22822 9570 22874
rect 9570 22822 9582 22874
rect 9582 22822 9612 22874
rect 9636 22822 9646 22874
rect 9646 22822 9692 22874
rect 9396 22820 9452 22822
rect 9476 22820 9532 22822
rect 9556 22820 9612 22822
rect 9636 22820 9692 22822
rect 9396 21786 9452 21788
rect 9476 21786 9532 21788
rect 9556 21786 9612 21788
rect 9636 21786 9692 21788
rect 9396 21734 9442 21786
rect 9442 21734 9452 21786
rect 9476 21734 9506 21786
rect 9506 21734 9518 21786
rect 9518 21734 9532 21786
rect 9556 21734 9570 21786
rect 9570 21734 9582 21786
rect 9582 21734 9612 21786
rect 9636 21734 9646 21786
rect 9646 21734 9692 21786
rect 9396 21732 9452 21734
rect 9476 21732 9532 21734
rect 9556 21732 9612 21734
rect 9636 21732 9692 21734
rect 9396 20698 9452 20700
rect 9476 20698 9532 20700
rect 9556 20698 9612 20700
rect 9636 20698 9692 20700
rect 9396 20646 9442 20698
rect 9442 20646 9452 20698
rect 9476 20646 9506 20698
rect 9506 20646 9518 20698
rect 9518 20646 9532 20698
rect 9556 20646 9570 20698
rect 9570 20646 9582 20698
rect 9582 20646 9612 20698
rect 9636 20646 9646 20698
rect 9646 20646 9692 20698
rect 9396 20644 9452 20646
rect 9476 20644 9532 20646
rect 9556 20644 9612 20646
rect 9636 20644 9692 20646
rect 9396 19610 9452 19612
rect 9476 19610 9532 19612
rect 9556 19610 9612 19612
rect 9636 19610 9692 19612
rect 9396 19558 9442 19610
rect 9442 19558 9452 19610
rect 9476 19558 9506 19610
rect 9506 19558 9518 19610
rect 9518 19558 9532 19610
rect 9556 19558 9570 19610
rect 9570 19558 9582 19610
rect 9582 19558 9612 19610
rect 9636 19558 9646 19610
rect 9646 19558 9692 19610
rect 9396 19556 9452 19558
rect 9476 19556 9532 19558
rect 9556 19556 9612 19558
rect 9636 19556 9692 19558
rect 13617 27770 13673 27772
rect 13697 27770 13753 27772
rect 13777 27770 13833 27772
rect 13857 27770 13913 27772
rect 13617 27718 13663 27770
rect 13663 27718 13673 27770
rect 13697 27718 13727 27770
rect 13727 27718 13739 27770
rect 13739 27718 13753 27770
rect 13777 27718 13791 27770
rect 13791 27718 13803 27770
rect 13803 27718 13833 27770
rect 13857 27718 13867 27770
rect 13867 27718 13913 27770
rect 13617 27716 13673 27718
rect 13697 27716 13753 27718
rect 13777 27716 13833 27718
rect 13857 27716 13913 27718
rect 13617 26682 13673 26684
rect 13697 26682 13753 26684
rect 13777 26682 13833 26684
rect 13857 26682 13913 26684
rect 13617 26630 13663 26682
rect 13663 26630 13673 26682
rect 13697 26630 13727 26682
rect 13727 26630 13739 26682
rect 13739 26630 13753 26682
rect 13777 26630 13791 26682
rect 13791 26630 13803 26682
rect 13803 26630 13833 26682
rect 13857 26630 13867 26682
rect 13867 26630 13913 26682
rect 13617 26628 13673 26630
rect 13697 26628 13753 26630
rect 13777 26628 13833 26630
rect 13857 26628 13913 26630
rect 15474 36080 15530 36136
rect 15658 34604 15714 34640
rect 17837 39194 17893 39196
rect 17917 39194 17973 39196
rect 17997 39194 18053 39196
rect 18077 39194 18133 39196
rect 17837 39142 17883 39194
rect 17883 39142 17893 39194
rect 17917 39142 17947 39194
rect 17947 39142 17959 39194
rect 17959 39142 17973 39194
rect 17997 39142 18011 39194
rect 18011 39142 18023 39194
rect 18023 39142 18053 39194
rect 18077 39142 18087 39194
rect 18087 39142 18133 39194
rect 17837 39140 17893 39142
rect 17917 39140 17973 39142
rect 17997 39140 18053 39142
rect 18077 39140 18133 39142
rect 17837 38106 17893 38108
rect 17917 38106 17973 38108
rect 17997 38106 18053 38108
rect 18077 38106 18133 38108
rect 17837 38054 17883 38106
rect 17883 38054 17893 38106
rect 17917 38054 17947 38106
rect 17947 38054 17959 38106
rect 17959 38054 17973 38106
rect 17997 38054 18011 38106
rect 18011 38054 18023 38106
rect 18023 38054 18053 38106
rect 18077 38054 18087 38106
rect 18087 38054 18133 38106
rect 17837 38052 17893 38054
rect 17917 38052 17973 38054
rect 17997 38052 18053 38054
rect 18077 38052 18133 38054
rect 22058 39738 22114 39740
rect 22138 39738 22194 39740
rect 22218 39738 22274 39740
rect 22298 39738 22354 39740
rect 22058 39686 22104 39738
rect 22104 39686 22114 39738
rect 22138 39686 22168 39738
rect 22168 39686 22180 39738
rect 22180 39686 22194 39738
rect 22218 39686 22232 39738
rect 22232 39686 22244 39738
rect 22244 39686 22274 39738
rect 22298 39686 22308 39738
rect 22308 39686 22354 39738
rect 22058 39684 22114 39686
rect 22138 39684 22194 39686
rect 22218 39684 22274 39686
rect 22298 39684 22354 39686
rect 17837 37018 17893 37020
rect 17917 37018 17973 37020
rect 17997 37018 18053 37020
rect 18077 37018 18133 37020
rect 17837 36966 17883 37018
rect 17883 36966 17893 37018
rect 17917 36966 17947 37018
rect 17947 36966 17959 37018
rect 17959 36966 17973 37018
rect 17997 36966 18011 37018
rect 18011 36966 18023 37018
rect 18023 36966 18053 37018
rect 18077 36966 18087 37018
rect 18087 36966 18133 37018
rect 17837 36964 17893 36966
rect 17917 36964 17973 36966
rect 17997 36964 18053 36966
rect 18077 36964 18133 36966
rect 15658 34584 15660 34604
rect 15660 34584 15712 34604
rect 15712 34584 15714 34604
rect 16486 34584 16542 34640
rect 15290 32308 15292 32328
rect 15292 32308 15344 32328
rect 15344 32308 15346 32328
rect 15290 32272 15346 32308
rect 13617 25594 13673 25596
rect 13697 25594 13753 25596
rect 13777 25594 13833 25596
rect 13857 25594 13913 25596
rect 13617 25542 13663 25594
rect 13663 25542 13673 25594
rect 13697 25542 13727 25594
rect 13727 25542 13739 25594
rect 13739 25542 13753 25594
rect 13777 25542 13791 25594
rect 13791 25542 13803 25594
rect 13803 25542 13833 25594
rect 13857 25542 13867 25594
rect 13867 25542 13913 25594
rect 13617 25540 13673 25542
rect 13697 25540 13753 25542
rect 13777 25540 13833 25542
rect 13857 25540 13913 25542
rect 13617 24506 13673 24508
rect 13697 24506 13753 24508
rect 13777 24506 13833 24508
rect 13857 24506 13913 24508
rect 13617 24454 13663 24506
rect 13663 24454 13673 24506
rect 13697 24454 13727 24506
rect 13727 24454 13739 24506
rect 13739 24454 13753 24506
rect 13777 24454 13791 24506
rect 13791 24454 13803 24506
rect 13803 24454 13833 24506
rect 13857 24454 13867 24506
rect 13867 24454 13913 24506
rect 13617 24452 13673 24454
rect 13697 24452 13753 24454
rect 13777 24452 13833 24454
rect 13857 24452 13913 24454
rect 13726 23724 13782 23760
rect 13726 23704 13728 23724
rect 13728 23704 13780 23724
rect 13780 23704 13782 23724
rect 13617 23418 13673 23420
rect 13697 23418 13753 23420
rect 13777 23418 13833 23420
rect 13857 23418 13913 23420
rect 13617 23366 13663 23418
rect 13663 23366 13673 23418
rect 13697 23366 13727 23418
rect 13727 23366 13739 23418
rect 13739 23366 13753 23418
rect 13777 23366 13791 23418
rect 13791 23366 13803 23418
rect 13803 23366 13833 23418
rect 13857 23366 13867 23418
rect 13867 23366 13913 23418
rect 13617 23364 13673 23366
rect 13697 23364 13753 23366
rect 13777 23364 13833 23366
rect 13857 23364 13913 23366
rect 16578 32816 16634 32872
rect 22058 38650 22114 38652
rect 22138 38650 22194 38652
rect 22218 38650 22274 38652
rect 22298 38650 22354 38652
rect 22058 38598 22104 38650
rect 22104 38598 22114 38650
rect 22138 38598 22168 38650
rect 22168 38598 22180 38650
rect 22180 38598 22194 38650
rect 22218 38598 22232 38650
rect 22232 38598 22244 38650
rect 22244 38598 22274 38650
rect 22298 38598 22308 38650
rect 22308 38598 22354 38650
rect 22058 38596 22114 38598
rect 22138 38596 22194 38598
rect 22218 38596 22274 38598
rect 22298 38596 22354 38598
rect 22058 37562 22114 37564
rect 22138 37562 22194 37564
rect 22218 37562 22274 37564
rect 22298 37562 22354 37564
rect 22058 37510 22104 37562
rect 22104 37510 22114 37562
rect 22138 37510 22168 37562
rect 22168 37510 22180 37562
rect 22180 37510 22194 37562
rect 22218 37510 22232 37562
rect 22232 37510 22244 37562
rect 22244 37510 22274 37562
rect 22298 37510 22308 37562
rect 22308 37510 22354 37562
rect 22058 37508 22114 37510
rect 22138 37508 22194 37510
rect 22218 37508 22274 37510
rect 22298 37508 22354 37510
rect 18510 36080 18566 36136
rect 17837 35930 17893 35932
rect 17917 35930 17973 35932
rect 17997 35930 18053 35932
rect 18077 35930 18133 35932
rect 17837 35878 17883 35930
rect 17883 35878 17893 35930
rect 17917 35878 17947 35930
rect 17947 35878 17959 35930
rect 17959 35878 17973 35930
rect 17997 35878 18011 35930
rect 18011 35878 18023 35930
rect 18023 35878 18053 35930
rect 18077 35878 18087 35930
rect 18087 35878 18133 35930
rect 17837 35876 17893 35878
rect 17917 35876 17973 35878
rect 17997 35876 18053 35878
rect 18077 35876 18133 35878
rect 17837 34842 17893 34844
rect 17917 34842 17973 34844
rect 17997 34842 18053 34844
rect 18077 34842 18133 34844
rect 17837 34790 17883 34842
rect 17883 34790 17893 34842
rect 17917 34790 17947 34842
rect 17947 34790 17959 34842
rect 17959 34790 17973 34842
rect 17997 34790 18011 34842
rect 18011 34790 18023 34842
rect 18023 34790 18053 34842
rect 18077 34790 18087 34842
rect 18087 34790 18133 34842
rect 17837 34788 17893 34790
rect 17917 34788 17973 34790
rect 17997 34788 18053 34790
rect 18077 34788 18133 34790
rect 18786 34584 18842 34640
rect 17837 33754 17893 33756
rect 17917 33754 17973 33756
rect 17997 33754 18053 33756
rect 18077 33754 18133 33756
rect 17837 33702 17883 33754
rect 17883 33702 17893 33754
rect 17917 33702 17947 33754
rect 17947 33702 17959 33754
rect 17959 33702 17973 33754
rect 17997 33702 18011 33754
rect 18011 33702 18023 33754
rect 18023 33702 18053 33754
rect 18077 33702 18087 33754
rect 18087 33702 18133 33754
rect 17837 33700 17893 33702
rect 17917 33700 17973 33702
rect 17997 33700 18053 33702
rect 18077 33700 18133 33702
rect 17590 32408 17646 32464
rect 15934 29552 15990 29608
rect 17866 32816 17922 32872
rect 18142 32852 18144 32872
rect 18144 32852 18196 32872
rect 18196 32852 18198 32872
rect 18142 32816 18198 32852
rect 17837 32666 17893 32668
rect 17917 32666 17973 32668
rect 17997 32666 18053 32668
rect 18077 32666 18133 32668
rect 17837 32614 17883 32666
rect 17883 32614 17893 32666
rect 17917 32614 17947 32666
rect 17947 32614 17959 32666
rect 17959 32614 17973 32666
rect 17997 32614 18011 32666
rect 18011 32614 18023 32666
rect 18023 32614 18053 32666
rect 18077 32614 18087 32666
rect 18087 32614 18133 32666
rect 17837 32612 17893 32614
rect 17917 32612 17973 32614
rect 17997 32612 18053 32614
rect 18077 32612 18133 32614
rect 18234 32308 18236 32328
rect 18236 32308 18288 32328
rect 18288 32308 18290 32328
rect 18234 32272 18290 32308
rect 17837 31578 17893 31580
rect 17917 31578 17973 31580
rect 17997 31578 18053 31580
rect 18077 31578 18133 31580
rect 17837 31526 17883 31578
rect 17883 31526 17893 31578
rect 17917 31526 17947 31578
rect 17947 31526 17959 31578
rect 17959 31526 17973 31578
rect 17997 31526 18011 31578
rect 18011 31526 18023 31578
rect 18023 31526 18053 31578
rect 18077 31526 18087 31578
rect 18087 31526 18133 31578
rect 17837 31524 17893 31526
rect 17917 31524 17973 31526
rect 17997 31524 18053 31526
rect 18077 31524 18133 31526
rect 17837 30490 17893 30492
rect 17917 30490 17973 30492
rect 17997 30490 18053 30492
rect 18077 30490 18133 30492
rect 17837 30438 17883 30490
rect 17883 30438 17893 30490
rect 17917 30438 17947 30490
rect 17947 30438 17959 30490
rect 17959 30438 17973 30490
rect 17997 30438 18011 30490
rect 18011 30438 18023 30490
rect 18023 30438 18053 30490
rect 18077 30438 18087 30490
rect 18087 30438 18133 30490
rect 17837 30436 17893 30438
rect 17917 30436 17973 30438
rect 17997 30436 18053 30438
rect 18077 30436 18133 30438
rect 18142 29572 18198 29608
rect 18142 29552 18144 29572
rect 18144 29552 18196 29572
rect 18196 29552 18198 29572
rect 17837 29402 17893 29404
rect 17917 29402 17973 29404
rect 17997 29402 18053 29404
rect 18077 29402 18133 29404
rect 17837 29350 17883 29402
rect 17883 29350 17893 29402
rect 17917 29350 17947 29402
rect 17947 29350 17959 29402
rect 17959 29350 17973 29402
rect 17997 29350 18011 29402
rect 18011 29350 18023 29402
rect 18023 29350 18053 29402
rect 18077 29350 18087 29402
rect 18087 29350 18133 29402
rect 17837 29348 17893 29350
rect 17917 29348 17973 29350
rect 17997 29348 18053 29350
rect 18077 29348 18133 29350
rect 17498 29144 17554 29200
rect 18326 30368 18382 30424
rect 19154 34992 19210 35048
rect 19154 32408 19210 32464
rect 13617 22330 13673 22332
rect 13697 22330 13753 22332
rect 13777 22330 13833 22332
rect 13857 22330 13913 22332
rect 13617 22278 13663 22330
rect 13663 22278 13673 22330
rect 13697 22278 13727 22330
rect 13727 22278 13739 22330
rect 13739 22278 13753 22330
rect 13777 22278 13791 22330
rect 13791 22278 13803 22330
rect 13803 22278 13833 22330
rect 13857 22278 13867 22330
rect 13867 22278 13913 22330
rect 13617 22276 13673 22278
rect 13697 22276 13753 22278
rect 13777 22276 13833 22278
rect 13857 22276 13913 22278
rect 13617 21242 13673 21244
rect 13697 21242 13753 21244
rect 13777 21242 13833 21244
rect 13857 21242 13913 21244
rect 13617 21190 13663 21242
rect 13663 21190 13673 21242
rect 13697 21190 13727 21242
rect 13727 21190 13739 21242
rect 13739 21190 13753 21242
rect 13777 21190 13791 21242
rect 13791 21190 13803 21242
rect 13803 21190 13833 21242
rect 13857 21190 13867 21242
rect 13867 21190 13913 21242
rect 13617 21188 13673 21190
rect 13697 21188 13753 21190
rect 13777 21188 13833 21190
rect 13857 21188 13913 21190
rect 13617 20154 13673 20156
rect 13697 20154 13753 20156
rect 13777 20154 13833 20156
rect 13857 20154 13913 20156
rect 13617 20102 13663 20154
rect 13663 20102 13673 20154
rect 13697 20102 13727 20154
rect 13727 20102 13739 20154
rect 13739 20102 13753 20154
rect 13777 20102 13791 20154
rect 13791 20102 13803 20154
rect 13803 20102 13833 20154
rect 13857 20102 13867 20154
rect 13867 20102 13913 20154
rect 13617 20100 13673 20102
rect 13697 20100 13753 20102
rect 13777 20100 13833 20102
rect 13857 20100 13913 20102
rect 15566 23724 15622 23760
rect 15566 23704 15568 23724
rect 15568 23704 15620 23724
rect 15620 23704 15622 23724
rect 17837 28314 17893 28316
rect 17917 28314 17973 28316
rect 17997 28314 18053 28316
rect 18077 28314 18133 28316
rect 17837 28262 17883 28314
rect 17883 28262 17893 28314
rect 17917 28262 17947 28314
rect 17947 28262 17959 28314
rect 17959 28262 17973 28314
rect 17997 28262 18011 28314
rect 18011 28262 18023 28314
rect 18023 28262 18053 28314
rect 18077 28262 18087 28314
rect 18087 28262 18133 28314
rect 17837 28260 17893 28262
rect 17917 28260 17973 28262
rect 17997 28260 18053 28262
rect 18077 28260 18133 28262
rect 17837 27226 17893 27228
rect 17917 27226 17973 27228
rect 17997 27226 18053 27228
rect 18077 27226 18133 27228
rect 17837 27174 17883 27226
rect 17883 27174 17893 27226
rect 17917 27174 17947 27226
rect 17947 27174 17959 27226
rect 17959 27174 17973 27226
rect 17997 27174 18011 27226
rect 18011 27174 18023 27226
rect 18023 27174 18053 27226
rect 18077 27174 18087 27226
rect 18087 27174 18133 27226
rect 17837 27172 17893 27174
rect 17917 27172 17973 27174
rect 17997 27172 18053 27174
rect 18077 27172 18133 27174
rect 17837 26138 17893 26140
rect 17917 26138 17973 26140
rect 17997 26138 18053 26140
rect 18077 26138 18133 26140
rect 17837 26086 17883 26138
rect 17883 26086 17893 26138
rect 17917 26086 17947 26138
rect 17947 26086 17959 26138
rect 17959 26086 17973 26138
rect 17997 26086 18011 26138
rect 18011 26086 18023 26138
rect 18023 26086 18053 26138
rect 18077 26086 18087 26138
rect 18087 26086 18133 26138
rect 17837 26084 17893 26086
rect 17917 26084 17973 26086
rect 17997 26084 18053 26086
rect 18077 26084 18133 26086
rect 19522 32852 19524 32872
rect 19524 32852 19576 32872
rect 19576 32852 19578 32872
rect 19522 32816 19578 32852
rect 19430 32272 19486 32328
rect 22058 36474 22114 36476
rect 22138 36474 22194 36476
rect 22218 36474 22274 36476
rect 22298 36474 22354 36476
rect 22058 36422 22104 36474
rect 22104 36422 22114 36474
rect 22138 36422 22168 36474
rect 22168 36422 22180 36474
rect 22180 36422 22194 36474
rect 22218 36422 22232 36474
rect 22232 36422 22244 36474
rect 22244 36422 22274 36474
rect 22298 36422 22308 36474
rect 22308 36422 22354 36474
rect 22058 36420 22114 36422
rect 22138 36420 22194 36422
rect 22218 36420 22274 36422
rect 22298 36420 22354 36422
rect 22058 35386 22114 35388
rect 22138 35386 22194 35388
rect 22218 35386 22274 35388
rect 22298 35386 22354 35388
rect 22058 35334 22104 35386
rect 22104 35334 22114 35386
rect 22138 35334 22168 35386
rect 22168 35334 22180 35386
rect 22180 35334 22194 35386
rect 22218 35334 22232 35386
rect 22232 35334 22244 35386
rect 22244 35334 22274 35386
rect 22298 35334 22308 35386
rect 22308 35334 22354 35386
rect 22058 35332 22114 35334
rect 22138 35332 22194 35334
rect 22218 35332 22274 35334
rect 22298 35332 22354 35334
rect 22058 34298 22114 34300
rect 22138 34298 22194 34300
rect 22218 34298 22274 34300
rect 22298 34298 22354 34300
rect 22058 34246 22104 34298
rect 22104 34246 22114 34298
rect 22138 34246 22168 34298
rect 22168 34246 22180 34298
rect 22180 34246 22194 34298
rect 22218 34246 22232 34298
rect 22232 34246 22244 34298
rect 22244 34246 22274 34298
rect 22298 34246 22308 34298
rect 22308 34246 22354 34298
rect 22058 34244 22114 34246
rect 22138 34244 22194 34246
rect 22218 34244 22274 34246
rect 22298 34244 22354 34246
rect 19982 30368 20038 30424
rect 20534 30368 20590 30424
rect 17837 25050 17893 25052
rect 17917 25050 17973 25052
rect 17997 25050 18053 25052
rect 18077 25050 18133 25052
rect 17837 24998 17883 25050
rect 17883 24998 17893 25050
rect 17917 24998 17947 25050
rect 17947 24998 17959 25050
rect 17959 24998 17973 25050
rect 17997 24998 18011 25050
rect 18011 24998 18023 25050
rect 18023 24998 18053 25050
rect 18077 24998 18087 25050
rect 18087 24998 18133 25050
rect 17837 24996 17893 24998
rect 17917 24996 17973 24998
rect 17997 24996 18053 24998
rect 18077 24996 18133 24998
rect 17837 23962 17893 23964
rect 17917 23962 17973 23964
rect 17997 23962 18053 23964
rect 18077 23962 18133 23964
rect 17837 23910 17883 23962
rect 17883 23910 17893 23962
rect 17917 23910 17947 23962
rect 17947 23910 17959 23962
rect 17959 23910 17973 23962
rect 17997 23910 18011 23962
rect 18011 23910 18023 23962
rect 18023 23910 18053 23962
rect 18077 23910 18087 23962
rect 18087 23910 18133 23962
rect 17837 23908 17893 23910
rect 17917 23908 17973 23910
rect 17997 23908 18053 23910
rect 18077 23908 18133 23910
rect 19338 29164 19394 29200
rect 19338 29144 19340 29164
rect 19340 29144 19392 29164
rect 19392 29144 19394 29164
rect 22058 33210 22114 33212
rect 22138 33210 22194 33212
rect 22218 33210 22274 33212
rect 22298 33210 22354 33212
rect 22058 33158 22104 33210
rect 22104 33158 22114 33210
rect 22138 33158 22168 33210
rect 22168 33158 22180 33210
rect 22180 33158 22194 33210
rect 22218 33158 22232 33210
rect 22232 33158 22244 33210
rect 22244 33158 22274 33210
rect 22298 33158 22308 33210
rect 22308 33158 22354 33210
rect 22058 33156 22114 33158
rect 22138 33156 22194 33158
rect 22218 33156 22274 33158
rect 22298 33156 22354 33158
rect 22058 32122 22114 32124
rect 22138 32122 22194 32124
rect 22218 32122 22274 32124
rect 22298 32122 22354 32124
rect 22058 32070 22104 32122
rect 22104 32070 22114 32122
rect 22138 32070 22168 32122
rect 22168 32070 22180 32122
rect 22180 32070 22194 32122
rect 22218 32070 22232 32122
rect 22232 32070 22244 32122
rect 22244 32070 22274 32122
rect 22298 32070 22308 32122
rect 22308 32070 22354 32122
rect 22058 32068 22114 32070
rect 22138 32068 22194 32070
rect 22218 32068 22274 32070
rect 22298 32068 22354 32070
rect 22058 31034 22114 31036
rect 22138 31034 22194 31036
rect 22218 31034 22274 31036
rect 22298 31034 22354 31036
rect 22058 30982 22104 31034
rect 22104 30982 22114 31034
rect 22138 30982 22168 31034
rect 22168 30982 22180 31034
rect 22180 30982 22194 31034
rect 22218 30982 22232 31034
rect 22232 30982 22244 31034
rect 22244 30982 22274 31034
rect 22298 30982 22308 31034
rect 22308 30982 22354 31034
rect 22058 30980 22114 30982
rect 22138 30980 22194 30982
rect 22218 30980 22274 30982
rect 22298 30980 22354 30982
rect 19798 27124 19854 27160
rect 19798 27104 19800 27124
rect 19800 27104 19852 27124
rect 19852 27104 19854 27124
rect 17837 22874 17893 22876
rect 17917 22874 17973 22876
rect 17997 22874 18053 22876
rect 18077 22874 18133 22876
rect 17837 22822 17883 22874
rect 17883 22822 17893 22874
rect 17917 22822 17947 22874
rect 17947 22822 17959 22874
rect 17959 22822 17973 22874
rect 17997 22822 18011 22874
rect 18011 22822 18023 22874
rect 18023 22822 18053 22874
rect 18077 22822 18087 22874
rect 18087 22822 18133 22874
rect 17837 22820 17893 22822
rect 17917 22820 17973 22822
rect 17997 22820 18053 22822
rect 18077 22820 18133 22822
rect 17837 21786 17893 21788
rect 17917 21786 17973 21788
rect 17997 21786 18053 21788
rect 18077 21786 18133 21788
rect 17837 21734 17883 21786
rect 17883 21734 17893 21786
rect 17917 21734 17947 21786
rect 17947 21734 17959 21786
rect 17959 21734 17973 21786
rect 17997 21734 18011 21786
rect 18011 21734 18023 21786
rect 18023 21734 18053 21786
rect 18077 21734 18087 21786
rect 18087 21734 18133 21786
rect 17837 21732 17893 21734
rect 17917 21732 17973 21734
rect 17997 21732 18053 21734
rect 18077 21732 18133 21734
rect 17837 20698 17893 20700
rect 17917 20698 17973 20700
rect 17997 20698 18053 20700
rect 18077 20698 18133 20700
rect 17837 20646 17883 20698
rect 17883 20646 17893 20698
rect 17917 20646 17947 20698
rect 17947 20646 17959 20698
rect 17959 20646 17973 20698
rect 17997 20646 18011 20698
rect 18011 20646 18023 20698
rect 18023 20646 18053 20698
rect 18077 20646 18087 20698
rect 18087 20646 18133 20698
rect 17837 20644 17893 20646
rect 17917 20644 17973 20646
rect 17997 20644 18053 20646
rect 18077 20644 18133 20646
rect 17837 19610 17893 19612
rect 17917 19610 17973 19612
rect 17997 19610 18053 19612
rect 18077 19610 18133 19612
rect 17837 19558 17883 19610
rect 17883 19558 17893 19610
rect 17917 19558 17947 19610
rect 17947 19558 17959 19610
rect 17959 19558 17973 19610
rect 17997 19558 18011 19610
rect 18011 19558 18023 19610
rect 18023 19558 18053 19610
rect 18077 19558 18087 19610
rect 18087 19558 18133 19610
rect 17837 19556 17893 19558
rect 17917 19556 17973 19558
rect 17997 19556 18053 19558
rect 18077 19556 18133 19558
rect 26278 39194 26334 39196
rect 26358 39194 26414 39196
rect 26438 39194 26494 39196
rect 26518 39194 26574 39196
rect 26278 39142 26324 39194
rect 26324 39142 26334 39194
rect 26358 39142 26388 39194
rect 26388 39142 26400 39194
rect 26400 39142 26414 39194
rect 26438 39142 26452 39194
rect 26452 39142 26464 39194
rect 26464 39142 26494 39194
rect 26518 39142 26528 39194
rect 26528 39142 26574 39194
rect 26278 39140 26334 39142
rect 26358 39140 26414 39142
rect 26438 39140 26494 39142
rect 26518 39140 26574 39142
rect 26278 38106 26334 38108
rect 26358 38106 26414 38108
rect 26438 38106 26494 38108
rect 26518 38106 26574 38108
rect 26278 38054 26324 38106
rect 26324 38054 26334 38106
rect 26358 38054 26388 38106
rect 26388 38054 26400 38106
rect 26400 38054 26414 38106
rect 26438 38054 26452 38106
rect 26452 38054 26464 38106
rect 26464 38054 26494 38106
rect 26518 38054 26528 38106
rect 26528 38054 26574 38106
rect 26278 38052 26334 38054
rect 26358 38052 26414 38054
rect 26438 38052 26494 38054
rect 26518 38052 26574 38054
rect 26278 37018 26334 37020
rect 26358 37018 26414 37020
rect 26438 37018 26494 37020
rect 26518 37018 26574 37020
rect 26278 36966 26324 37018
rect 26324 36966 26334 37018
rect 26358 36966 26388 37018
rect 26388 36966 26400 37018
rect 26400 36966 26414 37018
rect 26438 36966 26452 37018
rect 26452 36966 26464 37018
rect 26464 36966 26494 37018
rect 26518 36966 26528 37018
rect 26528 36966 26574 37018
rect 26278 36964 26334 36966
rect 26358 36964 26414 36966
rect 26438 36964 26494 36966
rect 26518 36964 26574 36966
rect 26278 35930 26334 35932
rect 26358 35930 26414 35932
rect 26438 35930 26494 35932
rect 26518 35930 26574 35932
rect 26278 35878 26324 35930
rect 26324 35878 26334 35930
rect 26358 35878 26388 35930
rect 26388 35878 26400 35930
rect 26400 35878 26414 35930
rect 26438 35878 26452 35930
rect 26452 35878 26464 35930
rect 26464 35878 26494 35930
rect 26518 35878 26528 35930
rect 26528 35878 26574 35930
rect 26278 35876 26334 35878
rect 26358 35876 26414 35878
rect 26438 35876 26494 35878
rect 26518 35876 26574 35878
rect 26278 34842 26334 34844
rect 26358 34842 26414 34844
rect 26438 34842 26494 34844
rect 26518 34842 26574 34844
rect 26278 34790 26324 34842
rect 26324 34790 26334 34842
rect 26358 34790 26388 34842
rect 26388 34790 26400 34842
rect 26400 34790 26414 34842
rect 26438 34790 26452 34842
rect 26452 34790 26464 34842
rect 26464 34790 26494 34842
rect 26518 34790 26528 34842
rect 26528 34790 26574 34842
rect 26278 34788 26334 34790
rect 26358 34788 26414 34790
rect 26438 34788 26494 34790
rect 26518 34788 26574 34790
rect 26278 33754 26334 33756
rect 26358 33754 26414 33756
rect 26438 33754 26494 33756
rect 26518 33754 26574 33756
rect 26278 33702 26324 33754
rect 26324 33702 26334 33754
rect 26358 33702 26388 33754
rect 26388 33702 26400 33754
rect 26400 33702 26414 33754
rect 26438 33702 26452 33754
rect 26452 33702 26464 33754
rect 26464 33702 26494 33754
rect 26518 33702 26528 33754
rect 26528 33702 26574 33754
rect 26278 33700 26334 33702
rect 26358 33700 26414 33702
rect 26438 33700 26494 33702
rect 26518 33700 26574 33702
rect 26278 32666 26334 32668
rect 26358 32666 26414 32668
rect 26438 32666 26494 32668
rect 26518 32666 26574 32668
rect 26278 32614 26324 32666
rect 26324 32614 26334 32666
rect 26358 32614 26388 32666
rect 26388 32614 26400 32666
rect 26400 32614 26414 32666
rect 26438 32614 26452 32666
rect 26452 32614 26464 32666
rect 26464 32614 26494 32666
rect 26518 32614 26528 32666
rect 26528 32614 26574 32666
rect 26278 32612 26334 32614
rect 26358 32612 26414 32614
rect 26438 32612 26494 32614
rect 26518 32612 26574 32614
rect 22058 29946 22114 29948
rect 22138 29946 22194 29948
rect 22218 29946 22274 29948
rect 22298 29946 22354 29948
rect 22058 29894 22104 29946
rect 22104 29894 22114 29946
rect 22138 29894 22168 29946
rect 22168 29894 22180 29946
rect 22180 29894 22194 29946
rect 22218 29894 22232 29946
rect 22232 29894 22244 29946
rect 22244 29894 22274 29946
rect 22298 29894 22308 29946
rect 22308 29894 22354 29946
rect 22058 29892 22114 29894
rect 22138 29892 22194 29894
rect 22218 29892 22274 29894
rect 22298 29892 22354 29894
rect 21086 26424 21142 26480
rect 5176 19066 5232 19068
rect 5256 19066 5312 19068
rect 5336 19066 5392 19068
rect 5416 19066 5472 19068
rect 5176 19014 5222 19066
rect 5222 19014 5232 19066
rect 5256 19014 5286 19066
rect 5286 19014 5298 19066
rect 5298 19014 5312 19066
rect 5336 19014 5350 19066
rect 5350 19014 5362 19066
rect 5362 19014 5392 19066
rect 5416 19014 5426 19066
rect 5426 19014 5472 19066
rect 5176 19012 5232 19014
rect 5256 19012 5312 19014
rect 5336 19012 5392 19014
rect 5416 19012 5472 19014
rect 13617 19066 13673 19068
rect 13697 19066 13753 19068
rect 13777 19066 13833 19068
rect 13857 19066 13913 19068
rect 13617 19014 13663 19066
rect 13663 19014 13673 19066
rect 13697 19014 13727 19066
rect 13727 19014 13739 19066
rect 13739 19014 13753 19066
rect 13777 19014 13791 19066
rect 13791 19014 13803 19066
rect 13803 19014 13833 19066
rect 13857 19014 13867 19066
rect 13867 19014 13913 19066
rect 13617 19012 13673 19014
rect 13697 19012 13753 19014
rect 13777 19012 13833 19014
rect 13857 19012 13913 19014
rect 9396 18522 9452 18524
rect 9476 18522 9532 18524
rect 9556 18522 9612 18524
rect 9636 18522 9692 18524
rect 9396 18470 9442 18522
rect 9442 18470 9452 18522
rect 9476 18470 9506 18522
rect 9506 18470 9518 18522
rect 9518 18470 9532 18522
rect 9556 18470 9570 18522
rect 9570 18470 9582 18522
rect 9582 18470 9612 18522
rect 9636 18470 9646 18522
rect 9646 18470 9692 18522
rect 9396 18468 9452 18470
rect 9476 18468 9532 18470
rect 9556 18468 9612 18470
rect 9636 18468 9692 18470
rect 17837 18522 17893 18524
rect 17917 18522 17973 18524
rect 17997 18522 18053 18524
rect 18077 18522 18133 18524
rect 17837 18470 17883 18522
rect 17883 18470 17893 18522
rect 17917 18470 17947 18522
rect 17947 18470 17959 18522
rect 17959 18470 17973 18522
rect 17997 18470 18011 18522
rect 18011 18470 18023 18522
rect 18023 18470 18053 18522
rect 18077 18470 18087 18522
rect 18087 18470 18133 18522
rect 17837 18468 17893 18470
rect 17917 18468 17973 18470
rect 17997 18468 18053 18470
rect 18077 18468 18133 18470
rect 5176 17978 5232 17980
rect 5256 17978 5312 17980
rect 5336 17978 5392 17980
rect 5416 17978 5472 17980
rect 5176 17926 5222 17978
rect 5222 17926 5232 17978
rect 5256 17926 5286 17978
rect 5286 17926 5298 17978
rect 5298 17926 5312 17978
rect 5336 17926 5350 17978
rect 5350 17926 5362 17978
rect 5362 17926 5392 17978
rect 5416 17926 5426 17978
rect 5426 17926 5472 17978
rect 5176 17924 5232 17926
rect 5256 17924 5312 17926
rect 5336 17924 5392 17926
rect 5416 17924 5472 17926
rect 13617 17978 13673 17980
rect 13697 17978 13753 17980
rect 13777 17978 13833 17980
rect 13857 17978 13913 17980
rect 13617 17926 13663 17978
rect 13663 17926 13673 17978
rect 13697 17926 13727 17978
rect 13727 17926 13739 17978
rect 13739 17926 13753 17978
rect 13777 17926 13791 17978
rect 13791 17926 13803 17978
rect 13803 17926 13833 17978
rect 13857 17926 13867 17978
rect 13867 17926 13913 17978
rect 13617 17924 13673 17926
rect 13697 17924 13753 17926
rect 13777 17924 13833 17926
rect 13857 17924 13913 17926
rect 9396 17434 9452 17436
rect 9476 17434 9532 17436
rect 9556 17434 9612 17436
rect 9636 17434 9692 17436
rect 9396 17382 9442 17434
rect 9442 17382 9452 17434
rect 9476 17382 9506 17434
rect 9506 17382 9518 17434
rect 9518 17382 9532 17434
rect 9556 17382 9570 17434
rect 9570 17382 9582 17434
rect 9582 17382 9612 17434
rect 9636 17382 9646 17434
rect 9646 17382 9692 17434
rect 9396 17380 9452 17382
rect 9476 17380 9532 17382
rect 9556 17380 9612 17382
rect 9636 17380 9692 17382
rect 17837 17434 17893 17436
rect 17917 17434 17973 17436
rect 17997 17434 18053 17436
rect 18077 17434 18133 17436
rect 17837 17382 17883 17434
rect 17883 17382 17893 17434
rect 17917 17382 17947 17434
rect 17947 17382 17959 17434
rect 17959 17382 17973 17434
rect 17997 17382 18011 17434
rect 18011 17382 18023 17434
rect 18023 17382 18053 17434
rect 18077 17382 18087 17434
rect 18087 17382 18133 17434
rect 17837 17380 17893 17382
rect 17917 17380 17973 17382
rect 17997 17380 18053 17382
rect 18077 17380 18133 17382
rect 5176 16890 5232 16892
rect 5256 16890 5312 16892
rect 5336 16890 5392 16892
rect 5416 16890 5472 16892
rect 5176 16838 5222 16890
rect 5222 16838 5232 16890
rect 5256 16838 5286 16890
rect 5286 16838 5298 16890
rect 5298 16838 5312 16890
rect 5336 16838 5350 16890
rect 5350 16838 5362 16890
rect 5362 16838 5392 16890
rect 5416 16838 5426 16890
rect 5426 16838 5472 16890
rect 5176 16836 5232 16838
rect 5256 16836 5312 16838
rect 5336 16836 5392 16838
rect 5416 16836 5472 16838
rect 13617 16890 13673 16892
rect 13697 16890 13753 16892
rect 13777 16890 13833 16892
rect 13857 16890 13913 16892
rect 13617 16838 13663 16890
rect 13663 16838 13673 16890
rect 13697 16838 13727 16890
rect 13727 16838 13739 16890
rect 13739 16838 13753 16890
rect 13777 16838 13791 16890
rect 13791 16838 13803 16890
rect 13803 16838 13833 16890
rect 13857 16838 13867 16890
rect 13867 16838 13913 16890
rect 13617 16836 13673 16838
rect 13697 16836 13753 16838
rect 13777 16836 13833 16838
rect 13857 16836 13913 16838
rect 9396 16346 9452 16348
rect 9476 16346 9532 16348
rect 9556 16346 9612 16348
rect 9636 16346 9692 16348
rect 9396 16294 9442 16346
rect 9442 16294 9452 16346
rect 9476 16294 9506 16346
rect 9506 16294 9518 16346
rect 9518 16294 9532 16346
rect 9556 16294 9570 16346
rect 9570 16294 9582 16346
rect 9582 16294 9612 16346
rect 9636 16294 9646 16346
rect 9646 16294 9692 16346
rect 9396 16292 9452 16294
rect 9476 16292 9532 16294
rect 9556 16292 9612 16294
rect 9636 16292 9692 16294
rect 17837 16346 17893 16348
rect 17917 16346 17973 16348
rect 17997 16346 18053 16348
rect 18077 16346 18133 16348
rect 17837 16294 17883 16346
rect 17883 16294 17893 16346
rect 17917 16294 17947 16346
rect 17947 16294 17959 16346
rect 17959 16294 17973 16346
rect 17997 16294 18011 16346
rect 18011 16294 18023 16346
rect 18023 16294 18053 16346
rect 18077 16294 18087 16346
rect 18087 16294 18133 16346
rect 17837 16292 17893 16294
rect 17917 16292 17973 16294
rect 17997 16292 18053 16294
rect 18077 16292 18133 16294
rect 5176 15802 5232 15804
rect 5256 15802 5312 15804
rect 5336 15802 5392 15804
rect 5416 15802 5472 15804
rect 5176 15750 5222 15802
rect 5222 15750 5232 15802
rect 5256 15750 5286 15802
rect 5286 15750 5298 15802
rect 5298 15750 5312 15802
rect 5336 15750 5350 15802
rect 5350 15750 5362 15802
rect 5362 15750 5392 15802
rect 5416 15750 5426 15802
rect 5426 15750 5472 15802
rect 5176 15748 5232 15750
rect 5256 15748 5312 15750
rect 5336 15748 5392 15750
rect 5416 15748 5472 15750
rect 13617 15802 13673 15804
rect 13697 15802 13753 15804
rect 13777 15802 13833 15804
rect 13857 15802 13913 15804
rect 13617 15750 13663 15802
rect 13663 15750 13673 15802
rect 13697 15750 13727 15802
rect 13727 15750 13739 15802
rect 13739 15750 13753 15802
rect 13777 15750 13791 15802
rect 13791 15750 13803 15802
rect 13803 15750 13833 15802
rect 13857 15750 13867 15802
rect 13867 15750 13913 15802
rect 13617 15748 13673 15750
rect 13697 15748 13753 15750
rect 13777 15748 13833 15750
rect 13857 15748 13913 15750
rect 9396 15258 9452 15260
rect 9476 15258 9532 15260
rect 9556 15258 9612 15260
rect 9636 15258 9692 15260
rect 9396 15206 9442 15258
rect 9442 15206 9452 15258
rect 9476 15206 9506 15258
rect 9506 15206 9518 15258
rect 9518 15206 9532 15258
rect 9556 15206 9570 15258
rect 9570 15206 9582 15258
rect 9582 15206 9612 15258
rect 9636 15206 9646 15258
rect 9646 15206 9692 15258
rect 9396 15204 9452 15206
rect 9476 15204 9532 15206
rect 9556 15204 9612 15206
rect 9636 15204 9692 15206
rect 17837 15258 17893 15260
rect 17917 15258 17973 15260
rect 17997 15258 18053 15260
rect 18077 15258 18133 15260
rect 17837 15206 17883 15258
rect 17883 15206 17893 15258
rect 17917 15206 17947 15258
rect 17947 15206 17959 15258
rect 17959 15206 17973 15258
rect 17997 15206 18011 15258
rect 18011 15206 18023 15258
rect 18023 15206 18053 15258
rect 18077 15206 18087 15258
rect 18087 15206 18133 15258
rect 17837 15204 17893 15206
rect 17917 15204 17973 15206
rect 17997 15204 18053 15206
rect 18077 15204 18133 15206
rect 5176 14714 5232 14716
rect 5256 14714 5312 14716
rect 5336 14714 5392 14716
rect 5416 14714 5472 14716
rect 5176 14662 5222 14714
rect 5222 14662 5232 14714
rect 5256 14662 5286 14714
rect 5286 14662 5298 14714
rect 5298 14662 5312 14714
rect 5336 14662 5350 14714
rect 5350 14662 5362 14714
rect 5362 14662 5392 14714
rect 5416 14662 5426 14714
rect 5426 14662 5472 14714
rect 5176 14660 5232 14662
rect 5256 14660 5312 14662
rect 5336 14660 5392 14662
rect 5416 14660 5472 14662
rect 13617 14714 13673 14716
rect 13697 14714 13753 14716
rect 13777 14714 13833 14716
rect 13857 14714 13913 14716
rect 13617 14662 13663 14714
rect 13663 14662 13673 14714
rect 13697 14662 13727 14714
rect 13727 14662 13739 14714
rect 13739 14662 13753 14714
rect 13777 14662 13791 14714
rect 13791 14662 13803 14714
rect 13803 14662 13833 14714
rect 13857 14662 13867 14714
rect 13867 14662 13913 14714
rect 13617 14660 13673 14662
rect 13697 14660 13753 14662
rect 13777 14660 13833 14662
rect 13857 14660 13913 14662
rect 938 14356 940 14376
rect 940 14356 992 14376
rect 992 14356 994 14376
rect 938 14320 994 14356
rect 9396 14170 9452 14172
rect 9476 14170 9532 14172
rect 9556 14170 9612 14172
rect 9636 14170 9692 14172
rect 9396 14118 9442 14170
rect 9442 14118 9452 14170
rect 9476 14118 9506 14170
rect 9506 14118 9518 14170
rect 9518 14118 9532 14170
rect 9556 14118 9570 14170
rect 9570 14118 9582 14170
rect 9582 14118 9612 14170
rect 9636 14118 9646 14170
rect 9646 14118 9692 14170
rect 9396 14116 9452 14118
rect 9476 14116 9532 14118
rect 9556 14116 9612 14118
rect 9636 14116 9692 14118
rect 17837 14170 17893 14172
rect 17917 14170 17973 14172
rect 17997 14170 18053 14172
rect 18077 14170 18133 14172
rect 17837 14118 17883 14170
rect 17883 14118 17893 14170
rect 17917 14118 17947 14170
rect 17947 14118 17959 14170
rect 17959 14118 17973 14170
rect 17997 14118 18011 14170
rect 18011 14118 18023 14170
rect 18023 14118 18053 14170
rect 18077 14118 18087 14170
rect 18087 14118 18133 14170
rect 17837 14116 17893 14118
rect 17917 14116 17973 14118
rect 17997 14116 18053 14118
rect 18077 14116 18133 14118
rect 5176 13626 5232 13628
rect 5256 13626 5312 13628
rect 5336 13626 5392 13628
rect 5416 13626 5472 13628
rect 5176 13574 5222 13626
rect 5222 13574 5232 13626
rect 5256 13574 5286 13626
rect 5286 13574 5298 13626
rect 5298 13574 5312 13626
rect 5336 13574 5350 13626
rect 5350 13574 5362 13626
rect 5362 13574 5392 13626
rect 5416 13574 5426 13626
rect 5426 13574 5472 13626
rect 5176 13572 5232 13574
rect 5256 13572 5312 13574
rect 5336 13572 5392 13574
rect 5416 13572 5472 13574
rect 13617 13626 13673 13628
rect 13697 13626 13753 13628
rect 13777 13626 13833 13628
rect 13857 13626 13913 13628
rect 13617 13574 13663 13626
rect 13663 13574 13673 13626
rect 13697 13574 13727 13626
rect 13727 13574 13739 13626
rect 13739 13574 13753 13626
rect 13777 13574 13791 13626
rect 13791 13574 13803 13626
rect 13803 13574 13833 13626
rect 13857 13574 13867 13626
rect 13867 13574 13913 13626
rect 13617 13572 13673 13574
rect 13697 13572 13753 13574
rect 13777 13572 13833 13574
rect 13857 13572 13913 13574
rect 9396 13082 9452 13084
rect 9476 13082 9532 13084
rect 9556 13082 9612 13084
rect 9636 13082 9692 13084
rect 9396 13030 9442 13082
rect 9442 13030 9452 13082
rect 9476 13030 9506 13082
rect 9506 13030 9518 13082
rect 9518 13030 9532 13082
rect 9556 13030 9570 13082
rect 9570 13030 9582 13082
rect 9582 13030 9612 13082
rect 9636 13030 9646 13082
rect 9646 13030 9692 13082
rect 9396 13028 9452 13030
rect 9476 13028 9532 13030
rect 9556 13028 9612 13030
rect 9636 13028 9692 13030
rect 17837 13082 17893 13084
rect 17917 13082 17973 13084
rect 17997 13082 18053 13084
rect 18077 13082 18133 13084
rect 17837 13030 17883 13082
rect 17883 13030 17893 13082
rect 17917 13030 17947 13082
rect 17947 13030 17959 13082
rect 17959 13030 17973 13082
rect 17997 13030 18011 13082
rect 18011 13030 18023 13082
rect 18023 13030 18053 13082
rect 18077 13030 18087 13082
rect 18087 13030 18133 13082
rect 17837 13028 17893 13030
rect 17917 13028 17973 13030
rect 17997 13028 18053 13030
rect 18077 13028 18133 13030
rect 5176 12538 5232 12540
rect 5256 12538 5312 12540
rect 5336 12538 5392 12540
rect 5416 12538 5472 12540
rect 5176 12486 5222 12538
rect 5222 12486 5232 12538
rect 5256 12486 5286 12538
rect 5286 12486 5298 12538
rect 5298 12486 5312 12538
rect 5336 12486 5350 12538
rect 5350 12486 5362 12538
rect 5362 12486 5392 12538
rect 5416 12486 5426 12538
rect 5426 12486 5472 12538
rect 5176 12484 5232 12486
rect 5256 12484 5312 12486
rect 5336 12484 5392 12486
rect 5416 12484 5472 12486
rect 13617 12538 13673 12540
rect 13697 12538 13753 12540
rect 13777 12538 13833 12540
rect 13857 12538 13913 12540
rect 13617 12486 13663 12538
rect 13663 12486 13673 12538
rect 13697 12486 13727 12538
rect 13727 12486 13739 12538
rect 13739 12486 13753 12538
rect 13777 12486 13791 12538
rect 13791 12486 13803 12538
rect 13803 12486 13833 12538
rect 13857 12486 13867 12538
rect 13867 12486 13913 12538
rect 13617 12484 13673 12486
rect 13697 12484 13753 12486
rect 13777 12484 13833 12486
rect 13857 12484 13913 12486
rect 20534 23160 20590 23216
rect 22058 28858 22114 28860
rect 22138 28858 22194 28860
rect 22218 28858 22274 28860
rect 22298 28858 22354 28860
rect 22058 28806 22104 28858
rect 22104 28806 22114 28858
rect 22138 28806 22168 28858
rect 22168 28806 22180 28858
rect 22180 28806 22194 28858
rect 22218 28806 22232 28858
rect 22232 28806 22244 28858
rect 22244 28806 22274 28858
rect 22298 28806 22308 28858
rect 22308 28806 22354 28858
rect 22058 28804 22114 28806
rect 22138 28804 22194 28806
rect 22218 28804 22274 28806
rect 22298 28804 22354 28806
rect 26278 31578 26334 31580
rect 26358 31578 26414 31580
rect 26438 31578 26494 31580
rect 26518 31578 26574 31580
rect 26278 31526 26324 31578
rect 26324 31526 26334 31578
rect 26358 31526 26388 31578
rect 26388 31526 26400 31578
rect 26400 31526 26414 31578
rect 26438 31526 26452 31578
rect 26452 31526 26464 31578
rect 26464 31526 26494 31578
rect 26518 31526 26528 31578
rect 26528 31526 26574 31578
rect 26278 31524 26334 31526
rect 26358 31524 26414 31526
rect 26438 31524 26494 31526
rect 26518 31524 26574 31526
rect 26278 30490 26334 30492
rect 26358 30490 26414 30492
rect 26438 30490 26494 30492
rect 26518 30490 26574 30492
rect 26278 30438 26324 30490
rect 26324 30438 26334 30490
rect 26358 30438 26388 30490
rect 26388 30438 26400 30490
rect 26400 30438 26414 30490
rect 26438 30438 26452 30490
rect 26452 30438 26464 30490
rect 26464 30438 26494 30490
rect 26518 30438 26528 30490
rect 26528 30438 26574 30490
rect 26278 30436 26334 30438
rect 26358 30436 26414 30438
rect 26438 30436 26494 30438
rect 26518 30436 26574 30438
rect 30499 39738 30555 39740
rect 30579 39738 30635 39740
rect 30659 39738 30715 39740
rect 30739 39738 30795 39740
rect 30499 39686 30545 39738
rect 30545 39686 30555 39738
rect 30579 39686 30609 39738
rect 30609 39686 30621 39738
rect 30621 39686 30635 39738
rect 30659 39686 30673 39738
rect 30673 39686 30685 39738
rect 30685 39686 30715 39738
rect 30739 39686 30749 39738
rect 30749 39686 30795 39738
rect 30499 39684 30555 39686
rect 30579 39684 30635 39686
rect 30659 39684 30715 39686
rect 30739 39684 30795 39686
rect 34719 39194 34775 39196
rect 34799 39194 34855 39196
rect 34879 39194 34935 39196
rect 34959 39194 35015 39196
rect 34719 39142 34765 39194
rect 34765 39142 34775 39194
rect 34799 39142 34829 39194
rect 34829 39142 34841 39194
rect 34841 39142 34855 39194
rect 34879 39142 34893 39194
rect 34893 39142 34905 39194
rect 34905 39142 34935 39194
rect 34959 39142 34969 39194
rect 34969 39142 35015 39194
rect 34719 39140 34775 39142
rect 34799 39140 34855 39142
rect 34879 39140 34935 39142
rect 34959 39140 35015 39142
rect 30499 38650 30555 38652
rect 30579 38650 30635 38652
rect 30659 38650 30715 38652
rect 30739 38650 30795 38652
rect 30499 38598 30545 38650
rect 30545 38598 30555 38650
rect 30579 38598 30609 38650
rect 30609 38598 30621 38650
rect 30621 38598 30635 38650
rect 30659 38598 30673 38650
rect 30673 38598 30685 38650
rect 30685 38598 30715 38650
rect 30739 38598 30749 38650
rect 30749 38598 30795 38650
rect 30499 38596 30555 38598
rect 30579 38596 30635 38598
rect 30659 38596 30715 38598
rect 30739 38596 30795 38598
rect 34719 38106 34775 38108
rect 34799 38106 34855 38108
rect 34879 38106 34935 38108
rect 34959 38106 35015 38108
rect 34719 38054 34765 38106
rect 34765 38054 34775 38106
rect 34799 38054 34829 38106
rect 34829 38054 34841 38106
rect 34841 38054 34855 38106
rect 34879 38054 34893 38106
rect 34893 38054 34905 38106
rect 34905 38054 34935 38106
rect 34959 38054 34969 38106
rect 34969 38054 35015 38106
rect 34719 38052 34775 38054
rect 34799 38052 34855 38054
rect 34879 38052 34935 38054
rect 34959 38052 35015 38054
rect 30499 37562 30555 37564
rect 30579 37562 30635 37564
rect 30659 37562 30715 37564
rect 30739 37562 30795 37564
rect 30499 37510 30545 37562
rect 30545 37510 30555 37562
rect 30579 37510 30609 37562
rect 30609 37510 30621 37562
rect 30621 37510 30635 37562
rect 30659 37510 30673 37562
rect 30673 37510 30685 37562
rect 30685 37510 30715 37562
rect 30739 37510 30749 37562
rect 30749 37510 30795 37562
rect 30499 37508 30555 37510
rect 30579 37508 30635 37510
rect 30659 37508 30715 37510
rect 30739 37508 30795 37510
rect 34719 37018 34775 37020
rect 34799 37018 34855 37020
rect 34879 37018 34935 37020
rect 34959 37018 35015 37020
rect 34719 36966 34765 37018
rect 34765 36966 34775 37018
rect 34799 36966 34829 37018
rect 34829 36966 34841 37018
rect 34841 36966 34855 37018
rect 34879 36966 34893 37018
rect 34893 36966 34905 37018
rect 34905 36966 34935 37018
rect 34959 36966 34969 37018
rect 34969 36966 35015 37018
rect 34719 36964 34775 36966
rect 34799 36964 34855 36966
rect 34879 36964 34935 36966
rect 34959 36964 35015 36966
rect 30499 36474 30555 36476
rect 30579 36474 30635 36476
rect 30659 36474 30715 36476
rect 30739 36474 30795 36476
rect 30499 36422 30545 36474
rect 30545 36422 30555 36474
rect 30579 36422 30609 36474
rect 30609 36422 30621 36474
rect 30621 36422 30635 36474
rect 30659 36422 30673 36474
rect 30673 36422 30685 36474
rect 30685 36422 30715 36474
rect 30739 36422 30749 36474
rect 30749 36422 30795 36474
rect 30499 36420 30555 36422
rect 30579 36420 30635 36422
rect 30659 36420 30715 36422
rect 30739 36420 30795 36422
rect 34719 35930 34775 35932
rect 34799 35930 34855 35932
rect 34879 35930 34935 35932
rect 34959 35930 35015 35932
rect 34719 35878 34765 35930
rect 34765 35878 34775 35930
rect 34799 35878 34829 35930
rect 34829 35878 34841 35930
rect 34841 35878 34855 35930
rect 34879 35878 34893 35930
rect 34893 35878 34905 35930
rect 34905 35878 34935 35930
rect 34959 35878 34969 35930
rect 34969 35878 35015 35930
rect 34719 35876 34775 35878
rect 34799 35876 34855 35878
rect 34879 35876 34935 35878
rect 34959 35876 35015 35878
rect 30499 35386 30555 35388
rect 30579 35386 30635 35388
rect 30659 35386 30715 35388
rect 30739 35386 30795 35388
rect 30499 35334 30545 35386
rect 30545 35334 30555 35386
rect 30579 35334 30609 35386
rect 30609 35334 30621 35386
rect 30621 35334 30635 35386
rect 30659 35334 30673 35386
rect 30673 35334 30685 35386
rect 30685 35334 30715 35386
rect 30739 35334 30749 35386
rect 30749 35334 30795 35386
rect 30499 35332 30555 35334
rect 30579 35332 30635 35334
rect 30659 35332 30715 35334
rect 30739 35332 30795 35334
rect 34719 34842 34775 34844
rect 34799 34842 34855 34844
rect 34879 34842 34935 34844
rect 34959 34842 35015 34844
rect 34719 34790 34765 34842
rect 34765 34790 34775 34842
rect 34799 34790 34829 34842
rect 34829 34790 34841 34842
rect 34841 34790 34855 34842
rect 34879 34790 34893 34842
rect 34893 34790 34905 34842
rect 34905 34790 34935 34842
rect 34959 34790 34969 34842
rect 34969 34790 35015 34842
rect 34719 34788 34775 34790
rect 34799 34788 34855 34790
rect 34879 34788 34935 34790
rect 34959 34788 35015 34790
rect 35162 34720 35218 34776
rect 30499 34298 30555 34300
rect 30579 34298 30635 34300
rect 30659 34298 30715 34300
rect 30739 34298 30795 34300
rect 30499 34246 30545 34298
rect 30545 34246 30555 34298
rect 30579 34246 30609 34298
rect 30609 34246 30621 34298
rect 30621 34246 30635 34298
rect 30659 34246 30673 34298
rect 30673 34246 30685 34298
rect 30685 34246 30715 34298
rect 30739 34246 30749 34298
rect 30749 34246 30795 34298
rect 30499 34244 30555 34246
rect 30579 34244 30635 34246
rect 30659 34244 30715 34246
rect 30739 34244 30795 34246
rect 34719 33754 34775 33756
rect 34799 33754 34855 33756
rect 34879 33754 34935 33756
rect 34959 33754 35015 33756
rect 34719 33702 34765 33754
rect 34765 33702 34775 33754
rect 34799 33702 34829 33754
rect 34829 33702 34841 33754
rect 34841 33702 34855 33754
rect 34879 33702 34893 33754
rect 34893 33702 34905 33754
rect 34905 33702 34935 33754
rect 34959 33702 34969 33754
rect 34969 33702 35015 33754
rect 34719 33700 34775 33702
rect 34799 33700 34855 33702
rect 34879 33700 34935 33702
rect 34959 33700 35015 33702
rect 30499 33210 30555 33212
rect 30579 33210 30635 33212
rect 30659 33210 30715 33212
rect 30739 33210 30795 33212
rect 30499 33158 30545 33210
rect 30545 33158 30555 33210
rect 30579 33158 30609 33210
rect 30609 33158 30621 33210
rect 30621 33158 30635 33210
rect 30659 33158 30673 33210
rect 30673 33158 30685 33210
rect 30685 33158 30715 33210
rect 30739 33158 30749 33210
rect 30749 33158 30795 33210
rect 30499 33156 30555 33158
rect 30579 33156 30635 33158
rect 30659 33156 30715 33158
rect 30739 33156 30795 33158
rect 34719 32666 34775 32668
rect 34799 32666 34855 32668
rect 34879 32666 34935 32668
rect 34959 32666 35015 32668
rect 34719 32614 34765 32666
rect 34765 32614 34775 32666
rect 34799 32614 34829 32666
rect 34829 32614 34841 32666
rect 34841 32614 34855 32666
rect 34879 32614 34893 32666
rect 34893 32614 34905 32666
rect 34905 32614 34935 32666
rect 34959 32614 34969 32666
rect 34969 32614 35015 32666
rect 34719 32612 34775 32614
rect 34799 32612 34855 32614
rect 34879 32612 34935 32614
rect 34959 32612 35015 32614
rect 30499 32122 30555 32124
rect 30579 32122 30635 32124
rect 30659 32122 30715 32124
rect 30739 32122 30795 32124
rect 30499 32070 30545 32122
rect 30545 32070 30555 32122
rect 30579 32070 30609 32122
rect 30609 32070 30621 32122
rect 30621 32070 30635 32122
rect 30659 32070 30673 32122
rect 30673 32070 30685 32122
rect 30685 32070 30715 32122
rect 30739 32070 30749 32122
rect 30749 32070 30795 32122
rect 30499 32068 30555 32070
rect 30579 32068 30635 32070
rect 30659 32068 30715 32070
rect 30739 32068 30795 32070
rect 34719 31578 34775 31580
rect 34799 31578 34855 31580
rect 34879 31578 34935 31580
rect 34959 31578 35015 31580
rect 34719 31526 34765 31578
rect 34765 31526 34775 31578
rect 34799 31526 34829 31578
rect 34829 31526 34841 31578
rect 34841 31526 34855 31578
rect 34879 31526 34893 31578
rect 34893 31526 34905 31578
rect 34905 31526 34935 31578
rect 34959 31526 34969 31578
rect 34969 31526 35015 31578
rect 34719 31524 34775 31526
rect 34799 31524 34855 31526
rect 34879 31524 34935 31526
rect 34959 31524 35015 31526
rect 30499 31034 30555 31036
rect 30579 31034 30635 31036
rect 30659 31034 30715 31036
rect 30739 31034 30795 31036
rect 30499 30982 30545 31034
rect 30545 30982 30555 31034
rect 30579 30982 30609 31034
rect 30609 30982 30621 31034
rect 30621 30982 30635 31034
rect 30659 30982 30673 31034
rect 30673 30982 30685 31034
rect 30685 30982 30715 31034
rect 30739 30982 30749 31034
rect 30749 30982 30795 31034
rect 30499 30980 30555 30982
rect 30579 30980 30635 30982
rect 30659 30980 30715 30982
rect 30739 30980 30795 30982
rect 34719 30490 34775 30492
rect 34799 30490 34855 30492
rect 34879 30490 34935 30492
rect 34959 30490 35015 30492
rect 34719 30438 34765 30490
rect 34765 30438 34775 30490
rect 34799 30438 34829 30490
rect 34829 30438 34841 30490
rect 34841 30438 34855 30490
rect 34879 30438 34893 30490
rect 34893 30438 34905 30490
rect 34905 30438 34935 30490
rect 34959 30438 34969 30490
rect 34969 30438 35015 30490
rect 34719 30436 34775 30438
rect 34799 30436 34855 30438
rect 34879 30436 34935 30438
rect 34959 30436 35015 30438
rect 30499 29946 30555 29948
rect 30579 29946 30635 29948
rect 30659 29946 30715 29948
rect 30739 29946 30795 29948
rect 30499 29894 30545 29946
rect 30545 29894 30555 29946
rect 30579 29894 30609 29946
rect 30609 29894 30621 29946
rect 30621 29894 30635 29946
rect 30659 29894 30673 29946
rect 30673 29894 30685 29946
rect 30685 29894 30715 29946
rect 30739 29894 30749 29946
rect 30749 29894 30795 29946
rect 30499 29892 30555 29894
rect 30579 29892 30635 29894
rect 30659 29892 30715 29894
rect 30739 29892 30795 29894
rect 26278 29402 26334 29404
rect 26358 29402 26414 29404
rect 26438 29402 26494 29404
rect 26518 29402 26574 29404
rect 26278 29350 26324 29402
rect 26324 29350 26334 29402
rect 26358 29350 26388 29402
rect 26388 29350 26400 29402
rect 26400 29350 26414 29402
rect 26438 29350 26452 29402
rect 26452 29350 26464 29402
rect 26464 29350 26494 29402
rect 26518 29350 26528 29402
rect 26528 29350 26574 29402
rect 26278 29348 26334 29350
rect 26358 29348 26414 29350
rect 26438 29348 26494 29350
rect 26518 29348 26574 29350
rect 34719 29402 34775 29404
rect 34799 29402 34855 29404
rect 34879 29402 34935 29404
rect 34959 29402 35015 29404
rect 34719 29350 34765 29402
rect 34765 29350 34775 29402
rect 34799 29350 34829 29402
rect 34829 29350 34841 29402
rect 34841 29350 34855 29402
rect 34879 29350 34893 29402
rect 34893 29350 34905 29402
rect 34905 29350 34935 29402
rect 34959 29350 34969 29402
rect 34969 29350 35015 29402
rect 34719 29348 34775 29350
rect 34799 29348 34855 29350
rect 34879 29348 34935 29350
rect 34959 29348 35015 29350
rect 22058 27770 22114 27772
rect 22138 27770 22194 27772
rect 22218 27770 22274 27772
rect 22298 27770 22354 27772
rect 22058 27718 22104 27770
rect 22104 27718 22114 27770
rect 22138 27718 22168 27770
rect 22168 27718 22180 27770
rect 22180 27718 22194 27770
rect 22218 27718 22232 27770
rect 22232 27718 22244 27770
rect 22244 27718 22274 27770
rect 22298 27718 22308 27770
rect 22308 27718 22354 27770
rect 22058 27716 22114 27718
rect 22138 27716 22194 27718
rect 22218 27716 22274 27718
rect 22298 27716 22354 27718
rect 21730 27104 21786 27160
rect 22058 26682 22114 26684
rect 22138 26682 22194 26684
rect 22218 26682 22274 26684
rect 22298 26682 22354 26684
rect 22058 26630 22104 26682
rect 22104 26630 22114 26682
rect 22138 26630 22168 26682
rect 22168 26630 22180 26682
rect 22180 26630 22194 26682
rect 22218 26630 22232 26682
rect 22232 26630 22244 26682
rect 22244 26630 22274 26682
rect 22298 26630 22308 26682
rect 22308 26630 22354 26682
rect 22058 26628 22114 26630
rect 22138 26628 22194 26630
rect 22218 26628 22274 26630
rect 22298 26628 22354 26630
rect 22058 25594 22114 25596
rect 22138 25594 22194 25596
rect 22218 25594 22274 25596
rect 22298 25594 22354 25596
rect 22058 25542 22104 25594
rect 22104 25542 22114 25594
rect 22138 25542 22168 25594
rect 22168 25542 22180 25594
rect 22180 25542 22194 25594
rect 22218 25542 22232 25594
rect 22232 25542 22244 25594
rect 22244 25542 22274 25594
rect 22298 25542 22308 25594
rect 22308 25542 22354 25594
rect 22058 25540 22114 25542
rect 22138 25540 22194 25542
rect 22218 25540 22274 25542
rect 22298 25540 22354 25542
rect 20810 22888 20866 22944
rect 22058 24506 22114 24508
rect 22138 24506 22194 24508
rect 22218 24506 22274 24508
rect 22298 24506 22354 24508
rect 22058 24454 22104 24506
rect 22104 24454 22114 24506
rect 22138 24454 22168 24506
rect 22168 24454 22180 24506
rect 22180 24454 22194 24506
rect 22218 24454 22232 24506
rect 22232 24454 22244 24506
rect 22244 24454 22274 24506
rect 22298 24454 22308 24506
rect 22308 24454 22354 24506
rect 22058 24452 22114 24454
rect 22138 24452 22194 24454
rect 22218 24452 22274 24454
rect 22298 24452 22354 24454
rect 30499 28858 30555 28860
rect 30579 28858 30635 28860
rect 30659 28858 30715 28860
rect 30739 28858 30795 28860
rect 30499 28806 30545 28858
rect 30545 28806 30555 28858
rect 30579 28806 30609 28858
rect 30609 28806 30621 28858
rect 30621 28806 30635 28858
rect 30659 28806 30673 28858
rect 30673 28806 30685 28858
rect 30685 28806 30715 28858
rect 30739 28806 30749 28858
rect 30749 28806 30795 28858
rect 30499 28804 30555 28806
rect 30579 28804 30635 28806
rect 30659 28804 30715 28806
rect 30739 28804 30795 28806
rect 26278 28314 26334 28316
rect 26358 28314 26414 28316
rect 26438 28314 26494 28316
rect 26518 28314 26574 28316
rect 26278 28262 26324 28314
rect 26324 28262 26334 28314
rect 26358 28262 26388 28314
rect 26388 28262 26400 28314
rect 26400 28262 26414 28314
rect 26438 28262 26452 28314
rect 26452 28262 26464 28314
rect 26464 28262 26494 28314
rect 26518 28262 26528 28314
rect 26528 28262 26574 28314
rect 26278 28260 26334 28262
rect 26358 28260 26414 28262
rect 26438 28260 26494 28262
rect 26518 28260 26574 28262
rect 34719 28314 34775 28316
rect 34799 28314 34855 28316
rect 34879 28314 34935 28316
rect 34959 28314 35015 28316
rect 34719 28262 34765 28314
rect 34765 28262 34775 28314
rect 34799 28262 34829 28314
rect 34829 28262 34841 28314
rect 34841 28262 34855 28314
rect 34879 28262 34893 28314
rect 34893 28262 34905 28314
rect 34905 28262 34935 28314
rect 34959 28262 34969 28314
rect 34969 28262 35015 28314
rect 34719 28260 34775 28262
rect 34799 28260 34855 28262
rect 34879 28260 34935 28262
rect 34959 28260 35015 28262
rect 30499 27770 30555 27772
rect 30579 27770 30635 27772
rect 30659 27770 30715 27772
rect 30739 27770 30795 27772
rect 30499 27718 30545 27770
rect 30545 27718 30555 27770
rect 30579 27718 30609 27770
rect 30609 27718 30621 27770
rect 30621 27718 30635 27770
rect 30659 27718 30673 27770
rect 30673 27718 30685 27770
rect 30685 27718 30715 27770
rect 30739 27718 30749 27770
rect 30749 27718 30795 27770
rect 30499 27716 30555 27718
rect 30579 27716 30635 27718
rect 30659 27716 30715 27718
rect 30739 27716 30795 27718
rect 22282 23568 22338 23624
rect 22058 23418 22114 23420
rect 22138 23418 22194 23420
rect 22218 23418 22274 23420
rect 22298 23418 22354 23420
rect 22058 23366 22104 23418
rect 22104 23366 22114 23418
rect 22138 23366 22168 23418
rect 22168 23366 22180 23418
rect 22180 23366 22194 23418
rect 22218 23366 22232 23418
rect 22232 23366 22244 23418
rect 22244 23366 22274 23418
rect 22298 23366 22308 23418
rect 22308 23366 22354 23418
rect 22058 23364 22114 23366
rect 22138 23364 22194 23366
rect 22218 23364 22274 23366
rect 22298 23364 22354 23366
rect 22006 22772 22062 22808
rect 22006 22752 22008 22772
rect 22008 22752 22060 22772
rect 22060 22752 22062 22772
rect 22374 22888 22430 22944
rect 23018 23568 23074 23624
rect 22058 22330 22114 22332
rect 22138 22330 22194 22332
rect 22218 22330 22274 22332
rect 22298 22330 22354 22332
rect 22058 22278 22104 22330
rect 22104 22278 22114 22330
rect 22138 22278 22168 22330
rect 22168 22278 22180 22330
rect 22180 22278 22194 22330
rect 22218 22278 22232 22330
rect 22232 22278 22244 22330
rect 22244 22278 22274 22330
rect 22298 22278 22308 22330
rect 22308 22278 22354 22330
rect 22058 22276 22114 22278
rect 22138 22276 22194 22278
rect 22218 22276 22274 22278
rect 22298 22276 22354 22278
rect 22058 21242 22114 21244
rect 22138 21242 22194 21244
rect 22218 21242 22274 21244
rect 22298 21242 22354 21244
rect 22058 21190 22104 21242
rect 22104 21190 22114 21242
rect 22138 21190 22168 21242
rect 22168 21190 22180 21242
rect 22180 21190 22194 21242
rect 22218 21190 22232 21242
rect 22232 21190 22244 21242
rect 22244 21190 22274 21242
rect 22298 21190 22308 21242
rect 22308 21190 22354 21242
rect 22058 21188 22114 21190
rect 22138 21188 22194 21190
rect 22218 21188 22274 21190
rect 22298 21188 22354 21190
rect 22058 20154 22114 20156
rect 22138 20154 22194 20156
rect 22218 20154 22274 20156
rect 22298 20154 22354 20156
rect 22058 20102 22104 20154
rect 22104 20102 22114 20154
rect 22138 20102 22168 20154
rect 22168 20102 22180 20154
rect 22180 20102 22194 20154
rect 22218 20102 22232 20154
rect 22232 20102 22244 20154
rect 22244 20102 22274 20154
rect 22298 20102 22308 20154
rect 22308 20102 22354 20154
rect 22058 20100 22114 20102
rect 22138 20100 22194 20102
rect 22218 20100 22274 20102
rect 22298 20100 22354 20102
rect 23846 22752 23902 22808
rect 22058 19066 22114 19068
rect 22138 19066 22194 19068
rect 22218 19066 22274 19068
rect 22298 19066 22354 19068
rect 22058 19014 22104 19066
rect 22104 19014 22114 19066
rect 22138 19014 22168 19066
rect 22168 19014 22180 19066
rect 22180 19014 22194 19066
rect 22218 19014 22232 19066
rect 22232 19014 22244 19066
rect 22244 19014 22274 19066
rect 22298 19014 22308 19066
rect 22308 19014 22354 19066
rect 22058 19012 22114 19014
rect 22138 19012 22194 19014
rect 22218 19012 22274 19014
rect 22298 19012 22354 19014
rect 22058 17978 22114 17980
rect 22138 17978 22194 17980
rect 22218 17978 22274 17980
rect 22298 17978 22354 17980
rect 22058 17926 22104 17978
rect 22104 17926 22114 17978
rect 22138 17926 22168 17978
rect 22168 17926 22180 17978
rect 22180 17926 22194 17978
rect 22218 17926 22232 17978
rect 22232 17926 22244 17978
rect 22244 17926 22274 17978
rect 22298 17926 22308 17978
rect 22308 17926 22354 17978
rect 22058 17924 22114 17926
rect 22138 17924 22194 17926
rect 22218 17924 22274 17926
rect 22298 17924 22354 17926
rect 22058 16890 22114 16892
rect 22138 16890 22194 16892
rect 22218 16890 22274 16892
rect 22298 16890 22354 16892
rect 22058 16838 22104 16890
rect 22104 16838 22114 16890
rect 22138 16838 22168 16890
rect 22168 16838 22180 16890
rect 22180 16838 22194 16890
rect 22218 16838 22232 16890
rect 22232 16838 22244 16890
rect 22244 16838 22274 16890
rect 22298 16838 22308 16890
rect 22308 16838 22354 16890
rect 22058 16836 22114 16838
rect 22138 16836 22194 16838
rect 22218 16836 22274 16838
rect 22298 16836 22354 16838
rect 22058 15802 22114 15804
rect 22138 15802 22194 15804
rect 22218 15802 22274 15804
rect 22298 15802 22354 15804
rect 22058 15750 22104 15802
rect 22104 15750 22114 15802
rect 22138 15750 22168 15802
rect 22168 15750 22180 15802
rect 22180 15750 22194 15802
rect 22218 15750 22232 15802
rect 22232 15750 22244 15802
rect 22244 15750 22274 15802
rect 22298 15750 22308 15802
rect 22308 15750 22354 15802
rect 22058 15748 22114 15750
rect 22138 15748 22194 15750
rect 22218 15748 22274 15750
rect 22298 15748 22354 15750
rect 22058 14714 22114 14716
rect 22138 14714 22194 14716
rect 22218 14714 22274 14716
rect 22298 14714 22354 14716
rect 22058 14662 22104 14714
rect 22104 14662 22114 14714
rect 22138 14662 22168 14714
rect 22168 14662 22180 14714
rect 22180 14662 22194 14714
rect 22218 14662 22232 14714
rect 22232 14662 22244 14714
rect 22244 14662 22274 14714
rect 22298 14662 22308 14714
rect 22308 14662 22354 14714
rect 22058 14660 22114 14662
rect 22138 14660 22194 14662
rect 22218 14660 22274 14662
rect 22298 14660 22354 14662
rect 22058 13626 22114 13628
rect 22138 13626 22194 13628
rect 22218 13626 22274 13628
rect 22298 13626 22354 13628
rect 22058 13574 22104 13626
rect 22104 13574 22114 13626
rect 22138 13574 22168 13626
rect 22168 13574 22180 13626
rect 22180 13574 22194 13626
rect 22218 13574 22232 13626
rect 22232 13574 22244 13626
rect 22244 13574 22274 13626
rect 22298 13574 22308 13626
rect 22308 13574 22354 13626
rect 22058 13572 22114 13574
rect 22138 13572 22194 13574
rect 22218 13572 22274 13574
rect 22298 13572 22354 13574
rect 34518 27412 34520 27432
rect 34520 27412 34572 27432
rect 34572 27412 34574 27432
rect 34518 27376 34574 27412
rect 26278 27226 26334 27228
rect 26358 27226 26414 27228
rect 26438 27226 26494 27228
rect 26518 27226 26574 27228
rect 26278 27174 26324 27226
rect 26324 27174 26334 27226
rect 26358 27174 26388 27226
rect 26388 27174 26400 27226
rect 26400 27174 26414 27226
rect 26438 27174 26452 27226
rect 26452 27174 26464 27226
rect 26464 27174 26494 27226
rect 26518 27174 26528 27226
rect 26528 27174 26574 27226
rect 26278 27172 26334 27174
rect 26358 27172 26414 27174
rect 26438 27172 26494 27174
rect 26518 27172 26574 27174
rect 34719 27226 34775 27228
rect 34799 27226 34855 27228
rect 34879 27226 34935 27228
rect 34959 27226 35015 27228
rect 34719 27174 34765 27226
rect 34765 27174 34775 27226
rect 34799 27174 34829 27226
rect 34829 27174 34841 27226
rect 34841 27174 34855 27226
rect 34879 27174 34893 27226
rect 34893 27174 34905 27226
rect 34905 27174 34935 27226
rect 34959 27174 34969 27226
rect 34969 27174 35015 27226
rect 34719 27172 34775 27174
rect 34799 27172 34855 27174
rect 34879 27172 34935 27174
rect 34959 27172 35015 27174
rect 30499 26682 30555 26684
rect 30579 26682 30635 26684
rect 30659 26682 30715 26684
rect 30739 26682 30795 26684
rect 30499 26630 30545 26682
rect 30545 26630 30555 26682
rect 30579 26630 30609 26682
rect 30609 26630 30621 26682
rect 30621 26630 30635 26682
rect 30659 26630 30673 26682
rect 30673 26630 30685 26682
rect 30685 26630 30715 26682
rect 30739 26630 30749 26682
rect 30749 26630 30795 26682
rect 30499 26628 30555 26630
rect 30579 26628 30635 26630
rect 30659 26628 30715 26630
rect 30739 26628 30795 26630
rect 24582 26424 24638 26480
rect 26278 26138 26334 26140
rect 26358 26138 26414 26140
rect 26438 26138 26494 26140
rect 26518 26138 26574 26140
rect 26278 26086 26324 26138
rect 26324 26086 26334 26138
rect 26358 26086 26388 26138
rect 26388 26086 26400 26138
rect 26400 26086 26414 26138
rect 26438 26086 26452 26138
rect 26452 26086 26464 26138
rect 26464 26086 26494 26138
rect 26518 26086 26528 26138
rect 26528 26086 26574 26138
rect 26278 26084 26334 26086
rect 26358 26084 26414 26086
rect 26438 26084 26494 26086
rect 26518 26084 26574 26086
rect 34719 26138 34775 26140
rect 34799 26138 34855 26140
rect 34879 26138 34935 26140
rect 34959 26138 35015 26140
rect 34719 26086 34765 26138
rect 34765 26086 34775 26138
rect 34799 26086 34829 26138
rect 34829 26086 34841 26138
rect 34841 26086 34855 26138
rect 34879 26086 34893 26138
rect 34893 26086 34905 26138
rect 34905 26086 34935 26138
rect 34959 26086 34969 26138
rect 34969 26086 35015 26138
rect 34719 26084 34775 26086
rect 34799 26084 34855 26086
rect 34879 26084 34935 26086
rect 34959 26084 35015 26086
rect 30499 25594 30555 25596
rect 30579 25594 30635 25596
rect 30659 25594 30715 25596
rect 30739 25594 30795 25596
rect 30499 25542 30545 25594
rect 30545 25542 30555 25594
rect 30579 25542 30609 25594
rect 30609 25542 30621 25594
rect 30621 25542 30635 25594
rect 30659 25542 30673 25594
rect 30673 25542 30685 25594
rect 30685 25542 30715 25594
rect 30739 25542 30749 25594
rect 30749 25542 30795 25594
rect 30499 25540 30555 25542
rect 30579 25540 30635 25542
rect 30659 25540 30715 25542
rect 30739 25540 30795 25542
rect 26278 25050 26334 25052
rect 26358 25050 26414 25052
rect 26438 25050 26494 25052
rect 26518 25050 26574 25052
rect 26278 24998 26324 25050
rect 26324 24998 26334 25050
rect 26358 24998 26388 25050
rect 26388 24998 26400 25050
rect 26400 24998 26414 25050
rect 26438 24998 26452 25050
rect 26452 24998 26464 25050
rect 26464 24998 26494 25050
rect 26518 24998 26528 25050
rect 26528 24998 26574 25050
rect 26278 24996 26334 24998
rect 26358 24996 26414 24998
rect 26438 24996 26494 24998
rect 26518 24996 26574 24998
rect 34719 25050 34775 25052
rect 34799 25050 34855 25052
rect 34879 25050 34935 25052
rect 34959 25050 35015 25052
rect 34719 24998 34765 25050
rect 34765 24998 34775 25050
rect 34799 24998 34829 25050
rect 34829 24998 34841 25050
rect 34841 24998 34855 25050
rect 34879 24998 34893 25050
rect 34893 24998 34905 25050
rect 34905 24998 34935 25050
rect 34959 24998 34969 25050
rect 34969 24998 35015 25050
rect 34719 24996 34775 24998
rect 34799 24996 34855 24998
rect 34879 24996 34935 24998
rect 34959 24996 35015 24998
rect 30499 24506 30555 24508
rect 30579 24506 30635 24508
rect 30659 24506 30715 24508
rect 30739 24506 30795 24508
rect 30499 24454 30545 24506
rect 30545 24454 30555 24506
rect 30579 24454 30609 24506
rect 30609 24454 30621 24506
rect 30621 24454 30635 24506
rect 30659 24454 30673 24506
rect 30673 24454 30685 24506
rect 30685 24454 30715 24506
rect 30739 24454 30749 24506
rect 30749 24454 30795 24506
rect 30499 24452 30555 24454
rect 30579 24452 30635 24454
rect 30659 24452 30715 24454
rect 30739 24452 30795 24454
rect 26278 23962 26334 23964
rect 26358 23962 26414 23964
rect 26438 23962 26494 23964
rect 26518 23962 26574 23964
rect 26278 23910 26324 23962
rect 26324 23910 26334 23962
rect 26358 23910 26388 23962
rect 26388 23910 26400 23962
rect 26400 23910 26414 23962
rect 26438 23910 26452 23962
rect 26452 23910 26464 23962
rect 26464 23910 26494 23962
rect 26518 23910 26528 23962
rect 26528 23910 26574 23962
rect 26278 23908 26334 23910
rect 26358 23908 26414 23910
rect 26438 23908 26494 23910
rect 26518 23908 26574 23910
rect 34719 23962 34775 23964
rect 34799 23962 34855 23964
rect 34879 23962 34935 23964
rect 34959 23962 35015 23964
rect 34719 23910 34765 23962
rect 34765 23910 34775 23962
rect 34799 23910 34829 23962
rect 34829 23910 34841 23962
rect 34841 23910 34855 23962
rect 34879 23910 34893 23962
rect 34893 23910 34905 23962
rect 34905 23910 34935 23962
rect 34959 23910 34969 23962
rect 34969 23910 35015 23962
rect 34719 23908 34775 23910
rect 34799 23908 34855 23910
rect 34879 23908 34935 23910
rect 34959 23908 35015 23910
rect 30499 23418 30555 23420
rect 30579 23418 30635 23420
rect 30659 23418 30715 23420
rect 30739 23418 30795 23420
rect 30499 23366 30545 23418
rect 30545 23366 30555 23418
rect 30579 23366 30609 23418
rect 30609 23366 30621 23418
rect 30621 23366 30635 23418
rect 30659 23366 30673 23418
rect 30673 23366 30685 23418
rect 30685 23366 30715 23418
rect 30739 23366 30749 23418
rect 30749 23366 30795 23418
rect 30499 23364 30555 23366
rect 30579 23364 30635 23366
rect 30659 23364 30715 23366
rect 30739 23364 30795 23366
rect 24490 23160 24546 23216
rect 26278 22874 26334 22876
rect 26358 22874 26414 22876
rect 26438 22874 26494 22876
rect 26518 22874 26574 22876
rect 26278 22822 26324 22874
rect 26324 22822 26334 22874
rect 26358 22822 26388 22874
rect 26388 22822 26400 22874
rect 26400 22822 26414 22874
rect 26438 22822 26452 22874
rect 26452 22822 26464 22874
rect 26464 22822 26494 22874
rect 26518 22822 26528 22874
rect 26528 22822 26574 22874
rect 26278 22820 26334 22822
rect 26358 22820 26414 22822
rect 26438 22820 26494 22822
rect 26518 22820 26574 22822
rect 34719 22874 34775 22876
rect 34799 22874 34855 22876
rect 34879 22874 34935 22876
rect 34959 22874 35015 22876
rect 34719 22822 34765 22874
rect 34765 22822 34775 22874
rect 34799 22822 34829 22874
rect 34829 22822 34841 22874
rect 34841 22822 34855 22874
rect 34879 22822 34893 22874
rect 34893 22822 34905 22874
rect 34905 22822 34935 22874
rect 34959 22822 34969 22874
rect 34969 22822 35015 22874
rect 34719 22820 34775 22822
rect 34799 22820 34855 22822
rect 34879 22820 34935 22822
rect 34959 22820 35015 22822
rect 30499 22330 30555 22332
rect 30579 22330 30635 22332
rect 30659 22330 30715 22332
rect 30739 22330 30795 22332
rect 30499 22278 30545 22330
rect 30545 22278 30555 22330
rect 30579 22278 30609 22330
rect 30609 22278 30621 22330
rect 30621 22278 30635 22330
rect 30659 22278 30673 22330
rect 30673 22278 30685 22330
rect 30685 22278 30715 22330
rect 30739 22278 30749 22330
rect 30749 22278 30795 22330
rect 30499 22276 30555 22278
rect 30579 22276 30635 22278
rect 30659 22276 30715 22278
rect 30739 22276 30795 22278
rect 26278 21786 26334 21788
rect 26358 21786 26414 21788
rect 26438 21786 26494 21788
rect 26518 21786 26574 21788
rect 26278 21734 26324 21786
rect 26324 21734 26334 21786
rect 26358 21734 26388 21786
rect 26388 21734 26400 21786
rect 26400 21734 26414 21786
rect 26438 21734 26452 21786
rect 26452 21734 26464 21786
rect 26464 21734 26494 21786
rect 26518 21734 26528 21786
rect 26528 21734 26574 21786
rect 26278 21732 26334 21734
rect 26358 21732 26414 21734
rect 26438 21732 26494 21734
rect 26518 21732 26574 21734
rect 34719 21786 34775 21788
rect 34799 21786 34855 21788
rect 34879 21786 34935 21788
rect 34959 21786 35015 21788
rect 34719 21734 34765 21786
rect 34765 21734 34775 21786
rect 34799 21734 34829 21786
rect 34829 21734 34841 21786
rect 34841 21734 34855 21786
rect 34879 21734 34893 21786
rect 34893 21734 34905 21786
rect 34905 21734 34935 21786
rect 34959 21734 34969 21786
rect 34969 21734 35015 21786
rect 34719 21732 34775 21734
rect 34799 21732 34855 21734
rect 34879 21732 34935 21734
rect 34959 21732 35015 21734
rect 30499 21242 30555 21244
rect 30579 21242 30635 21244
rect 30659 21242 30715 21244
rect 30739 21242 30795 21244
rect 30499 21190 30545 21242
rect 30545 21190 30555 21242
rect 30579 21190 30609 21242
rect 30609 21190 30621 21242
rect 30621 21190 30635 21242
rect 30659 21190 30673 21242
rect 30673 21190 30685 21242
rect 30685 21190 30715 21242
rect 30739 21190 30749 21242
rect 30749 21190 30795 21242
rect 30499 21188 30555 21190
rect 30579 21188 30635 21190
rect 30659 21188 30715 21190
rect 30739 21188 30795 21190
rect 26278 20698 26334 20700
rect 26358 20698 26414 20700
rect 26438 20698 26494 20700
rect 26518 20698 26574 20700
rect 26278 20646 26324 20698
rect 26324 20646 26334 20698
rect 26358 20646 26388 20698
rect 26388 20646 26400 20698
rect 26400 20646 26414 20698
rect 26438 20646 26452 20698
rect 26452 20646 26464 20698
rect 26464 20646 26494 20698
rect 26518 20646 26528 20698
rect 26528 20646 26574 20698
rect 26278 20644 26334 20646
rect 26358 20644 26414 20646
rect 26438 20644 26494 20646
rect 26518 20644 26574 20646
rect 34719 20698 34775 20700
rect 34799 20698 34855 20700
rect 34879 20698 34935 20700
rect 34959 20698 35015 20700
rect 34719 20646 34765 20698
rect 34765 20646 34775 20698
rect 34799 20646 34829 20698
rect 34829 20646 34841 20698
rect 34841 20646 34855 20698
rect 34879 20646 34893 20698
rect 34893 20646 34905 20698
rect 34905 20646 34935 20698
rect 34959 20646 34969 20698
rect 34969 20646 35015 20698
rect 34719 20644 34775 20646
rect 34799 20644 34855 20646
rect 34879 20644 34935 20646
rect 34959 20644 35015 20646
rect 30499 20154 30555 20156
rect 30579 20154 30635 20156
rect 30659 20154 30715 20156
rect 30739 20154 30795 20156
rect 30499 20102 30545 20154
rect 30545 20102 30555 20154
rect 30579 20102 30609 20154
rect 30609 20102 30621 20154
rect 30621 20102 30635 20154
rect 30659 20102 30673 20154
rect 30673 20102 30685 20154
rect 30685 20102 30715 20154
rect 30739 20102 30749 20154
rect 30749 20102 30795 20154
rect 30499 20100 30555 20102
rect 30579 20100 30635 20102
rect 30659 20100 30715 20102
rect 30739 20100 30795 20102
rect 34610 19780 34666 19816
rect 34610 19760 34612 19780
rect 34612 19760 34664 19780
rect 34664 19760 34666 19780
rect 26278 19610 26334 19612
rect 26358 19610 26414 19612
rect 26438 19610 26494 19612
rect 26518 19610 26574 19612
rect 26278 19558 26324 19610
rect 26324 19558 26334 19610
rect 26358 19558 26388 19610
rect 26388 19558 26400 19610
rect 26400 19558 26414 19610
rect 26438 19558 26452 19610
rect 26452 19558 26464 19610
rect 26464 19558 26494 19610
rect 26518 19558 26528 19610
rect 26528 19558 26574 19610
rect 26278 19556 26334 19558
rect 26358 19556 26414 19558
rect 26438 19556 26494 19558
rect 26518 19556 26574 19558
rect 34719 19610 34775 19612
rect 34799 19610 34855 19612
rect 34879 19610 34935 19612
rect 34959 19610 35015 19612
rect 34719 19558 34765 19610
rect 34765 19558 34775 19610
rect 34799 19558 34829 19610
rect 34829 19558 34841 19610
rect 34841 19558 34855 19610
rect 34879 19558 34893 19610
rect 34893 19558 34905 19610
rect 34905 19558 34935 19610
rect 34959 19558 34969 19610
rect 34969 19558 35015 19610
rect 34719 19556 34775 19558
rect 34799 19556 34855 19558
rect 34879 19556 34935 19558
rect 34959 19556 35015 19558
rect 30499 19066 30555 19068
rect 30579 19066 30635 19068
rect 30659 19066 30715 19068
rect 30739 19066 30795 19068
rect 30499 19014 30545 19066
rect 30545 19014 30555 19066
rect 30579 19014 30609 19066
rect 30609 19014 30621 19066
rect 30621 19014 30635 19066
rect 30659 19014 30673 19066
rect 30673 19014 30685 19066
rect 30685 19014 30715 19066
rect 30739 19014 30749 19066
rect 30749 19014 30795 19066
rect 30499 19012 30555 19014
rect 30579 19012 30635 19014
rect 30659 19012 30715 19014
rect 30739 19012 30795 19014
rect 26278 18522 26334 18524
rect 26358 18522 26414 18524
rect 26438 18522 26494 18524
rect 26518 18522 26574 18524
rect 26278 18470 26324 18522
rect 26324 18470 26334 18522
rect 26358 18470 26388 18522
rect 26388 18470 26400 18522
rect 26400 18470 26414 18522
rect 26438 18470 26452 18522
rect 26452 18470 26464 18522
rect 26464 18470 26494 18522
rect 26518 18470 26528 18522
rect 26528 18470 26574 18522
rect 26278 18468 26334 18470
rect 26358 18468 26414 18470
rect 26438 18468 26494 18470
rect 26518 18468 26574 18470
rect 34719 18522 34775 18524
rect 34799 18522 34855 18524
rect 34879 18522 34935 18524
rect 34959 18522 35015 18524
rect 34719 18470 34765 18522
rect 34765 18470 34775 18522
rect 34799 18470 34829 18522
rect 34829 18470 34841 18522
rect 34841 18470 34855 18522
rect 34879 18470 34893 18522
rect 34893 18470 34905 18522
rect 34905 18470 34935 18522
rect 34959 18470 34969 18522
rect 34969 18470 35015 18522
rect 34719 18468 34775 18470
rect 34799 18468 34855 18470
rect 34879 18468 34935 18470
rect 34959 18468 35015 18470
rect 30499 17978 30555 17980
rect 30579 17978 30635 17980
rect 30659 17978 30715 17980
rect 30739 17978 30795 17980
rect 30499 17926 30545 17978
rect 30545 17926 30555 17978
rect 30579 17926 30609 17978
rect 30609 17926 30621 17978
rect 30621 17926 30635 17978
rect 30659 17926 30673 17978
rect 30673 17926 30685 17978
rect 30685 17926 30715 17978
rect 30739 17926 30749 17978
rect 30749 17926 30795 17978
rect 30499 17924 30555 17926
rect 30579 17924 30635 17926
rect 30659 17924 30715 17926
rect 30739 17924 30795 17926
rect 26278 17434 26334 17436
rect 26358 17434 26414 17436
rect 26438 17434 26494 17436
rect 26518 17434 26574 17436
rect 26278 17382 26324 17434
rect 26324 17382 26334 17434
rect 26358 17382 26388 17434
rect 26388 17382 26400 17434
rect 26400 17382 26414 17434
rect 26438 17382 26452 17434
rect 26452 17382 26464 17434
rect 26464 17382 26494 17434
rect 26518 17382 26528 17434
rect 26528 17382 26574 17434
rect 26278 17380 26334 17382
rect 26358 17380 26414 17382
rect 26438 17380 26494 17382
rect 26518 17380 26574 17382
rect 34719 17434 34775 17436
rect 34799 17434 34855 17436
rect 34879 17434 34935 17436
rect 34959 17434 35015 17436
rect 34719 17382 34765 17434
rect 34765 17382 34775 17434
rect 34799 17382 34829 17434
rect 34829 17382 34841 17434
rect 34841 17382 34855 17434
rect 34879 17382 34893 17434
rect 34893 17382 34905 17434
rect 34905 17382 34935 17434
rect 34959 17382 34969 17434
rect 34969 17382 35015 17434
rect 34719 17380 34775 17382
rect 34799 17380 34855 17382
rect 34879 17380 34935 17382
rect 34959 17380 35015 17382
rect 30499 16890 30555 16892
rect 30579 16890 30635 16892
rect 30659 16890 30715 16892
rect 30739 16890 30795 16892
rect 30499 16838 30545 16890
rect 30545 16838 30555 16890
rect 30579 16838 30609 16890
rect 30609 16838 30621 16890
rect 30621 16838 30635 16890
rect 30659 16838 30673 16890
rect 30673 16838 30685 16890
rect 30685 16838 30715 16890
rect 30739 16838 30749 16890
rect 30749 16838 30795 16890
rect 30499 16836 30555 16838
rect 30579 16836 30635 16838
rect 30659 16836 30715 16838
rect 30739 16836 30795 16838
rect 26278 16346 26334 16348
rect 26358 16346 26414 16348
rect 26438 16346 26494 16348
rect 26518 16346 26574 16348
rect 26278 16294 26324 16346
rect 26324 16294 26334 16346
rect 26358 16294 26388 16346
rect 26388 16294 26400 16346
rect 26400 16294 26414 16346
rect 26438 16294 26452 16346
rect 26452 16294 26464 16346
rect 26464 16294 26494 16346
rect 26518 16294 26528 16346
rect 26528 16294 26574 16346
rect 26278 16292 26334 16294
rect 26358 16292 26414 16294
rect 26438 16292 26494 16294
rect 26518 16292 26574 16294
rect 34719 16346 34775 16348
rect 34799 16346 34855 16348
rect 34879 16346 34935 16348
rect 34959 16346 35015 16348
rect 34719 16294 34765 16346
rect 34765 16294 34775 16346
rect 34799 16294 34829 16346
rect 34829 16294 34841 16346
rect 34841 16294 34855 16346
rect 34879 16294 34893 16346
rect 34893 16294 34905 16346
rect 34905 16294 34935 16346
rect 34959 16294 34969 16346
rect 34969 16294 35015 16346
rect 34719 16292 34775 16294
rect 34799 16292 34855 16294
rect 34879 16292 34935 16294
rect 34959 16292 35015 16294
rect 30499 15802 30555 15804
rect 30579 15802 30635 15804
rect 30659 15802 30715 15804
rect 30739 15802 30795 15804
rect 30499 15750 30545 15802
rect 30545 15750 30555 15802
rect 30579 15750 30609 15802
rect 30609 15750 30621 15802
rect 30621 15750 30635 15802
rect 30659 15750 30673 15802
rect 30673 15750 30685 15802
rect 30685 15750 30715 15802
rect 30739 15750 30749 15802
rect 30749 15750 30795 15802
rect 30499 15748 30555 15750
rect 30579 15748 30635 15750
rect 30659 15748 30715 15750
rect 30739 15748 30795 15750
rect 26278 15258 26334 15260
rect 26358 15258 26414 15260
rect 26438 15258 26494 15260
rect 26518 15258 26574 15260
rect 26278 15206 26324 15258
rect 26324 15206 26334 15258
rect 26358 15206 26388 15258
rect 26388 15206 26400 15258
rect 26400 15206 26414 15258
rect 26438 15206 26452 15258
rect 26452 15206 26464 15258
rect 26464 15206 26494 15258
rect 26518 15206 26528 15258
rect 26528 15206 26574 15258
rect 26278 15204 26334 15206
rect 26358 15204 26414 15206
rect 26438 15204 26494 15206
rect 26518 15204 26574 15206
rect 34719 15258 34775 15260
rect 34799 15258 34855 15260
rect 34879 15258 34935 15260
rect 34959 15258 35015 15260
rect 34719 15206 34765 15258
rect 34765 15206 34775 15258
rect 34799 15206 34829 15258
rect 34829 15206 34841 15258
rect 34841 15206 34855 15258
rect 34879 15206 34893 15258
rect 34893 15206 34905 15258
rect 34905 15206 34935 15258
rect 34959 15206 34969 15258
rect 34969 15206 35015 15258
rect 34719 15204 34775 15206
rect 34799 15204 34855 15206
rect 34879 15204 34935 15206
rect 34959 15204 35015 15206
rect 30499 14714 30555 14716
rect 30579 14714 30635 14716
rect 30659 14714 30715 14716
rect 30739 14714 30795 14716
rect 30499 14662 30545 14714
rect 30545 14662 30555 14714
rect 30579 14662 30609 14714
rect 30609 14662 30621 14714
rect 30621 14662 30635 14714
rect 30659 14662 30673 14714
rect 30673 14662 30685 14714
rect 30685 14662 30715 14714
rect 30739 14662 30749 14714
rect 30749 14662 30795 14714
rect 30499 14660 30555 14662
rect 30579 14660 30635 14662
rect 30659 14660 30715 14662
rect 30739 14660 30795 14662
rect 26278 14170 26334 14172
rect 26358 14170 26414 14172
rect 26438 14170 26494 14172
rect 26518 14170 26574 14172
rect 26278 14118 26324 14170
rect 26324 14118 26334 14170
rect 26358 14118 26388 14170
rect 26388 14118 26400 14170
rect 26400 14118 26414 14170
rect 26438 14118 26452 14170
rect 26452 14118 26464 14170
rect 26464 14118 26494 14170
rect 26518 14118 26528 14170
rect 26528 14118 26574 14170
rect 26278 14116 26334 14118
rect 26358 14116 26414 14118
rect 26438 14116 26494 14118
rect 26518 14116 26574 14118
rect 34719 14170 34775 14172
rect 34799 14170 34855 14172
rect 34879 14170 34935 14172
rect 34959 14170 35015 14172
rect 34719 14118 34765 14170
rect 34765 14118 34775 14170
rect 34799 14118 34829 14170
rect 34829 14118 34841 14170
rect 34841 14118 34855 14170
rect 34879 14118 34893 14170
rect 34893 14118 34905 14170
rect 34905 14118 34935 14170
rect 34959 14118 34969 14170
rect 34969 14118 35015 14170
rect 34719 14116 34775 14118
rect 34799 14116 34855 14118
rect 34879 14116 34935 14118
rect 34959 14116 35015 14118
rect 30499 13626 30555 13628
rect 30579 13626 30635 13628
rect 30659 13626 30715 13628
rect 30739 13626 30795 13628
rect 30499 13574 30545 13626
rect 30545 13574 30555 13626
rect 30579 13574 30609 13626
rect 30609 13574 30621 13626
rect 30621 13574 30635 13626
rect 30659 13574 30673 13626
rect 30673 13574 30685 13626
rect 30685 13574 30715 13626
rect 30739 13574 30749 13626
rect 30749 13574 30795 13626
rect 30499 13572 30555 13574
rect 30579 13572 30635 13574
rect 30659 13572 30715 13574
rect 30739 13572 30795 13574
rect 26278 13082 26334 13084
rect 26358 13082 26414 13084
rect 26438 13082 26494 13084
rect 26518 13082 26574 13084
rect 26278 13030 26324 13082
rect 26324 13030 26334 13082
rect 26358 13030 26388 13082
rect 26388 13030 26400 13082
rect 26400 13030 26414 13082
rect 26438 13030 26452 13082
rect 26452 13030 26464 13082
rect 26464 13030 26494 13082
rect 26518 13030 26528 13082
rect 26528 13030 26574 13082
rect 26278 13028 26334 13030
rect 26358 13028 26414 13030
rect 26438 13028 26494 13030
rect 26518 13028 26574 13030
rect 34719 13082 34775 13084
rect 34799 13082 34855 13084
rect 34879 13082 34935 13084
rect 34959 13082 35015 13084
rect 34719 13030 34765 13082
rect 34765 13030 34775 13082
rect 34799 13030 34829 13082
rect 34829 13030 34841 13082
rect 34841 13030 34855 13082
rect 34879 13030 34893 13082
rect 34893 13030 34905 13082
rect 34905 13030 34935 13082
rect 34959 13030 34969 13082
rect 34969 13030 35015 13082
rect 34719 13028 34775 13030
rect 34799 13028 34855 13030
rect 34879 13028 34935 13030
rect 34959 13028 35015 13030
rect 35162 12960 35218 13016
rect 22058 12538 22114 12540
rect 22138 12538 22194 12540
rect 22218 12538 22274 12540
rect 22298 12538 22354 12540
rect 22058 12486 22104 12538
rect 22104 12486 22114 12538
rect 22138 12486 22168 12538
rect 22168 12486 22180 12538
rect 22180 12486 22194 12538
rect 22218 12486 22232 12538
rect 22232 12486 22244 12538
rect 22244 12486 22274 12538
rect 22298 12486 22308 12538
rect 22308 12486 22354 12538
rect 22058 12484 22114 12486
rect 22138 12484 22194 12486
rect 22218 12484 22274 12486
rect 22298 12484 22354 12486
rect 30499 12538 30555 12540
rect 30579 12538 30635 12540
rect 30659 12538 30715 12540
rect 30739 12538 30795 12540
rect 30499 12486 30545 12538
rect 30545 12486 30555 12538
rect 30579 12486 30609 12538
rect 30609 12486 30621 12538
rect 30621 12486 30635 12538
rect 30659 12486 30673 12538
rect 30673 12486 30685 12538
rect 30685 12486 30715 12538
rect 30739 12486 30749 12538
rect 30749 12486 30795 12538
rect 30499 12484 30555 12486
rect 30579 12484 30635 12486
rect 30659 12484 30715 12486
rect 30739 12484 30795 12486
rect 9396 11994 9452 11996
rect 9476 11994 9532 11996
rect 9556 11994 9612 11996
rect 9636 11994 9692 11996
rect 9396 11942 9442 11994
rect 9442 11942 9452 11994
rect 9476 11942 9506 11994
rect 9506 11942 9518 11994
rect 9518 11942 9532 11994
rect 9556 11942 9570 11994
rect 9570 11942 9582 11994
rect 9582 11942 9612 11994
rect 9636 11942 9646 11994
rect 9646 11942 9692 11994
rect 9396 11940 9452 11942
rect 9476 11940 9532 11942
rect 9556 11940 9612 11942
rect 9636 11940 9692 11942
rect 17837 11994 17893 11996
rect 17917 11994 17973 11996
rect 17997 11994 18053 11996
rect 18077 11994 18133 11996
rect 17837 11942 17883 11994
rect 17883 11942 17893 11994
rect 17917 11942 17947 11994
rect 17947 11942 17959 11994
rect 17959 11942 17973 11994
rect 17997 11942 18011 11994
rect 18011 11942 18023 11994
rect 18023 11942 18053 11994
rect 18077 11942 18087 11994
rect 18087 11942 18133 11994
rect 17837 11940 17893 11942
rect 17917 11940 17973 11942
rect 17997 11940 18053 11942
rect 18077 11940 18133 11942
rect 5176 11450 5232 11452
rect 5256 11450 5312 11452
rect 5336 11450 5392 11452
rect 5416 11450 5472 11452
rect 5176 11398 5222 11450
rect 5222 11398 5232 11450
rect 5256 11398 5286 11450
rect 5286 11398 5298 11450
rect 5298 11398 5312 11450
rect 5336 11398 5350 11450
rect 5350 11398 5362 11450
rect 5362 11398 5392 11450
rect 5416 11398 5426 11450
rect 5426 11398 5472 11450
rect 5176 11396 5232 11398
rect 5256 11396 5312 11398
rect 5336 11396 5392 11398
rect 5416 11396 5472 11398
rect 13617 11450 13673 11452
rect 13697 11450 13753 11452
rect 13777 11450 13833 11452
rect 13857 11450 13913 11452
rect 13617 11398 13663 11450
rect 13663 11398 13673 11450
rect 13697 11398 13727 11450
rect 13727 11398 13739 11450
rect 13739 11398 13753 11450
rect 13777 11398 13791 11450
rect 13791 11398 13803 11450
rect 13803 11398 13833 11450
rect 13857 11398 13867 11450
rect 13867 11398 13913 11450
rect 13617 11396 13673 11398
rect 13697 11396 13753 11398
rect 13777 11396 13833 11398
rect 13857 11396 13913 11398
rect 9396 10906 9452 10908
rect 9476 10906 9532 10908
rect 9556 10906 9612 10908
rect 9636 10906 9692 10908
rect 9396 10854 9442 10906
rect 9442 10854 9452 10906
rect 9476 10854 9506 10906
rect 9506 10854 9518 10906
rect 9518 10854 9532 10906
rect 9556 10854 9570 10906
rect 9570 10854 9582 10906
rect 9582 10854 9612 10906
rect 9636 10854 9646 10906
rect 9646 10854 9692 10906
rect 9396 10852 9452 10854
rect 9476 10852 9532 10854
rect 9556 10852 9612 10854
rect 9636 10852 9692 10854
rect 17837 10906 17893 10908
rect 17917 10906 17973 10908
rect 17997 10906 18053 10908
rect 18077 10906 18133 10908
rect 17837 10854 17883 10906
rect 17883 10854 17893 10906
rect 17917 10854 17947 10906
rect 17947 10854 17959 10906
rect 17959 10854 17973 10906
rect 17997 10854 18011 10906
rect 18011 10854 18023 10906
rect 18023 10854 18053 10906
rect 18077 10854 18087 10906
rect 18087 10854 18133 10906
rect 17837 10852 17893 10854
rect 17917 10852 17973 10854
rect 17997 10852 18053 10854
rect 18077 10852 18133 10854
rect 5176 10362 5232 10364
rect 5256 10362 5312 10364
rect 5336 10362 5392 10364
rect 5416 10362 5472 10364
rect 5176 10310 5222 10362
rect 5222 10310 5232 10362
rect 5256 10310 5286 10362
rect 5286 10310 5298 10362
rect 5298 10310 5312 10362
rect 5336 10310 5350 10362
rect 5350 10310 5362 10362
rect 5362 10310 5392 10362
rect 5416 10310 5426 10362
rect 5426 10310 5472 10362
rect 5176 10308 5232 10310
rect 5256 10308 5312 10310
rect 5336 10308 5392 10310
rect 5416 10308 5472 10310
rect 13617 10362 13673 10364
rect 13697 10362 13753 10364
rect 13777 10362 13833 10364
rect 13857 10362 13913 10364
rect 13617 10310 13663 10362
rect 13663 10310 13673 10362
rect 13697 10310 13727 10362
rect 13727 10310 13739 10362
rect 13739 10310 13753 10362
rect 13777 10310 13791 10362
rect 13791 10310 13803 10362
rect 13803 10310 13833 10362
rect 13857 10310 13867 10362
rect 13867 10310 13913 10362
rect 13617 10308 13673 10310
rect 13697 10308 13753 10310
rect 13777 10308 13833 10310
rect 13857 10308 13913 10310
rect 9396 9818 9452 9820
rect 9476 9818 9532 9820
rect 9556 9818 9612 9820
rect 9636 9818 9692 9820
rect 9396 9766 9442 9818
rect 9442 9766 9452 9818
rect 9476 9766 9506 9818
rect 9506 9766 9518 9818
rect 9518 9766 9532 9818
rect 9556 9766 9570 9818
rect 9570 9766 9582 9818
rect 9582 9766 9612 9818
rect 9636 9766 9646 9818
rect 9646 9766 9692 9818
rect 9396 9764 9452 9766
rect 9476 9764 9532 9766
rect 9556 9764 9612 9766
rect 9636 9764 9692 9766
rect 17837 9818 17893 9820
rect 17917 9818 17973 9820
rect 17997 9818 18053 9820
rect 18077 9818 18133 9820
rect 17837 9766 17883 9818
rect 17883 9766 17893 9818
rect 17917 9766 17947 9818
rect 17947 9766 17959 9818
rect 17959 9766 17973 9818
rect 17997 9766 18011 9818
rect 18011 9766 18023 9818
rect 18023 9766 18053 9818
rect 18077 9766 18087 9818
rect 18087 9766 18133 9818
rect 17837 9764 17893 9766
rect 17917 9764 17973 9766
rect 17997 9764 18053 9766
rect 18077 9764 18133 9766
rect 5176 9274 5232 9276
rect 5256 9274 5312 9276
rect 5336 9274 5392 9276
rect 5416 9274 5472 9276
rect 5176 9222 5222 9274
rect 5222 9222 5232 9274
rect 5256 9222 5286 9274
rect 5286 9222 5298 9274
rect 5298 9222 5312 9274
rect 5336 9222 5350 9274
rect 5350 9222 5362 9274
rect 5362 9222 5392 9274
rect 5416 9222 5426 9274
rect 5426 9222 5472 9274
rect 5176 9220 5232 9222
rect 5256 9220 5312 9222
rect 5336 9220 5392 9222
rect 5416 9220 5472 9222
rect 13617 9274 13673 9276
rect 13697 9274 13753 9276
rect 13777 9274 13833 9276
rect 13857 9274 13913 9276
rect 13617 9222 13663 9274
rect 13663 9222 13673 9274
rect 13697 9222 13727 9274
rect 13727 9222 13739 9274
rect 13739 9222 13753 9274
rect 13777 9222 13791 9274
rect 13791 9222 13803 9274
rect 13803 9222 13833 9274
rect 13857 9222 13867 9274
rect 13867 9222 13913 9274
rect 13617 9220 13673 9222
rect 13697 9220 13753 9222
rect 13777 9220 13833 9222
rect 13857 9220 13913 9222
rect 9396 8730 9452 8732
rect 9476 8730 9532 8732
rect 9556 8730 9612 8732
rect 9636 8730 9692 8732
rect 9396 8678 9442 8730
rect 9442 8678 9452 8730
rect 9476 8678 9506 8730
rect 9506 8678 9518 8730
rect 9518 8678 9532 8730
rect 9556 8678 9570 8730
rect 9570 8678 9582 8730
rect 9582 8678 9612 8730
rect 9636 8678 9646 8730
rect 9646 8678 9692 8730
rect 9396 8676 9452 8678
rect 9476 8676 9532 8678
rect 9556 8676 9612 8678
rect 9636 8676 9692 8678
rect 17837 8730 17893 8732
rect 17917 8730 17973 8732
rect 17997 8730 18053 8732
rect 18077 8730 18133 8732
rect 17837 8678 17883 8730
rect 17883 8678 17893 8730
rect 17917 8678 17947 8730
rect 17947 8678 17959 8730
rect 17959 8678 17973 8730
rect 17997 8678 18011 8730
rect 18011 8678 18023 8730
rect 18023 8678 18053 8730
rect 18077 8678 18087 8730
rect 18087 8678 18133 8730
rect 17837 8676 17893 8678
rect 17917 8676 17973 8678
rect 17997 8676 18053 8678
rect 18077 8676 18133 8678
rect 5176 8186 5232 8188
rect 5256 8186 5312 8188
rect 5336 8186 5392 8188
rect 5416 8186 5472 8188
rect 5176 8134 5222 8186
rect 5222 8134 5232 8186
rect 5256 8134 5286 8186
rect 5286 8134 5298 8186
rect 5298 8134 5312 8186
rect 5336 8134 5350 8186
rect 5350 8134 5362 8186
rect 5362 8134 5392 8186
rect 5416 8134 5426 8186
rect 5426 8134 5472 8186
rect 5176 8132 5232 8134
rect 5256 8132 5312 8134
rect 5336 8132 5392 8134
rect 5416 8132 5472 8134
rect 13617 8186 13673 8188
rect 13697 8186 13753 8188
rect 13777 8186 13833 8188
rect 13857 8186 13913 8188
rect 13617 8134 13663 8186
rect 13663 8134 13673 8186
rect 13697 8134 13727 8186
rect 13727 8134 13739 8186
rect 13739 8134 13753 8186
rect 13777 8134 13791 8186
rect 13791 8134 13803 8186
rect 13803 8134 13833 8186
rect 13857 8134 13867 8186
rect 13867 8134 13913 8186
rect 13617 8132 13673 8134
rect 13697 8132 13753 8134
rect 13777 8132 13833 8134
rect 13857 8132 13913 8134
rect 9396 7642 9452 7644
rect 9476 7642 9532 7644
rect 9556 7642 9612 7644
rect 9636 7642 9692 7644
rect 9396 7590 9442 7642
rect 9442 7590 9452 7642
rect 9476 7590 9506 7642
rect 9506 7590 9518 7642
rect 9518 7590 9532 7642
rect 9556 7590 9570 7642
rect 9570 7590 9582 7642
rect 9582 7590 9612 7642
rect 9636 7590 9646 7642
rect 9646 7590 9692 7642
rect 9396 7588 9452 7590
rect 9476 7588 9532 7590
rect 9556 7588 9612 7590
rect 9636 7588 9692 7590
rect 17837 7642 17893 7644
rect 17917 7642 17973 7644
rect 17997 7642 18053 7644
rect 18077 7642 18133 7644
rect 17837 7590 17883 7642
rect 17883 7590 17893 7642
rect 17917 7590 17947 7642
rect 17947 7590 17959 7642
rect 17959 7590 17973 7642
rect 17997 7590 18011 7642
rect 18011 7590 18023 7642
rect 18023 7590 18053 7642
rect 18077 7590 18087 7642
rect 18087 7590 18133 7642
rect 17837 7588 17893 7590
rect 17917 7588 17973 7590
rect 17997 7588 18053 7590
rect 18077 7588 18133 7590
rect 5176 7098 5232 7100
rect 5256 7098 5312 7100
rect 5336 7098 5392 7100
rect 5416 7098 5472 7100
rect 5176 7046 5222 7098
rect 5222 7046 5232 7098
rect 5256 7046 5286 7098
rect 5286 7046 5298 7098
rect 5298 7046 5312 7098
rect 5336 7046 5350 7098
rect 5350 7046 5362 7098
rect 5362 7046 5392 7098
rect 5416 7046 5426 7098
rect 5426 7046 5472 7098
rect 5176 7044 5232 7046
rect 5256 7044 5312 7046
rect 5336 7044 5392 7046
rect 5416 7044 5472 7046
rect 13617 7098 13673 7100
rect 13697 7098 13753 7100
rect 13777 7098 13833 7100
rect 13857 7098 13913 7100
rect 13617 7046 13663 7098
rect 13663 7046 13673 7098
rect 13697 7046 13727 7098
rect 13727 7046 13739 7098
rect 13739 7046 13753 7098
rect 13777 7046 13791 7098
rect 13791 7046 13803 7098
rect 13803 7046 13833 7098
rect 13857 7046 13867 7098
rect 13867 7046 13913 7098
rect 13617 7044 13673 7046
rect 13697 7044 13753 7046
rect 13777 7044 13833 7046
rect 13857 7044 13913 7046
rect 1398 6840 1454 6896
rect 9396 6554 9452 6556
rect 9476 6554 9532 6556
rect 9556 6554 9612 6556
rect 9636 6554 9692 6556
rect 9396 6502 9442 6554
rect 9442 6502 9452 6554
rect 9476 6502 9506 6554
rect 9506 6502 9518 6554
rect 9518 6502 9532 6554
rect 9556 6502 9570 6554
rect 9570 6502 9582 6554
rect 9582 6502 9612 6554
rect 9636 6502 9646 6554
rect 9646 6502 9692 6554
rect 9396 6500 9452 6502
rect 9476 6500 9532 6502
rect 9556 6500 9612 6502
rect 9636 6500 9692 6502
rect 17837 6554 17893 6556
rect 17917 6554 17973 6556
rect 17997 6554 18053 6556
rect 18077 6554 18133 6556
rect 17837 6502 17883 6554
rect 17883 6502 17893 6554
rect 17917 6502 17947 6554
rect 17947 6502 17959 6554
rect 17959 6502 17973 6554
rect 17997 6502 18011 6554
rect 18011 6502 18023 6554
rect 18023 6502 18053 6554
rect 18077 6502 18087 6554
rect 18087 6502 18133 6554
rect 17837 6500 17893 6502
rect 17917 6500 17973 6502
rect 17997 6500 18053 6502
rect 18077 6500 18133 6502
rect 5176 6010 5232 6012
rect 5256 6010 5312 6012
rect 5336 6010 5392 6012
rect 5416 6010 5472 6012
rect 5176 5958 5222 6010
rect 5222 5958 5232 6010
rect 5256 5958 5286 6010
rect 5286 5958 5298 6010
rect 5298 5958 5312 6010
rect 5336 5958 5350 6010
rect 5350 5958 5362 6010
rect 5362 5958 5392 6010
rect 5416 5958 5426 6010
rect 5426 5958 5472 6010
rect 5176 5956 5232 5958
rect 5256 5956 5312 5958
rect 5336 5956 5392 5958
rect 5416 5956 5472 5958
rect 13617 6010 13673 6012
rect 13697 6010 13753 6012
rect 13777 6010 13833 6012
rect 13857 6010 13913 6012
rect 13617 5958 13663 6010
rect 13663 5958 13673 6010
rect 13697 5958 13727 6010
rect 13727 5958 13739 6010
rect 13739 5958 13753 6010
rect 13777 5958 13791 6010
rect 13791 5958 13803 6010
rect 13803 5958 13833 6010
rect 13857 5958 13867 6010
rect 13867 5958 13913 6010
rect 13617 5956 13673 5958
rect 13697 5956 13753 5958
rect 13777 5956 13833 5958
rect 13857 5956 13913 5958
rect 9396 5466 9452 5468
rect 9476 5466 9532 5468
rect 9556 5466 9612 5468
rect 9636 5466 9692 5468
rect 9396 5414 9442 5466
rect 9442 5414 9452 5466
rect 9476 5414 9506 5466
rect 9506 5414 9518 5466
rect 9518 5414 9532 5466
rect 9556 5414 9570 5466
rect 9570 5414 9582 5466
rect 9582 5414 9612 5466
rect 9636 5414 9646 5466
rect 9646 5414 9692 5466
rect 9396 5412 9452 5414
rect 9476 5412 9532 5414
rect 9556 5412 9612 5414
rect 9636 5412 9692 5414
rect 17837 5466 17893 5468
rect 17917 5466 17973 5468
rect 17997 5466 18053 5468
rect 18077 5466 18133 5468
rect 17837 5414 17883 5466
rect 17883 5414 17893 5466
rect 17917 5414 17947 5466
rect 17947 5414 17959 5466
rect 17959 5414 17973 5466
rect 17997 5414 18011 5466
rect 18011 5414 18023 5466
rect 18023 5414 18053 5466
rect 18077 5414 18087 5466
rect 18087 5414 18133 5466
rect 17837 5412 17893 5414
rect 17917 5412 17973 5414
rect 17997 5412 18053 5414
rect 18077 5412 18133 5414
rect 5176 4922 5232 4924
rect 5256 4922 5312 4924
rect 5336 4922 5392 4924
rect 5416 4922 5472 4924
rect 5176 4870 5222 4922
rect 5222 4870 5232 4922
rect 5256 4870 5286 4922
rect 5286 4870 5298 4922
rect 5298 4870 5312 4922
rect 5336 4870 5350 4922
rect 5350 4870 5362 4922
rect 5362 4870 5392 4922
rect 5416 4870 5426 4922
rect 5426 4870 5472 4922
rect 5176 4868 5232 4870
rect 5256 4868 5312 4870
rect 5336 4868 5392 4870
rect 5416 4868 5472 4870
rect 13617 4922 13673 4924
rect 13697 4922 13753 4924
rect 13777 4922 13833 4924
rect 13857 4922 13913 4924
rect 13617 4870 13663 4922
rect 13663 4870 13673 4922
rect 13697 4870 13727 4922
rect 13727 4870 13739 4922
rect 13739 4870 13753 4922
rect 13777 4870 13791 4922
rect 13791 4870 13803 4922
rect 13803 4870 13833 4922
rect 13857 4870 13867 4922
rect 13867 4870 13913 4922
rect 13617 4868 13673 4870
rect 13697 4868 13753 4870
rect 13777 4868 13833 4870
rect 13857 4868 13913 4870
rect 9396 4378 9452 4380
rect 9476 4378 9532 4380
rect 9556 4378 9612 4380
rect 9636 4378 9692 4380
rect 9396 4326 9442 4378
rect 9442 4326 9452 4378
rect 9476 4326 9506 4378
rect 9506 4326 9518 4378
rect 9518 4326 9532 4378
rect 9556 4326 9570 4378
rect 9570 4326 9582 4378
rect 9582 4326 9612 4378
rect 9636 4326 9646 4378
rect 9646 4326 9692 4378
rect 9396 4324 9452 4326
rect 9476 4324 9532 4326
rect 9556 4324 9612 4326
rect 9636 4324 9692 4326
rect 17837 4378 17893 4380
rect 17917 4378 17973 4380
rect 17997 4378 18053 4380
rect 18077 4378 18133 4380
rect 17837 4326 17883 4378
rect 17883 4326 17893 4378
rect 17917 4326 17947 4378
rect 17947 4326 17959 4378
rect 17959 4326 17973 4378
rect 17997 4326 18011 4378
rect 18011 4326 18023 4378
rect 18023 4326 18053 4378
rect 18077 4326 18087 4378
rect 18087 4326 18133 4378
rect 17837 4324 17893 4326
rect 17917 4324 17973 4326
rect 17997 4324 18053 4326
rect 18077 4324 18133 4326
rect 5176 3834 5232 3836
rect 5256 3834 5312 3836
rect 5336 3834 5392 3836
rect 5416 3834 5472 3836
rect 5176 3782 5222 3834
rect 5222 3782 5232 3834
rect 5256 3782 5286 3834
rect 5286 3782 5298 3834
rect 5298 3782 5312 3834
rect 5336 3782 5350 3834
rect 5350 3782 5362 3834
rect 5362 3782 5392 3834
rect 5416 3782 5426 3834
rect 5426 3782 5472 3834
rect 5176 3780 5232 3782
rect 5256 3780 5312 3782
rect 5336 3780 5392 3782
rect 5416 3780 5472 3782
rect 13617 3834 13673 3836
rect 13697 3834 13753 3836
rect 13777 3834 13833 3836
rect 13857 3834 13913 3836
rect 13617 3782 13663 3834
rect 13663 3782 13673 3834
rect 13697 3782 13727 3834
rect 13727 3782 13739 3834
rect 13739 3782 13753 3834
rect 13777 3782 13791 3834
rect 13791 3782 13803 3834
rect 13803 3782 13833 3834
rect 13857 3782 13867 3834
rect 13867 3782 13913 3834
rect 13617 3780 13673 3782
rect 13697 3780 13753 3782
rect 13777 3780 13833 3782
rect 13857 3780 13913 3782
rect 9396 3290 9452 3292
rect 9476 3290 9532 3292
rect 9556 3290 9612 3292
rect 9636 3290 9692 3292
rect 9396 3238 9442 3290
rect 9442 3238 9452 3290
rect 9476 3238 9506 3290
rect 9506 3238 9518 3290
rect 9518 3238 9532 3290
rect 9556 3238 9570 3290
rect 9570 3238 9582 3290
rect 9582 3238 9612 3290
rect 9636 3238 9646 3290
rect 9646 3238 9692 3290
rect 9396 3236 9452 3238
rect 9476 3236 9532 3238
rect 9556 3236 9612 3238
rect 9636 3236 9692 3238
rect 17837 3290 17893 3292
rect 17917 3290 17973 3292
rect 17997 3290 18053 3292
rect 18077 3290 18133 3292
rect 17837 3238 17883 3290
rect 17883 3238 17893 3290
rect 17917 3238 17947 3290
rect 17947 3238 17959 3290
rect 17959 3238 17973 3290
rect 17997 3238 18011 3290
rect 18011 3238 18023 3290
rect 18023 3238 18053 3290
rect 18077 3238 18087 3290
rect 18087 3238 18133 3290
rect 17837 3236 17893 3238
rect 17917 3236 17973 3238
rect 17997 3236 18053 3238
rect 18077 3236 18133 3238
rect 5176 2746 5232 2748
rect 5256 2746 5312 2748
rect 5336 2746 5392 2748
rect 5416 2746 5472 2748
rect 5176 2694 5222 2746
rect 5222 2694 5232 2746
rect 5256 2694 5286 2746
rect 5286 2694 5298 2746
rect 5298 2694 5312 2746
rect 5336 2694 5350 2746
rect 5350 2694 5362 2746
rect 5362 2694 5392 2746
rect 5416 2694 5426 2746
rect 5426 2694 5472 2746
rect 5176 2692 5232 2694
rect 5256 2692 5312 2694
rect 5336 2692 5392 2694
rect 5416 2692 5472 2694
rect 13617 2746 13673 2748
rect 13697 2746 13753 2748
rect 13777 2746 13833 2748
rect 13857 2746 13913 2748
rect 13617 2694 13663 2746
rect 13663 2694 13673 2746
rect 13697 2694 13727 2746
rect 13727 2694 13739 2746
rect 13739 2694 13753 2746
rect 13777 2694 13791 2746
rect 13791 2694 13803 2746
rect 13803 2694 13833 2746
rect 13857 2694 13867 2746
rect 13867 2694 13913 2746
rect 13617 2692 13673 2694
rect 13697 2692 13753 2694
rect 13777 2692 13833 2694
rect 13857 2692 13913 2694
rect 26278 11994 26334 11996
rect 26358 11994 26414 11996
rect 26438 11994 26494 11996
rect 26518 11994 26574 11996
rect 26278 11942 26324 11994
rect 26324 11942 26334 11994
rect 26358 11942 26388 11994
rect 26388 11942 26400 11994
rect 26400 11942 26414 11994
rect 26438 11942 26452 11994
rect 26452 11942 26464 11994
rect 26464 11942 26494 11994
rect 26518 11942 26528 11994
rect 26528 11942 26574 11994
rect 26278 11940 26334 11942
rect 26358 11940 26414 11942
rect 26438 11940 26494 11942
rect 26518 11940 26574 11942
rect 34719 11994 34775 11996
rect 34799 11994 34855 11996
rect 34879 11994 34935 11996
rect 34959 11994 35015 11996
rect 34719 11942 34765 11994
rect 34765 11942 34775 11994
rect 34799 11942 34829 11994
rect 34829 11942 34841 11994
rect 34841 11942 34855 11994
rect 34879 11942 34893 11994
rect 34893 11942 34905 11994
rect 34905 11942 34935 11994
rect 34959 11942 34969 11994
rect 34969 11942 35015 11994
rect 34719 11940 34775 11942
rect 34799 11940 34855 11942
rect 34879 11940 34935 11942
rect 34959 11940 35015 11942
rect 22058 11450 22114 11452
rect 22138 11450 22194 11452
rect 22218 11450 22274 11452
rect 22298 11450 22354 11452
rect 22058 11398 22104 11450
rect 22104 11398 22114 11450
rect 22138 11398 22168 11450
rect 22168 11398 22180 11450
rect 22180 11398 22194 11450
rect 22218 11398 22232 11450
rect 22232 11398 22244 11450
rect 22244 11398 22274 11450
rect 22298 11398 22308 11450
rect 22308 11398 22354 11450
rect 22058 11396 22114 11398
rect 22138 11396 22194 11398
rect 22218 11396 22274 11398
rect 22298 11396 22354 11398
rect 30499 11450 30555 11452
rect 30579 11450 30635 11452
rect 30659 11450 30715 11452
rect 30739 11450 30795 11452
rect 30499 11398 30545 11450
rect 30545 11398 30555 11450
rect 30579 11398 30609 11450
rect 30609 11398 30621 11450
rect 30621 11398 30635 11450
rect 30659 11398 30673 11450
rect 30673 11398 30685 11450
rect 30685 11398 30715 11450
rect 30739 11398 30749 11450
rect 30749 11398 30795 11450
rect 30499 11396 30555 11398
rect 30579 11396 30635 11398
rect 30659 11396 30715 11398
rect 30739 11396 30795 11398
rect 26278 10906 26334 10908
rect 26358 10906 26414 10908
rect 26438 10906 26494 10908
rect 26518 10906 26574 10908
rect 26278 10854 26324 10906
rect 26324 10854 26334 10906
rect 26358 10854 26388 10906
rect 26388 10854 26400 10906
rect 26400 10854 26414 10906
rect 26438 10854 26452 10906
rect 26452 10854 26464 10906
rect 26464 10854 26494 10906
rect 26518 10854 26528 10906
rect 26528 10854 26574 10906
rect 26278 10852 26334 10854
rect 26358 10852 26414 10854
rect 26438 10852 26494 10854
rect 26518 10852 26574 10854
rect 34719 10906 34775 10908
rect 34799 10906 34855 10908
rect 34879 10906 34935 10908
rect 34959 10906 35015 10908
rect 34719 10854 34765 10906
rect 34765 10854 34775 10906
rect 34799 10854 34829 10906
rect 34829 10854 34841 10906
rect 34841 10854 34855 10906
rect 34879 10854 34893 10906
rect 34893 10854 34905 10906
rect 34905 10854 34935 10906
rect 34959 10854 34969 10906
rect 34969 10854 35015 10906
rect 34719 10852 34775 10854
rect 34799 10852 34855 10854
rect 34879 10852 34935 10854
rect 34959 10852 35015 10854
rect 22058 10362 22114 10364
rect 22138 10362 22194 10364
rect 22218 10362 22274 10364
rect 22298 10362 22354 10364
rect 22058 10310 22104 10362
rect 22104 10310 22114 10362
rect 22138 10310 22168 10362
rect 22168 10310 22180 10362
rect 22180 10310 22194 10362
rect 22218 10310 22232 10362
rect 22232 10310 22244 10362
rect 22244 10310 22274 10362
rect 22298 10310 22308 10362
rect 22308 10310 22354 10362
rect 22058 10308 22114 10310
rect 22138 10308 22194 10310
rect 22218 10308 22274 10310
rect 22298 10308 22354 10310
rect 30499 10362 30555 10364
rect 30579 10362 30635 10364
rect 30659 10362 30715 10364
rect 30739 10362 30795 10364
rect 30499 10310 30545 10362
rect 30545 10310 30555 10362
rect 30579 10310 30609 10362
rect 30609 10310 30621 10362
rect 30621 10310 30635 10362
rect 30659 10310 30673 10362
rect 30673 10310 30685 10362
rect 30685 10310 30715 10362
rect 30739 10310 30749 10362
rect 30749 10310 30795 10362
rect 30499 10308 30555 10310
rect 30579 10308 30635 10310
rect 30659 10308 30715 10310
rect 30739 10308 30795 10310
rect 26278 9818 26334 9820
rect 26358 9818 26414 9820
rect 26438 9818 26494 9820
rect 26518 9818 26574 9820
rect 26278 9766 26324 9818
rect 26324 9766 26334 9818
rect 26358 9766 26388 9818
rect 26388 9766 26400 9818
rect 26400 9766 26414 9818
rect 26438 9766 26452 9818
rect 26452 9766 26464 9818
rect 26464 9766 26494 9818
rect 26518 9766 26528 9818
rect 26528 9766 26574 9818
rect 26278 9764 26334 9766
rect 26358 9764 26414 9766
rect 26438 9764 26494 9766
rect 26518 9764 26574 9766
rect 34719 9818 34775 9820
rect 34799 9818 34855 9820
rect 34879 9818 34935 9820
rect 34959 9818 35015 9820
rect 34719 9766 34765 9818
rect 34765 9766 34775 9818
rect 34799 9766 34829 9818
rect 34829 9766 34841 9818
rect 34841 9766 34855 9818
rect 34879 9766 34893 9818
rect 34893 9766 34905 9818
rect 34905 9766 34935 9818
rect 34959 9766 34969 9818
rect 34969 9766 35015 9818
rect 34719 9764 34775 9766
rect 34799 9764 34855 9766
rect 34879 9764 34935 9766
rect 34959 9764 35015 9766
rect 22058 9274 22114 9276
rect 22138 9274 22194 9276
rect 22218 9274 22274 9276
rect 22298 9274 22354 9276
rect 22058 9222 22104 9274
rect 22104 9222 22114 9274
rect 22138 9222 22168 9274
rect 22168 9222 22180 9274
rect 22180 9222 22194 9274
rect 22218 9222 22232 9274
rect 22232 9222 22244 9274
rect 22244 9222 22274 9274
rect 22298 9222 22308 9274
rect 22308 9222 22354 9274
rect 22058 9220 22114 9222
rect 22138 9220 22194 9222
rect 22218 9220 22274 9222
rect 22298 9220 22354 9222
rect 30499 9274 30555 9276
rect 30579 9274 30635 9276
rect 30659 9274 30715 9276
rect 30739 9274 30795 9276
rect 30499 9222 30545 9274
rect 30545 9222 30555 9274
rect 30579 9222 30609 9274
rect 30609 9222 30621 9274
rect 30621 9222 30635 9274
rect 30659 9222 30673 9274
rect 30673 9222 30685 9274
rect 30685 9222 30715 9274
rect 30739 9222 30749 9274
rect 30749 9222 30795 9274
rect 30499 9220 30555 9222
rect 30579 9220 30635 9222
rect 30659 9220 30715 9222
rect 30739 9220 30795 9222
rect 26278 8730 26334 8732
rect 26358 8730 26414 8732
rect 26438 8730 26494 8732
rect 26518 8730 26574 8732
rect 26278 8678 26324 8730
rect 26324 8678 26334 8730
rect 26358 8678 26388 8730
rect 26388 8678 26400 8730
rect 26400 8678 26414 8730
rect 26438 8678 26452 8730
rect 26452 8678 26464 8730
rect 26464 8678 26494 8730
rect 26518 8678 26528 8730
rect 26528 8678 26574 8730
rect 26278 8676 26334 8678
rect 26358 8676 26414 8678
rect 26438 8676 26494 8678
rect 26518 8676 26574 8678
rect 34719 8730 34775 8732
rect 34799 8730 34855 8732
rect 34879 8730 34935 8732
rect 34959 8730 35015 8732
rect 34719 8678 34765 8730
rect 34765 8678 34775 8730
rect 34799 8678 34829 8730
rect 34829 8678 34841 8730
rect 34841 8678 34855 8730
rect 34879 8678 34893 8730
rect 34893 8678 34905 8730
rect 34905 8678 34935 8730
rect 34959 8678 34969 8730
rect 34969 8678 35015 8730
rect 34719 8676 34775 8678
rect 34799 8676 34855 8678
rect 34879 8676 34935 8678
rect 34959 8676 35015 8678
rect 22058 8186 22114 8188
rect 22138 8186 22194 8188
rect 22218 8186 22274 8188
rect 22298 8186 22354 8188
rect 22058 8134 22104 8186
rect 22104 8134 22114 8186
rect 22138 8134 22168 8186
rect 22168 8134 22180 8186
rect 22180 8134 22194 8186
rect 22218 8134 22232 8186
rect 22232 8134 22244 8186
rect 22244 8134 22274 8186
rect 22298 8134 22308 8186
rect 22308 8134 22354 8186
rect 22058 8132 22114 8134
rect 22138 8132 22194 8134
rect 22218 8132 22274 8134
rect 22298 8132 22354 8134
rect 30499 8186 30555 8188
rect 30579 8186 30635 8188
rect 30659 8186 30715 8188
rect 30739 8186 30795 8188
rect 30499 8134 30545 8186
rect 30545 8134 30555 8186
rect 30579 8134 30609 8186
rect 30609 8134 30621 8186
rect 30621 8134 30635 8186
rect 30659 8134 30673 8186
rect 30673 8134 30685 8186
rect 30685 8134 30715 8186
rect 30739 8134 30749 8186
rect 30749 8134 30795 8186
rect 30499 8132 30555 8134
rect 30579 8132 30635 8134
rect 30659 8132 30715 8134
rect 30739 8132 30795 8134
rect 26278 7642 26334 7644
rect 26358 7642 26414 7644
rect 26438 7642 26494 7644
rect 26518 7642 26574 7644
rect 26278 7590 26324 7642
rect 26324 7590 26334 7642
rect 26358 7590 26388 7642
rect 26388 7590 26400 7642
rect 26400 7590 26414 7642
rect 26438 7590 26452 7642
rect 26452 7590 26464 7642
rect 26464 7590 26494 7642
rect 26518 7590 26528 7642
rect 26528 7590 26574 7642
rect 26278 7588 26334 7590
rect 26358 7588 26414 7590
rect 26438 7588 26494 7590
rect 26518 7588 26574 7590
rect 34719 7642 34775 7644
rect 34799 7642 34855 7644
rect 34879 7642 34935 7644
rect 34959 7642 35015 7644
rect 34719 7590 34765 7642
rect 34765 7590 34775 7642
rect 34799 7590 34829 7642
rect 34829 7590 34841 7642
rect 34841 7590 34855 7642
rect 34879 7590 34893 7642
rect 34893 7590 34905 7642
rect 34905 7590 34935 7642
rect 34959 7590 34969 7642
rect 34969 7590 35015 7642
rect 34719 7588 34775 7590
rect 34799 7588 34855 7590
rect 34879 7588 34935 7590
rect 34959 7588 35015 7590
rect 22058 7098 22114 7100
rect 22138 7098 22194 7100
rect 22218 7098 22274 7100
rect 22298 7098 22354 7100
rect 22058 7046 22104 7098
rect 22104 7046 22114 7098
rect 22138 7046 22168 7098
rect 22168 7046 22180 7098
rect 22180 7046 22194 7098
rect 22218 7046 22232 7098
rect 22232 7046 22244 7098
rect 22244 7046 22274 7098
rect 22298 7046 22308 7098
rect 22308 7046 22354 7098
rect 22058 7044 22114 7046
rect 22138 7044 22194 7046
rect 22218 7044 22274 7046
rect 22298 7044 22354 7046
rect 30499 7098 30555 7100
rect 30579 7098 30635 7100
rect 30659 7098 30715 7100
rect 30739 7098 30795 7100
rect 30499 7046 30545 7098
rect 30545 7046 30555 7098
rect 30579 7046 30609 7098
rect 30609 7046 30621 7098
rect 30621 7046 30635 7098
rect 30659 7046 30673 7098
rect 30673 7046 30685 7098
rect 30685 7046 30715 7098
rect 30739 7046 30749 7098
rect 30749 7046 30795 7098
rect 30499 7044 30555 7046
rect 30579 7044 30635 7046
rect 30659 7044 30715 7046
rect 30739 7044 30795 7046
rect 26278 6554 26334 6556
rect 26358 6554 26414 6556
rect 26438 6554 26494 6556
rect 26518 6554 26574 6556
rect 26278 6502 26324 6554
rect 26324 6502 26334 6554
rect 26358 6502 26388 6554
rect 26388 6502 26400 6554
rect 26400 6502 26414 6554
rect 26438 6502 26452 6554
rect 26452 6502 26464 6554
rect 26464 6502 26494 6554
rect 26518 6502 26528 6554
rect 26528 6502 26574 6554
rect 26278 6500 26334 6502
rect 26358 6500 26414 6502
rect 26438 6500 26494 6502
rect 26518 6500 26574 6502
rect 34719 6554 34775 6556
rect 34799 6554 34855 6556
rect 34879 6554 34935 6556
rect 34959 6554 35015 6556
rect 34719 6502 34765 6554
rect 34765 6502 34775 6554
rect 34799 6502 34829 6554
rect 34829 6502 34841 6554
rect 34841 6502 34855 6554
rect 34879 6502 34893 6554
rect 34893 6502 34905 6554
rect 34905 6502 34935 6554
rect 34959 6502 34969 6554
rect 34969 6502 35015 6554
rect 34719 6500 34775 6502
rect 34799 6500 34855 6502
rect 34879 6500 34935 6502
rect 34959 6500 35015 6502
rect 22058 6010 22114 6012
rect 22138 6010 22194 6012
rect 22218 6010 22274 6012
rect 22298 6010 22354 6012
rect 22058 5958 22104 6010
rect 22104 5958 22114 6010
rect 22138 5958 22168 6010
rect 22168 5958 22180 6010
rect 22180 5958 22194 6010
rect 22218 5958 22232 6010
rect 22232 5958 22244 6010
rect 22244 5958 22274 6010
rect 22298 5958 22308 6010
rect 22308 5958 22354 6010
rect 22058 5956 22114 5958
rect 22138 5956 22194 5958
rect 22218 5956 22274 5958
rect 22298 5956 22354 5958
rect 30499 6010 30555 6012
rect 30579 6010 30635 6012
rect 30659 6010 30715 6012
rect 30739 6010 30795 6012
rect 30499 5958 30545 6010
rect 30545 5958 30555 6010
rect 30579 5958 30609 6010
rect 30609 5958 30621 6010
rect 30621 5958 30635 6010
rect 30659 5958 30673 6010
rect 30673 5958 30685 6010
rect 30685 5958 30715 6010
rect 30739 5958 30749 6010
rect 30749 5958 30795 6010
rect 30499 5956 30555 5958
rect 30579 5956 30635 5958
rect 30659 5956 30715 5958
rect 30739 5956 30795 5958
rect 34518 5636 34574 5672
rect 34518 5616 34520 5636
rect 34520 5616 34572 5636
rect 34572 5616 34574 5636
rect 26278 5466 26334 5468
rect 26358 5466 26414 5468
rect 26438 5466 26494 5468
rect 26518 5466 26574 5468
rect 26278 5414 26324 5466
rect 26324 5414 26334 5466
rect 26358 5414 26388 5466
rect 26388 5414 26400 5466
rect 26400 5414 26414 5466
rect 26438 5414 26452 5466
rect 26452 5414 26464 5466
rect 26464 5414 26494 5466
rect 26518 5414 26528 5466
rect 26528 5414 26574 5466
rect 26278 5412 26334 5414
rect 26358 5412 26414 5414
rect 26438 5412 26494 5414
rect 26518 5412 26574 5414
rect 34719 5466 34775 5468
rect 34799 5466 34855 5468
rect 34879 5466 34935 5468
rect 34959 5466 35015 5468
rect 34719 5414 34765 5466
rect 34765 5414 34775 5466
rect 34799 5414 34829 5466
rect 34829 5414 34841 5466
rect 34841 5414 34855 5466
rect 34879 5414 34893 5466
rect 34893 5414 34905 5466
rect 34905 5414 34935 5466
rect 34959 5414 34969 5466
rect 34969 5414 35015 5466
rect 34719 5412 34775 5414
rect 34799 5412 34855 5414
rect 34879 5412 34935 5414
rect 34959 5412 35015 5414
rect 22058 4922 22114 4924
rect 22138 4922 22194 4924
rect 22218 4922 22274 4924
rect 22298 4922 22354 4924
rect 22058 4870 22104 4922
rect 22104 4870 22114 4922
rect 22138 4870 22168 4922
rect 22168 4870 22180 4922
rect 22180 4870 22194 4922
rect 22218 4870 22232 4922
rect 22232 4870 22244 4922
rect 22244 4870 22274 4922
rect 22298 4870 22308 4922
rect 22308 4870 22354 4922
rect 22058 4868 22114 4870
rect 22138 4868 22194 4870
rect 22218 4868 22274 4870
rect 22298 4868 22354 4870
rect 30499 4922 30555 4924
rect 30579 4922 30635 4924
rect 30659 4922 30715 4924
rect 30739 4922 30795 4924
rect 30499 4870 30545 4922
rect 30545 4870 30555 4922
rect 30579 4870 30609 4922
rect 30609 4870 30621 4922
rect 30621 4870 30635 4922
rect 30659 4870 30673 4922
rect 30673 4870 30685 4922
rect 30685 4870 30715 4922
rect 30739 4870 30749 4922
rect 30749 4870 30795 4922
rect 30499 4868 30555 4870
rect 30579 4868 30635 4870
rect 30659 4868 30715 4870
rect 30739 4868 30795 4870
rect 26278 4378 26334 4380
rect 26358 4378 26414 4380
rect 26438 4378 26494 4380
rect 26518 4378 26574 4380
rect 26278 4326 26324 4378
rect 26324 4326 26334 4378
rect 26358 4326 26388 4378
rect 26388 4326 26400 4378
rect 26400 4326 26414 4378
rect 26438 4326 26452 4378
rect 26452 4326 26464 4378
rect 26464 4326 26494 4378
rect 26518 4326 26528 4378
rect 26528 4326 26574 4378
rect 26278 4324 26334 4326
rect 26358 4324 26414 4326
rect 26438 4324 26494 4326
rect 26518 4324 26574 4326
rect 34719 4378 34775 4380
rect 34799 4378 34855 4380
rect 34879 4378 34935 4380
rect 34959 4378 35015 4380
rect 34719 4326 34765 4378
rect 34765 4326 34775 4378
rect 34799 4326 34829 4378
rect 34829 4326 34841 4378
rect 34841 4326 34855 4378
rect 34879 4326 34893 4378
rect 34893 4326 34905 4378
rect 34905 4326 34935 4378
rect 34959 4326 34969 4378
rect 34969 4326 35015 4378
rect 34719 4324 34775 4326
rect 34799 4324 34855 4326
rect 34879 4324 34935 4326
rect 34959 4324 35015 4326
rect 22058 3834 22114 3836
rect 22138 3834 22194 3836
rect 22218 3834 22274 3836
rect 22298 3834 22354 3836
rect 22058 3782 22104 3834
rect 22104 3782 22114 3834
rect 22138 3782 22168 3834
rect 22168 3782 22180 3834
rect 22180 3782 22194 3834
rect 22218 3782 22232 3834
rect 22232 3782 22244 3834
rect 22244 3782 22274 3834
rect 22298 3782 22308 3834
rect 22308 3782 22354 3834
rect 22058 3780 22114 3782
rect 22138 3780 22194 3782
rect 22218 3780 22274 3782
rect 22298 3780 22354 3782
rect 30499 3834 30555 3836
rect 30579 3834 30635 3836
rect 30659 3834 30715 3836
rect 30739 3834 30795 3836
rect 30499 3782 30545 3834
rect 30545 3782 30555 3834
rect 30579 3782 30609 3834
rect 30609 3782 30621 3834
rect 30621 3782 30635 3834
rect 30659 3782 30673 3834
rect 30673 3782 30685 3834
rect 30685 3782 30715 3834
rect 30739 3782 30749 3834
rect 30749 3782 30795 3834
rect 30499 3780 30555 3782
rect 30579 3780 30635 3782
rect 30659 3780 30715 3782
rect 30739 3780 30795 3782
rect 26278 3290 26334 3292
rect 26358 3290 26414 3292
rect 26438 3290 26494 3292
rect 26518 3290 26574 3292
rect 26278 3238 26324 3290
rect 26324 3238 26334 3290
rect 26358 3238 26388 3290
rect 26388 3238 26400 3290
rect 26400 3238 26414 3290
rect 26438 3238 26452 3290
rect 26452 3238 26464 3290
rect 26464 3238 26494 3290
rect 26518 3238 26528 3290
rect 26528 3238 26574 3290
rect 26278 3236 26334 3238
rect 26358 3236 26414 3238
rect 26438 3236 26494 3238
rect 26518 3236 26574 3238
rect 34719 3290 34775 3292
rect 34799 3290 34855 3292
rect 34879 3290 34935 3292
rect 34959 3290 35015 3292
rect 34719 3238 34765 3290
rect 34765 3238 34775 3290
rect 34799 3238 34829 3290
rect 34829 3238 34841 3290
rect 34841 3238 34855 3290
rect 34879 3238 34893 3290
rect 34893 3238 34905 3290
rect 34905 3238 34935 3290
rect 34959 3238 34969 3290
rect 34969 3238 35015 3290
rect 34719 3236 34775 3238
rect 34799 3236 34855 3238
rect 34879 3236 34935 3238
rect 34959 3236 35015 3238
rect 22058 2746 22114 2748
rect 22138 2746 22194 2748
rect 22218 2746 22274 2748
rect 22298 2746 22354 2748
rect 22058 2694 22104 2746
rect 22104 2694 22114 2746
rect 22138 2694 22168 2746
rect 22168 2694 22180 2746
rect 22180 2694 22194 2746
rect 22218 2694 22232 2746
rect 22232 2694 22244 2746
rect 22244 2694 22274 2746
rect 22298 2694 22308 2746
rect 22308 2694 22354 2746
rect 22058 2692 22114 2694
rect 22138 2692 22194 2694
rect 22218 2692 22274 2694
rect 22298 2692 22354 2694
rect 30499 2746 30555 2748
rect 30579 2746 30635 2748
rect 30659 2746 30715 2748
rect 30739 2746 30795 2748
rect 30499 2694 30545 2746
rect 30545 2694 30555 2746
rect 30579 2694 30609 2746
rect 30609 2694 30621 2746
rect 30621 2694 30635 2746
rect 30659 2694 30673 2746
rect 30673 2694 30685 2746
rect 30685 2694 30715 2746
rect 30739 2694 30749 2746
rect 30749 2694 30795 2746
rect 30499 2692 30555 2694
rect 30579 2692 30635 2694
rect 30659 2692 30715 2694
rect 30739 2692 30795 2694
rect 9396 2202 9452 2204
rect 9476 2202 9532 2204
rect 9556 2202 9612 2204
rect 9636 2202 9692 2204
rect 9396 2150 9442 2202
rect 9442 2150 9452 2202
rect 9476 2150 9506 2202
rect 9506 2150 9518 2202
rect 9518 2150 9532 2202
rect 9556 2150 9570 2202
rect 9570 2150 9582 2202
rect 9582 2150 9612 2202
rect 9636 2150 9646 2202
rect 9646 2150 9692 2202
rect 9396 2148 9452 2150
rect 9476 2148 9532 2150
rect 9556 2148 9612 2150
rect 9636 2148 9692 2150
rect 17837 2202 17893 2204
rect 17917 2202 17973 2204
rect 17997 2202 18053 2204
rect 18077 2202 18133 2204
rect 17837 2150 17883 2202
rect 17883 2150 17893 2202
rect 17917 2150 17947 2202
rect 17947 2150 17959 2202
rect 17959 2150 17973 2202
rect 17997 2150 18011 2202
rect 18011 2150 18023 2202
rect 18023 2150 18053 2202
rect 18077 2150 18087 2202
rect 18087 2150 18133 2202
rect 17837 2148 17893 2150
rect 17917 2148 17973 2150
rect 17997 2148 18053 2150
rect 18077 2148 18133 2150
rect 26278 2202 26334 2204
rect 26358 2202 26414 2204
rect 26438 2202 26494 2204
rect 26518 2202 26574 2204
rect 26278 2150 26324 2202
rect 26324 2150 26334 2202
rect 26358 2150 26388 2202
rect 26388 2150 26400 2202
rect 26400 2150 26414 2202
rect 26438 2150 26452 2202
rect 26452 2150 26464 2202
rect 26464 2150 26494 2202
rect 26518 2150 26528 2202
rect 26528 2150 26574 2202
rect 26278 2148 26334 2150
rect 26358 2148 26414 2150
rect 26438 2148 26494 2150
rect 26518 2148 26574 2150
rect 34719 2202 34775 2204
rect 34799 2202 34855 2204
rect 34879 2202 34935 2204
rect 34959 2202 35015 2204
rect 34719 2150 34765 2202
rect 34765 2150 34775 2202
rect 34799 2150 34829 2202
rect 34829 2150 34841 2202
rect 34841 2150 34855 2202
rect 34879 2150 34893 2202
rect 34893 2150 34905 2202
rect 34905 2150 34935 2202
rect 34959 2150 34969 2202
rect 34969 2150 35015 2202
rect 34719 2148 34775 2150
rect 34799 2148 34855 2150
rect 34879 2148 34935 2150
rect 34959 2148 35015 2150
<< metal3 >>
rect 5166 39744 5482 39745
rect 5166 39680 5172 39744
rect 5236 39680 5252 39744
rect 5316 39680 5332 39744
rect 5396 39680 5412 39744
rect 5476 39680 5482 39744
rect 5166 39679 5482 39680
rect 13607 39744 13923 39745
rect 13607 39680 13613 39744
rect 13677 39680 13693 39744
rect 13757 39680 13773 39744
rect 13837 39680 13853 39744
rect 13917 39680 13923 39744
rect 13607 39679 13923 39680
rect 22048 39744 22364 39745
rect 22048 39680 22054 39744
rect 22118 39680 22134 39744
rect 22198 39680 22214 39744
rect 22278 39680 22294 39744
rect 22358 39680 22364 39744
rect 22048 39679 22364 39680
rect 30489 39744 30805 39745
rect 30489 39680 30495 39744
rect 30559 39680 30575 39744
rect 30639 39680 30655 39744
rect 30719 39680 30735 39744
rect 30799 39680 30805 39744
rect 30489 39679 30805 39680
rect 9386 39200 9702 39201
rect 9386 39136 9392 39200
rect 9456 39136 9472 39200
rect 9536 39136 9552 39200
rect 9616 39136 9632 39200
rect 9696 39136 9702 39200
rect 9386 39135 9702 39136
rect 17827 39200 18143 39201
rect 17827 39136 17833 39200
rect 17897 39136 17913 39200
rect 17977 39136 17993 39200
rect 18057 39136 18073 39200
rect 18137 39136 18143 39200
rect 17827 39135 18143 39136
rect 26268 39200 26584 39201
rect 26268 39136 26274 39200
rect 26338 39136 26354 39200
rect 26418 39136 26434 39200
rect 26498 39136 26514 39200
rect 26578 39136 26584 39200
rect 26268 39135 26584 39136
rect 34709 39200 35025 39201
rect 34709 39136 34715 39200
rect 34779 39136 34795 39200
rect 34859 39136 34875 39200
rect 34939 39136 34955 39200
rect 35019 39136 35025 39200
rect 34709 39135 35025 39136
rect 5166 38656 5482 38657
rect 5166 38592 5172 38656
rect 5236 38592 5252 38656
rect 5316 38592 5332 38656
rect 5396 38592 5412 38656
rect 5476 38592 5482 38656
rect 5166 38591 5482 38592
rect 13607 38656 13923 38657
rect 13607 38592 13613 38656
rect 13677 38592 13693 38656
rect 13757 38592 13773 38656
rect 13837 38592 13853 38656
rect 13917 38592 13923 38656
rect 13607 38591 13923 38592
rect 22048 38656 22364 38657
rect 22048 38592 22054 38656
rect 22118 38592 22134 38656
rect 22198 38592 22214 38656
rect 22278 38592 22294 38656
rect 22358 38592 22364 38656
rect 22048 38591 22364 38592
rect 30489 38656 30805 38657
rect 30489 38592 30495 38656
rect 30559 38592 30575 38656
rect 30639 38592 30655 38656
rect 30719 38592 30735 38656
rect 30799 38592 30805 38656
rect 30489 38591 30805 38592
rect 9386 38112 9702 38113
rect 9386 38048 9392 38112
rect 9456 38048 9472 38112
rect 9536 38048 9552 38112
rect 9616 38048 9632 38112
rect 9696 38048 9702 38112
rect 9386 38047 9702 38048
rect 17827 38112 18143 38113
rect 17827 38048 17833 38112
rect 17897 38048 17913 38112
rect 17977 38048 17993 38112
rect 18057 38048 18073 38112
rect 18137 38048 18143 38112
rect 17827 38047 18143 38048
rect 26268 38112 26584 38113
rect 26268 38048 26274 38112
rect 26338 38048 26354 38112
rect 26418 38048 26434 38112
rect 26498 38048 26514 38112
rect 26578 38048 26584 38112
rect 26268 38047 26584 38048
rect 34709 38112 35025 38113
rect 34709 38048 34715 38112
rect 34779 38048 34795 38112
rect 34859 38048 34875 38112
rect 34939 38048 34955 38112
rect 35019 38048 35025 38112
rect 34709 38047 35025 38048
rect 5166 37568 5482 37569
rect 5166 37504 5172 37568
rect 5236 37504 5252 37568
rect 5316 37504 5332 37568
rect 5396 37504 5412 37568
rect 5476 37504 5482 37568
rect 5166 37503 5482 37504
rect 13607 37568 13923 37569
rect 13607 37504 13613 37568
rect 13677 37504 13693 37568
rect 13757 37504 13773 37568
rect 13837 37504 13853 37568
rect 13917 37504 13923 37568
rect 13607 37503 13923 37504
rect 22048 37568 22364 37569
rect 22048 37504 22054 37568
rect 22118 37504 22134 37568
rect 22198 37504 22214 37568
rect 22278 37504 22294 37568
rect 22358 37504 22364 37568
rect 22048 37503 22364 37504
rect 30489 37568 30805 37569
rect 30489 37504 30495 37568
rect 30559 37504 30575 37568
rect 30639 37504 30655 37568
rect 30719 37504 30735 37568
rect 30799 37504 30805 37568
rect 30489 37503 30805 37504
rect 9386 37024 9702 37025
rect 9386 36960 9392 37024
rect 9456 36960 9472 37024
rect 9536 36960 9552 37024
rect 9616 36960 9632 37024
rect 9696 36960 9702 37024
rect 9386 36959 9702 36960
rect 17827 37024 18143 37025
rect 17827 36960 17833 37024
rect 17897 36960 17913 37024
rect 17977 36960 17993 37024
rect 18057 36960 18073 37024
rect 18137 36960 18143 37024
rect 17827 36959 18143 36960
rect 26268 37024 26584 37025
rect 26268 36960 26274 37024
rect 26338 36960 26354 37024
rect 26418 36960 26434 37024
rect 26498 36960 26514 37024
rect 26578 36960 26584 37024
rect 26268 36959 26584 36960
rect 34709 37024 35025 37025
rect 34709 36960 34715 37024
rect 34779 36960 34795 37024
rect 34859 36960 34875 37024
rect 34939 36960 34955 37024
rect 35019 36960 35025 37024
rect 34709 36959 35025 36960
rect 5166 36480 5482 36481
rect 5166 36416 5172 36480
rect 5236 36416 5252 36480
rect 5316 36416 5332 36480
rect 5396 36416 5412 36480
rect 5476 36416 5482 36480
rect 5166 36415 5482 36416
rect 13607 36480 13923 36481
rect 13607 36416 13613 36480
rect 13677 36416 13693 36480
rect 13757 36416 13773 36480
rect 13837 36416 13853 36480
rect 13917 36416 13923 36480
rect 13607 36415 13923 36416
rect 22048 36480 22364 36481
rect 22048 36416 22054 36480
rect 22118 36416 22134 36480
rect 22198 36416 22214 36480
rect 22278 36416 22294 36480
rect 22358 36416 22364 36480
rect 22048 36415 22364 36416
rect 30489 36480 30805 36481
rect 30489 36416 30495 36480
rect 30559 36416 30575 36480
rect 30639 36416 30655 36480
rect 30719 36416 30735 36480
rect 30799 36416 30805 36480
rect 30489 36415 30805 36416
rect 0 36138 800 36228
rect 933 36138 999 36141
rect 0 36136 999 36138
rect 0 36080 938 36136
rect 994 36080 999 36136
rect 0 36078 999 36080
rect 0 35988 800 36078
rect 933 36075 999 36078
rect 15469 36138 15535 36141
rect 18505 36138 18571 36141
rect 15469 36136 18571 36138
rect 15469 36080 15474 36136
rect 15530 36080 18510 36136
rect 18566 36080 18571 36136
rect 15469 36078 18571 36080
rect 15469 36075 15535 36078
rect 18505 36075 18571 36078
rect 9386 35936 9702 35937
rect 9386 35872 9392 35936
rect 9456 35872 9472 35936
rect 9536 35872 9552 35936
rect 9616 35872 9632 35936
rect 9696 35872 9702 35936
rect 9386 35871 9702 35872
rect 17827 35936 18143 35937
rect 17827 35872 17833 35936
rect 17897 35872 17913 35936
rect 17977 35872 17993 35936
rect 18057 35872 18073 35936
rect 18137 35872 18143 35936
rect 17827 35871 18143 35872
rect 26268 35936 26584 35937
rect 26268 35872 26274 35936
rect 26338 35872 26354 35936
rect 26418 35872 26434 35936
rect 26498 35872 26514 35936
rect 26578 35872 26584 35936
rect 26268 35871 26584 35872
rect 34709 35936 35025 35937
rect 34709 35872 34715 35936
rect 34779 35872 34795 35936
rect 34859 35872 34875 35936
rect 34939 35872 34955 35936
rect 35019 35872 35025 35936
rect 34709 35871 35025 35872
rect 5166 35392 5482 35393
rect 5166 35328 5172 35392
rect 5236 35328 5252 35392
rect 5316 35328 5332 35392
rect 5396 35328 5412 35392
rect 5476 35328 5482 35392
rect 5166 35327 5482 35328
rect 13607 35392 13923 35393
rect 13607 35328 13613 35392
rect 13677 35328 13693 35392
rect 13757 35328 13773 35392
rect 13837 35328 13853 35392
rect 13917 35328 13923 35392
rect 13607 35327 13923 35328
rect 22048 35392 22364 35393
rect 22048 35328 22054 35392
rect 22118 35328 22134 35392
rect 22198 35328 22214 35392
rect 22278 35328 22294 35392
rect 22358 35328 22364 35392
rect 22048 35327 22364 35328
rect 30489 35392 30805 35393
rect 30489 35328 30495 35392
rect 30559 35328 30575 35392
rect 30639 35328 30655 35392
rect 30719 35328 30735 35392
rect 30799 35328 30805 35392
rect 30489 35327 30805 35328
rect 11513 35050 11579 35053
rect 19149 35050 19215 35053
rect 11513 35048 19215 35050
rect 11513 34992 11518 35048
rect 11574 34992 19154 35048
rect 19210 34992 19215 35048
rect 11513 34990 19215 34992
rect 11513 34987 11579 34990
rect 19149 34987 19215 34990
rect 9386 34848 9702 34849
rect 9386 34784 9392 34848
rect 9456 34784 9472 34848
rect 9536 34784 9552 34848
rect 9616 34784 9632 34848
rect 9696 34784 9702 34848
rect 9386 34783 9702 34784
rect 17827 34848 18143 34849
rect 17827 34784 17833 34848
rect 17897 34784 17913 34848
rect 17977 34784 17993 34848
rect 18057 34784 18073 34848
rect 18137 34784 18143 34848
rect 17827 34783 18143 34784
rect 26268 34848 26584 34849
rect 26268 34784 26274 34848
rect 26338 34784 26354 34848
rect 26418 34784 26434 34848
rect 26498 34784 26514 34848
rect 26578 34784 26584 34848
rect 26268 34783 26584 34784
rect 34709 34848 35025 34849
rect 34709 34784 34715 34848
rect 34779 34784 34795 34848
rect 34859 34784 34875 34848
rect 34939 34784 34955 34848
rect 35019 34784 35025 34848
rect 34709 34783 35025 34784
rect 35200 34781 36000 34868
rect 35157 34776 36000 34781
rect 35157 34720 35162 34776
rect 35218 34720 36000 34776
rect 35157 34715 36000 34720
rect 11881 34642 11947 34645
rect 15193 34642 15259 34645
rect 11881 34640 15259 34642
rect 11881 34584 11886 34640
rect 11942 34584 15198 34640
rect 15254 34584 15259 34640
rect 11881 34582 15259 34584
rect 11881 34579 11947 34582
rect 15193 34579 15259 34582
rect 15653 34642 15719 34645
rect 16481 34642 16547 34645
rect 18781 34642 18847 34645
rect 15653 34640 18847 34642
rect 15653 34584 15658 34640
rect 15714 34584 16486 34640
rect 16542 34584 18786 34640
rect 18842 34584 18847 34640
rect 35200 34628 36000 34715
rect 15653 34582 18847 34584
rect 15653 34579 15719 34582
rect 16481 34579 16547 34582
rect 18781 34579 18847 34582
rect 5166 34304 5482 34305
rect 5166 34240 5172 34304
rect 5236 34240 5252 34304
rect 5316 34240 5332 34304
rect 5396 34240 5412 34304
rect 5476 34240 5482 34304
rect 5166 34239 5482 34240
rect 13607 34304 13923 34305
rect 13607 34240 13613 34304
rect 13677 34240 13693 34304
rect 13757 34240 13773 34304
rect 13837 34240 13853 34304
rect 13917 34240 13923 34304
rect 13607 34239 13923 34240
rect 22048 34304 22364 34305
rect 22048 34240 22054 34304
rect 22118 34240 22134 34304
rect 22198 34240 22214 34304
rect 22278 34240 22294 34304
rect 22358 34240 22364 34304
rect 22048 34239 22364 34240
rect 30489 34304 30805 34305
rect 30489 34240 30495 34304
rect 30559 34240 30575 34304
rect 30639 34240 30655 34304
rect 30719 34240 30735 34304
rect 30799 34240 30805 34304
rect 30489 34239 30805 34240
rect 9386 33760 9702 33761
rect 9386 33696 9392 33760
rect 9456 33696 9472 33760
rect 9536 33696 9552 33760
rect 9616 33696 9632 33760
rect 9696 33696 9702 33760
rect 9386 33695 9702 33696
rect 17827 33760 18143 33761
rect 17827 33696 17833 33760
rect 17897 33696 17913 33760
rect 17977 33696 17993 33760
rect 18057 33696 18073 33760
rect 18137 33696 18143 33760
rect 17827 33695 18143 33696
rect 26268 33760 26584 33761
rect 26268 33696 26274 33760
rect 26338 33696 26354 33760
rect 26418 33696 26434 33760
rect 26498 33696 26514 33760
rect 26578 33696 26584 33760
rect 26268 33695 26584 33696
rect 34709 33760 35025 33761
rect 34709 33696 34715 33760
rect 34779 33696 34795 33760
rect 34859 33696 34875 33760
rect 34939 33696 34955 33760
rect 35019 33696 35025 33760
rect 34709 33695 35025 33696
rect 5166 33216 5482 33217
rect 5166 33152 5172 33216
rect 5236 33152 5252 33216
rect 5316 33152 5332 33216
rect 5396 33152 5412 33216
rect 5476 33152 5482 33216
rect 5166 33151 5482 33152
rect 13607 33216 13923 33217
rect 13607 33152 13613 33216
rect 13677 33152 13693 33216
rect 13757 33152 13773 33216
rect 13837 33152 13853 33216
rect 13917 33152 13923 33216
rect 13607 33151 13923 33152
rect 22048 33216 22364 33217
rect 22048 33152 22054 33216
rect 22118 33152 22134 33216
rect 22198 33152 22214 33216
rect 22278 33152 22294 33216
rect 22358 33152 22364 33216
rect 22048 33151 22364 33152
rect 30489 33216 30805 33217
rect 30489 33152 30495 33216
rect 30559 33152 30575 33216
rect 30639 33152 30655 33216
rect 30719 33152 30735 33216
rect 30799 33152 30805 33216
rect 30489 33151 30805 33152
rect 14825 33010 14891 33013
rect 14782 33008 14891 33010
rect 14782 32952 14830 33008
rect 14886 32952 14891 33008
rect 14782 32947 14891 32952
rect 9386 32672 9702 32673
rect 9386 32608 9392 32672
rect 9456 32608 9472 32672
rect 9536 32608 9552 32672
rect 9616 32608 9632 32672
rect 9696 32608 9702 32672
rect 9386 32607 9702 32608
rect 10225 32602 10291 32605
rect 10501 32602 10567 32605
rect 10225 32600 10567 32602
rect 10225 32544 10230 32600
rect 10286 32544 10506 32600
rect 10562 32544 10567 32600
rect 10225 32542 10567 32544
rect 10225 32539 10291 32542
rect 10501 32539 10567 32542
rect 14782 32469 14842 32947
rect 16573 32874 16639 32877
rect 17861 32874 17927 32877
rect 16573 32872 17927 32874
rect 16573 32816 16578 32872
rect 16634 32816 17866 32872
rect 17922 32816 17927 32872
rect 16573 32814 17927 32816
rect 16573 32811 16639 32814
rect 17861 32811 17927 32814
rect 18137 32874 18203 32877
rect 19517 32874 19583 32877
rect 18137 32872 19583 32874
rect 18137 32816 18142 32872
rect 18198 32816 19522 32872
rect 19578 32816 19583 32872
rect 18137 32814 19583 32816
rect 18137 32811 18203 32814
rect 19517 32811 19583 32814
rect 17827 32672 18143 32673
rect 17827 32608 17833 32672
rect 17897 32608 17913 32672
rect 17977 32608 17993 32672
rect 18057 32608 18073 32672
rect 18137 32608 18143 32672
rect 17827 32607 18143 32608
rect 26268 32672 26584 32673
rect 26268 32608 26274 32672
rect 26338 32608 26354 32672
rect 26418 32608 26434 32672
rect 26498 32608 26514 32672
rect 26578 32608 26584 32672
rect 26268 32607 26584 32608
rect 34709 32672 35025 32673
rect 34709 32608 34715 32672
rect 34779 32608 34795 32672
rect 34859 32608 34875 32672
rect 34939 32608 34955 32672
rect 35019 32608 35025 32672
rect 34709 32607 35025 32608
rect 9949 32466 10015 32469
rect 10685 32466 10751 32469
rect 9949 32464 10751 32466
rect 9949 32408 9954 32464
rect 10010 32408 10690 32464
rect 10746 32408 10751 32464
rect 9949 32406 10751 32408
rect 9949 32403 10015 32406
rect 10685 32403 10751 32406
rect 14733 32464 14842 32469
rect 14733 32408 14738 32464
rect 14794 32408 14842 32464
rect 14733 32406 14842 32408
rect 17585 32466 17651 32469
rect 19149 32466 19215 32469
rect 17585 32464 19215 32466
rect 17585 32408 17590 32464
rect 17646 32408 19154 32464
rect 19210 32408 19215 32464
rect 17585 32406 19215 32408
rect 14733 32403 14799 32406
rect 17585 32403 17651 32406
rect 19149 32403 19215 32406
rect 13997 32330 14063 32333
rect 15285 32330 15351 32333
rect 18229 32330 18295 32333
rect 19425 32330 19491 32333
rect 13997 32328 19491 32330
rect 13997 32272 14002 32328
rect 14058 32272 15290 32328
rect 15346 32272 18234 32328
rect 18290 32272 19430 32328
rect 19486 32272 19491 32328
rect 13997 32270 19491 32272
rect 13997 32267 14063 32270
rect 15285 32267 15351 32270
rect 18229 32267 18295 32270
rect 19425 32267 19491 32270
rect 5166 32128 5482 32129
rect 5166 32064 5172 32128
rect 5236 32064 5252 32128
rect 5316 32064 5332 32128
rect 5396 32064 5412 32128
rect 5476 32064 5482 32128
rect 5166 32063 5482 32064
rect 13607 32128 13923 32129
rect 13607 32064 13613 32128
rect 13677 32064 13693 32128
rect 13757 32064 13773 32128
rect 13837 32064 13853 32128
rect 13917 32064 13923 32128
rect 13607 32063 13923 32064
rect 22048 32128 22364 32129
rect 22048 32064 22054 32128
rect 22118 32064 22134 32128
rect 22198 32064 22214 32128
rect 22278 32064 22294 32128
rect 22358 32064 22364 32128
rect 22048 32063 22364 32064
rect 30489 32128 30805 32129
rect 30489 32064 30495 32128
rect 30559 32064 30575 32128
rect 30639 32064 30655 32128
rect 30719 32064 30735 32128
rect 30799 32064 30805 32128
rect 30489 32063 30805 32064
rect 9386 31584 9702 31585
rect 9386 31520 9392 31584
rect 9456 31520 9472 31584
rect 9536 31520 9552 31584
rect 9616 31520 9632 31584
rect 9696 31520 9702 31584
rect 9386 31519 9702 31520
rect 17827 31584 18143 31585
rect 17827 31520 17833 31584
rect 17897 31520 17913 31584
rect 17977 31520 17993 31584
rect 18057 31520 18073 31584
rect 18137 31520 18143 31584
rect 17827 31519 18143 31520
rect 26268 31584 26584 31585
rect 26268 31520 26274 31584
rect 26338 31520 26354 31584
rect 26418 31520 26434 31584
rect 26498 31520 26514 31584
rect 26578 31520 26584 31584
rect 26268 31519 26584 31520
rect 34709 31584 35025 31585
rect 34709 31520 34715 31584
rect 34779 31520 34795 31584
rect 34859 31520 34875 31584
rect 34939 31520 34955 31584
rect 35019 31520 35025 31584
rect 34709 31519 35025 31520
rect 5166 31040 5482 31041
rect 5166 30976 5172 31040
rect 5236 30976 5252 31040
rect 5316 30976 5332 31040
rect 5396 30976 5412 31040
rect 5476 30976 5482 31040
rect 5166 30975 5482 30976
rect 13607 31040 13923 31041
rect 13607 30976 13613 31040
rect 13677 30976 13693 31040
rect 13757 30976 13773 31040
rect 13837 30976 13853 31040
rect 13917 30976 13923 31040
rect 13607 30975 13923 30976
rect 22048 31040 22364 31041
rect 22048 30976 22054 31040
rect 22118 30976 22134 31040
rect 22198 30976 22214 31040
rect 22278 30976 22294 31040
rect 22358 30976 22364 31040
rect 22048 30975 22364 30976
rect 30489 31040 30805 31041
rect 30489 30976 30495 31040
rect 30559 30976 30575 31040
rect 30639 30976 30655 31040
rect 30719 30976 30735 31040
rect 30799 30976 30805 31040
rect 30489 30975 30805 30976
rect 9386 30496 9702 30497
rect 9386 30432 9392 30496
rect 9456 30432 9472 30496
rect 9536 30432 9552 30496
rect 9616 30432 9632 30496
rect 9696 30432 9702 30496
rect 9386 30431 9702 30432
rect 17827 30496 18143 30497
rect 17827 30432 17833 30496
rect 17897 30432 17913 30496
rect 17977 30432 17993 30496
rect 18057 30432 18073 30496
rect 18137 30432 18143 30496
rect 17827 30431 18143 30432
rect 26268 30496 26584 30497
rect 26268 30432 26274 30496
rect 26338 30432 26354 30496
rect 26418 30432 26434 30496
rect 26498 30432 26514 30496
rect 26578 30432 26584 30496
rect 26268 30431 26584 30432
rect 34709 30496 35025 30497
rect 34709 30432 34715 30496
rect 34779 30432 34795 30496
rect 34859 30432 34875 30496
rect 34939 30432 34955 30496
rect 35019 30432 35025 30496
rect 34709 30431 35025 30432
rect 18321 30426 18387 30429
rect 19977 30426 20043 30429
rect 20529 30426 20595 30429
rect 18321 30424 20595 30426
rect 18321 30368 18326 30424
rect 18382 30368 19982 30424
rect 20038 30368 20534 30424
rect 20590 30368 20595 30424
rect 18321 30366 20595 30368
rect 18321 30363 18387 30366
rect 19977 30363 20043 30366
rect 20529 30363 20595 30366
rect 5166 29952 5482 29953
rect 5166 29888 5172 29952
rect 5236 29888 5252 29952
rect 5316 29888 5332 29952
rect 5396 29888 5412 29952
rect 5476 29888 5482 29952
rect 5166 29887 5482 29888
rect 13607 29952 13923 29953
rect 13607 29888 13613 29952
rect 13677 29888 13693 29952
rect 13757 29888 13773 29952
rect 13837 29888 13853 29952
rect 13917 29888 13923 29952
rect 13607 29887 13923 29888
rect 22048 29952 22364 29953
rect 22048 29888 22054 29952
rect 22118 29888 22134 29952
rect 22198 29888 22214 29952
rect 22278 29888 22294 29952
rect 22358 29888 22364 29952
rect 22048 29887 22364 29888
rect 30489 29952 30805 29953
rect 30489 29888 30495 29952
rect 30559 29888 30575 29952
rect 30639 29888 30655 29952
rect 30719 29888 30735 29952
rect 30799 29888 30805 29952
rect 30489 29887 30805 29888
rect 15929 29610 15995 29613
rect 18137 29610 18203 29613
rect 15929 29608 18203 29610
rect 15929 29552 15934 29608
rect 15990 29552 18142 29608
rect 18198 29552 18203 29608
rect 15929 29550 18203 29552
rect 15929 29547 15995 29550
rect 18137 29547 18203 29550
rect 9386 29408 9702 29409
rect 9386 29344 9392 29408
rect 9456 29344 9472 29408
rect 9536 29344 9552 29408
rect 9616 29344 9632 29408
rect 9696 29344 9702 29408
rect 9386 29343 9702 29344
rect 17827 29408 18143 29409
rect 17827 29344 17833 29408
rect 17897 29344 17913 29408
rect 17977 29344 17993 29408
rect 18057 29344 18073 29408
rect 18137 29344 18143 29408
rect 17827 29343 18143 29344
rect 26268 29408 26584 29409
rect 26268 29344 26274 29408
rect 26338 29344 26354 29408
rect 26418 29344 26434 29408
rect 26498 29344 26514 29408
rect 26578 29344 26584 29408
rect 26268 29343 26584 29344
rect 34709 29408 35025 29409
rect 34709 29344 34715 29408
rect 34779 29344 34795 29408
rect 34859 29344 34875 29408
rect 34939 29344 34955 29408
rect 35019 29344 35025 29408
rect 34709 29343 35025 29344
rect 17493 29202 17559 29205
rect 19333 29202 19399 29205
rect 17493 29200 19399 29202
rect 17493 29144 17498 29200
rect 17554 29144 19338 29200
rect 19394 29144 19399 29200
rect 17493 29142 19399 29144
rect 17493 29139 17559 29142
rect 19333 29139 19399 29142
rect 1393 28930 1459 28933
rect 798 28928 1459 28930
rect 798 28872 1398 28928
rect 1454 28872 1459 28928
rect 798 28870 1459 28872
rect 798 28748 858 28870
rect 1393 28867 1459 28870
rect 5166 28864 5482 28865
rect 5166 28800 5172 28864
rect 5236 28800 5252 28864
rect 5316 28800 5332 28864
rect 5396 28800 5412 28864
rect 5476 28800 5482 28864
rect 5166 28799 5482 28800
rect 13607 28864 13923 28865
rect 13607 28800 13613 28864
rect 13677 28800 13693 28864
rect 13757 28800 13773 28864
rect 13837 28800 13853 28864
rect 13917 28800 13923 28864
rect 13607 28799 13923 28800
rect 22048 28864 22364 28865
rect 22048 28800 22054 28864
rect 22118 28800 22134 28864
rect 22198 28800 22214 28864
rect 22278 28800 22294 28864
rect 22358 28800 22364 28864
rect 22048 28799 22364 28800
rect 30489 28864 30805 28865
rect 30489 28800 30495 28864
rect 30559 28800 30575 28864
rect 30639 28800 30655 28864
rect 30719 28800 30735 28864
rect 30799 28800 30805 28864
rect 30489 28799 30805 28800
rect 0 28598 858 28748
rect 0 28508 800 28598
rect 9386 28320 9702 28321
rect 9386 28256 9392 28320
rect 9456 28256 9472 28320
rect 9536 28256 9552 28320
rect 9616 28256 9632 28320
rect 9696 28256 9702 28320
rect 9386 28255 9702 28256
rect 17827 28320 18143 28321
rect 17827 28256 17833 28320
rect 17897 28256 17913 28320
rect 17977 28256 17993 28320
rect 18057 28256 18073 28320
rect 18137 28256 18143 28320
rect 17827 28255 18143 28256
rect 26268 28320 26584 28321
rect 26268 28256 26274 28320
rect 26338 28256 26354 28320
rect 26418 28256 26434 28320
rect 26498 28256 26514 28320
rect 26578 28256 26584 28320
rect 26268 28255 26584 28256
rect 34709 28320 35025 28321
rect 34709 28256 34715 28320
rect 34779 28256 34795 28320
rect 34859 28256 34875 28320
rect 34939 28256 34955 28320
rect 35019 28256 35025 28320
rect 34709 28255 35025 28256
rect 5166 27776 5482 27777
rect 5166 27712 5172 27776
rect 5236 27712 5252 27776
rect 5316 27712 5332 27776
rect 5396 27712 5412 27776
rect 5476 27712 5482 27776
rect 5166 27711 5482 27712
rect 13607 27776 13923 27777
rect 13607 27712 13613 27776
rect 13677 27712 13693 27776
rect 13757 27712 13773 27776
rect 13837 27712 13853 27776
rect 13917 27712 13923 27776
rect 13607 27711 13923 27712
rect 22048 27776 22364 27777
rect 22048 27712 22054 27776
rect 22118 27712 22134 27776
rect 22198 27712 22214 27776
rect 22278 27712 22294 27776
rect 22358 27712 22364 27776
rect 22048 27711 22364 27712
rect 30489 27776 30805 27777
rect 30489 27712 30495 27776
rect 30559 27712 30575 27776
rect 30639 27712 30655 27776
rect 30719 27712 30735 27776
rect 30799 27712 30805 27776
rect 30489 27711 30805 27712
rect 34513 27434 34579 27437
rect 34513 27432 35220 27434
rect 34513 27376 34518 27432
rect 34574 27388 35220 27432
rect 34574 27376 36000 27388
rect 34513 27374 36000 27376
rect 34513 27371 34579 27374
rect 35160 27238 36000 27374
rect 9386 27232 9702 27233
rect 9386 27168 9392 27232
rect 9456 27168 9472 27232
rect 9536 27168 9552 27232
rect 9616 27168 9632 27232
rect 9696 27168 9702 27232
rect 9386 27167 9702 27168
rect 17827 27232 18143 27233
rect 17827 27168 17833 27232
rect 17897 27168 17913 27232
rect 17977 27168 17993 27232
rect 18057 27168 18073 27232
rect 18137 27168 18143 27232
rect 17827 27167 18143 27168
rect 26268 27232 26584 27233
rect 26268 27168 26274 27232
rect 26338 27168 26354 27232
rect 26418 27168 26434 27232
rect 26498 27168 26514 27232
rect 26578 27168 26584 27232
rect 26268 27167 26584 27168
rect 34709 27232 35025 27233
rect 34709 27168 34715 27232
rect 34779 27168 34795 27232
rect 34859 27168 34875 27232
rect 34939 27168 34955 27232
rect 35019 27168 35025 27232
rect 34709 27167 35025 27168
rect 19793 27162 19859 27165
rect 21725 27162 21791 27165
rect 19793 27160 21791 27162
rect 19793 27104 19798 27160
rect 19854 27104 21730 27160
rect 21786 27104 21791 27160
rect 35200 27148 36000 27238
rect 19793 27102 21791 27104
rect 19793 27099 19859 27102
rect 21725 27099 21791 27102
rect 5166 26688 5482 26689
rect 5166 26624 5172 26688
rect 5236 26624 5252 26688
rect 5316 26624 5332 26688
rect 5396 26624 5412 26688
rect 5476 26624 5482 26688
rect 5166 26623 5482 26624
rect 13607 26688 13923 26689
rect 13607 26624 13613 26688
rect 13677 26624 13693 26688
rect 13757 26624 13773 26688
rect 13837 26624 13853 26688
rect 13917 26624 13923 26688
rect 13607 26623 13923 26624
rect 22048 26688 22364 26689
rect 22048 26624 22054 26688
rect 22118 26624 22134 26688
rect 22198 26624 22214 26688
rect 22278 26624 22294 26688
rect 22358 26624 22364 26688
rect 22048 26623 22364 26624
rect 30489 26688 30805 26689
rect 30489 26624 30495 26688
rect 30559 26624 30575 26688
rect 30639 26624 30655 26688
rect 30719 26624 30735 26688
rect 30799 26624 30805 26688
rect 30489 26623 30805 26624
rect 21081 26482 21147 26485
rect 24577 26482 24643 26485
rect 21081 26480 24643 26482
rect 21081 26424 21086 26480
rect 21142 26424 24582 26480
rect 24638 26424 24643 26480
rect 21081 26422 24643 26424
rect 21081 26419 21147 26422
rect 24577 26419 24643 26422
rect 9386 26144 9702 26145
rect 9386 26080 9392 26144
rect 9456 26080 9472 26144
rect 9536 26080 9552 26144
rect 9616 26080 9632 26144
rect 9696 26080 9702 26144
rect 9386 26079 9702 26080
rect 17827 26144 18143 26145
rect 17827 26080 17833 26144
rect 17897 26080 17913 26144
rect 17977 26080 17993 26144
rect 18057 26080 18073 26144
rect 18137 26080 18143 26144
rect 17827 26079 18143 26080
rect 26268 26144 26584 26145
rect 26268 26080 26274 26144
rect 26338 26080 26354 26144
rect 26418 26080 26434 26144
rect 26498 26080 26514 26144
rect 26578 26080 26584 26144
rect 26268 26079 26584 26080
rect 34709 26144 35025 26145
rect 34709 26080 34715 26144
rect 34779 26080 34795 26144
rect 34859 26080 34875 26144
rect 34939 26080 34955 26144
rect 35019 26080 35025 26144
rect 34709 26079 35025 26080
rect 5166 25600 5482 25601
rect 5166 25536 5172 25600
rect 5236 25536 5252 25600
rect 5316 25536 5332 25600
rect 5396 25536 5412 25600
rect 5476 25536 5482 25600
rect 5166 25535 5482 25536
rect 13607 25600 13923 25601
rect 13607 25536 13613 25600
rect 13677 25536 13693 25600
rect 13757 25536 13773 25600
rect 13837 25536 13853 25600
rect 13917 25536 13923 25600
rect 13607 25535 13923 25536
rect 22048 25600 22364 25601
rect 22048 25536 22054 25600
rect 22118 25536 22134 25600
rect 22198 25536 22214 25600
rect 22278 25536 22294 25600
rect 22358 25536 22364 25600
rect 22048 25535 22364 25536
rect 30489 25600 30805 25601
rect 30489 25536 30495 25600
rect 30559 25536 30575 25600
rect 30639 25536 30655 25600
rect 30719 25536 30735 25600
rect 30799 25536 30805 25600
rect 30489 25535 30805 25536
rect 9386 25056 9702 25057
rect 9386 24992 9392 25056
rect 9456 24992 9472 25056
rect 9536 24992 9552 25056
rect 9616 24992 9632 25056
rect 9696 24992 9702 25056
rect 9386 24991 9702 24992
rect 17827 25056 18143 25057
rect 17827 24992 17833 25056
rect 17897 24992 17913 25056
rect 17977 24992 17993 25056
rect 18057 24992 18073 25056
rect 18137 24992 18143 25056
rect 17827 24991 18143 24992
rect 26268 25056 26584 25057
rect 26268 24992 26274 25056
rect 26338 24992 26354 25056
rect 26418 24992 26434 25056
rect 26498 24992 26514 25056
rect 26578 24992 26584 25056
rect 26268 24991 26584 24992
rect 34709 25056 35025 25057
rect 34709 24992 34715 25056
rect 34779 24992 34795 25056
rect 34859 24992 34875 25056
rect 34939 24992 34955 25056
rect 35019 24992 35025 25056
rect 34709 24991 35025 24992
rect 5166 24512 5482 24513
rect 5166 24448 5172 24512
rect 5236 24448 5252 24512
rect 5316 24448 5332 24512
rect 5396 24448 5412 24512
rect 5476 24448 5482 24512
rect 5166 24447 5482 24448
rect 13607 24512 13923 24513
rect 13607 24448 13613 24512
rect 13677 24448 13693 24512
rect 13757 24448 13773 24512
rect 13837 24448 13853 24512
rect 13917 24448 13923 24512
rect 13607 24447 13923 24448
rect 22048 24512 22364 24513
rect 22048 24448 22054 24512
rect 22118 24448 22134 24512
rect 22198 24448 22214 24512
rect 22278 24448 22294 24512
rect 22358 24448 22364 24512
rect 22048 24447 22364 24448
rect 30489 24512 30805 24513
rect 30489 24448 30495 24512
rect 30559 24448 30575 24512
rect 30639 24448 30655 24512
rect 30719 24448 30735 24512
rect 30799 24448 30805 24512
rect 30489 24447 30805 24448
rect 9386 23968 9702 23969
rect 9386 23904 9392 23968
rect 9456 23904 9472 23968
rect 9536 23904 9552 23968
rect 9616 23904 9632 23968
rect 9696 23904 9702 23968
rect 9386 23903 9702 23904
rect 17827 23968 18143 23969
rect 17827 23904 17833 23968
rect 17897 23904 17913 23968
rect 17977 23904 17993 23968
rect 18057 23904 18073 23968
rect 18137 23904 18143 23968
rect 17827 23903 18143 23904
rect 26268 23968 26584 23969
rect 26268 23904 26274 23968
rect 26338 23904 26354 23968
rect 26418 23904 26434 23968
rect 26498 23904 26514 23968
rect 26578 23904 26584 23968
rect 26268 23903 26584 23904
rect 34709 23968 35025 23969
rect 34709 23904 34715 23968
rect 34779 23904 34795 23968
rect 34859 23904 34875 23968
rect 34939 23904 34955 23968
rect 35019 23904 35025 23968
rect 34709 23903 35025 23904
rect 13721 23762 13787 23765
rect 15561 23762 15627 23765
rect 13721 23760 15627 23762
rect 13721 23704 13726 23760
rect 13782 23704 15566 23760
rect 15622 23704 15627 23760
rect 13721 23702 15627 23704
rect 13721 23699 13787 23702
rect 15561 23699 15627 23702
rect 22277 23626 22343 23629
rect 23013 23626 23079 23629
rect 22277 23624 23079 23626
rect 22277 23568 22282 23624
rect 22338 23568 23018 23624
rect 23074 23568 23079 23624
rect 22277 23566 23079 23568
rect 22277 23563 22343 23566
rect 23013 23563 23079 23566
rect 5166 23424 5482 23425
rect 5166 23360 5172 23424
rect 5236 23360 5252 23424
rect 5316 23360 5332 23424
rect 5396 23360 5412 23424
rect 5476 23360 5482 23424
rect 5166 23359 5482 23360
rect 13607 23424 13923 23425
rect 13607 23360 13613 23424
rect 13677 23360 13693 23424
rect 13757 23360 13773 23424
rect 13837 23360 13853 23424
rect 13917 23360 13923 23424
rect 13607 23359 13923 23360
rect 22048 23424 22364 23425
rect 22048 23360 22054 23424
rect 22118 23360 22134 23424
rect 22198 23360 22214 23424
rect 22278 23360 22294 23424
rect 22358 23360 22364 23424
rect 22048 23359 22364 23360
rect 30489 23424 30805 23425
rect 30489 23360 30495 23424
rect 30559 23360 30575 23424
rect 30639 23360 30655 23424
rect 30719 23360 30735 23424
rect 30799 23360 30805 23424
rect 30489 23359 30805 23360
rect 20529 23218 20595 23221
rect 24485 23218 24551 23221
rect 20529 23216 24551 23218
rect 20529 23160 20534 23216
rect 20590 23160 24490 23216
rect 24546 23160 24551 23216
rect 20529 23158 24551 23160
rect 20529 23155 20595 23158
rect 24485 23155 24551 23158
rect 20805 22946 20871 22949
rect 22369 22946 22435 22949
rect 20805 22944 22435 22946
rect 20805 22888 20810 22944
rect 20866 22888 22374 22944
rect 22430 22888 22435 22944
rect 20805 22886 22435 22888
rect 20805 22883 20871 22886
rect 22369 22883 22435 22886
rect 9386 22880 9702 22881
rect 9386 22816 9392 22880
rect 9456 22816 9472 22880
rect 9536 22816 9552 22880
rect 9616 22816 9632 22880
rect 9696 22816 9702 22880
rect 9386 22815 9702 22816
rect 17827 22880 18143 22881
rect 17827 22816 17833 22880
rect 17897 22816 17913 22880
rect 17977 22816 17993 22880
rect 18057 22816 18073 22880
rect 18137 22816 18143 22880
rect 17827 22815 18143 22816
rect 26268 22880 26584 22881
rect 26268 22816 26274 22880
rect 26338 22816 26354 22880
rect 26418 22816 26434 22880
rect 26498 22816 26514 22880
rect 26578 22816 26584 22880
rect 26268 22815 26584 22816
rect 34709 22880 35025 22881
rect 34709 22816 34715 22880
rect 34779 22816 34795 22880
rect 34859 22816 34875 22880
rect 34939 22816 34955 22880
rect 35019 22816 35025 22880
rect 34709 22815 35025 22816
rect 22001 22810 22067 22813
rect 23841 22810 23907 22813
rect 22001 22808 23907 22810
rect 22001 22752 22006 22808
rect 22062 22752 23846 22808
rect 23902 22752 23907 22808
rect 22001 22750 23907 22752
rect 22001 22747 22067 22750
rect 23841 22747 23907 22750
rect 5166 22336 5482 22337
rect 5166 22272 5172 22336
rect 5236 22272 5252 22336
rect 5316 22272 5332 22336
rect 5396 22272 5412 22336
rect 5476 22272 5482 22336
rect 5166 22271 5482 22272
rect 13607 22336 13923 22337
rect 13607 22272 13613 22336
rect 13677 22272 13693 22336
rect 13757 22272 13773 22336
rect 13837 22272 13853 22336
rect 13917 22272 13923 22336
rect 13607 22271 13923 22272
rect 22048 22336 22364 22337
rect 22048 22272 22054 22336
rect 22118 22272 22134 22336
rect 22198 22272 22214 22336
rect 22278 22272 22294 22336
rect 22358 22272 22364 22336
rect 22048 22271 22364 22272
rect 30489 22336 30805 22337
rect 30489 22272 30495 22336
rect 30559 22272 30575 22336
rect 30639 22272 30655 22336
rect 30719 22272 30735 22336
rect 30799 22272 30805 22336
rect 30489 22271 30805 22272
rect 0 21858 800 21948
rect 933 21858 999 21861
rect 0 21856 999 21858
rect 0 21800 938 21856
rect 994 21800 999 21856
rect 0 21798 999 21800
rect 0 21708 800 21798
rect 933 21795 999 21798
rect 9386 21792 9702 21793
rect 9386 21728 9392 21792
rect 9456 21728 9472 21792
rect 9536 21728 9552 21792
rect 9616 21728 9632 21792
rect 9696 21728 9702 21792
rect 9386 21727 9702 21728
rect 17827 21792 18143 21793
rect 17827 21728 17833 21792
rect 17897 21728 17913 21792
rect 17977 21728 17993 21792
rect 18057 21728 18073 21792
rect 18137 21728 18143 21792
rect 17827 21727 18143 21728
rect 26268 21792 26584 21793
rect 26268 21728 26274 21792
rect 26338 21728 26354 21792
rect 26418 21728 26434 21792
rect 26498 21728 26514 21792
rect 26578 21728 26584 21792
rect 26268 21727 26584 21728
rect 34709 21792 35025 21793
rect 34709 21728 34715 21792
rect 34779 21728 34795 21792
rect 34859 21728 34875 21792
rect 34939 21728 34955 21792
rect 35019 21728 35025 21792
rect 34709 21727 35025 21728
rect 5166 21248 5482 21249
rect 5166 21184 5172 21248
rect 5236 21184 5252 21248
rect 5316 21184 5332 21248
rect 5396 21184 5412 21248
rect 5476 21184 5482 21248
rect 5166 21183 5482 21184
rect 13607 21248 13923 21249
rect 13607 21184 13613 21248
rect 13677 21184 13693 21248
rect 13757 21184 13773 21248
rect 13837 21184 13853 21248
rect 13917 21184 13923 21248
rect 13607 21183 13923 21184
rect 22048 21248 22364 21249
rect 22048 21184 22054 21248
rect 22118 21184 22134 21248
rect 22198 21184 22214 21248
rect 22278 21184 22294 21248
rect 22358 21184 22364 21248
rect 22048 21183 22364 21184
rect 30489 21248 30805 21249
rect 30489 21184 30495 21248
rect 30559 21184 30575 21248
rect 30639 21184 30655 21248
rect 30719 21184 30735 21248
rect 30799 21184 30805 21248
rect 30489 21183 30805 21184
rect 9386 20704 9702 20705
rect 9386 20640 9392 20704
rect 9456 20640 9472 20704
rect 9536 20640 9552 20704
rect 9616 20640 9632 20704
rect 9696 20640 9702 20704
rect 9386 20639 9702 20640
rect 17827 20704 18143 20705
rect 17827 20640 17833 20704
rect 17897 20640 17913 20704
rect 17977 20640 17993 20704
rect 18057 20640 18073 20704
rect 18137 20640 18143 20704
rect 17827 20639 18143 20640
rect 26268 20704 26584 20705
rect 26268 20640 26274 20704
rect 26338 20640 26354 20704
rect 26418 20640 26434 20704
rect 26498 20640 26514 20704
rect 26578 20640 26584 20704
rect 26268 20639 26584 20640
rect 34709 20704 35025 20705
rect 34709 20640 34715 20704
rect 34779 20640 34795 20704
rect 34859 20640 34875 20704
rect 34939 20640 34955 20704
rect 35019 20640 35025 20704
rect 34709 20639 35025 20640
rect 5166 20160 5482 20161
rect 5166 20096 5172 20160
rect 5236 20096 5252 20160
rect 5316 20096 5332 20160
rect 5396 20096 5412 20160
rect 5476 20096 5482 20160
rect 5166 20095 5482 20096
rect 13607 20160 13923 20161
rect 13607 20096 13613 20160
rect 13677 20096 13693 20160
rect 13757 20096 13773 20160
rect 13837 20096 13853 20160
rect 13917 20096 13923 20160
rect 13607 20095 13923 20096
rect 22048 20160 22364 20161
rect 22048 20096 22054 20160
rect 22118 20096 22134 20160
rect 22198 20096 22214 20160
rect 22278 20096 22294 20160
rect 22358 20096 22364 20160
rect 22048 20095 22364 20096
rect 30489 20160 30805 20161
rect 30489 20096 30495 20160
rect 30559 20096 30575 20160
rect 30639 20096 30655 20160
rect 30719 20096 30735 20160
rect 30799 20096 30805 20160
rect 30489 20095 30805 20096
rect 34605 19818 34671 19821
rect 35200 19818 36000 19908
rect 34605 19816 36000 19818
rect 34605 19760 34610 19816
rect 34666 19760 36000 19816
rect 34605 19758 36000 19760
rect 34605 19755 34671 19758
rect 35200 19668 36000 19758
rect 9386 19616 9702 19617
rect 9386 19552 9392 19616
rect 9456 19552 9472 19616
rect 9536 19552 9552 19616
rect 9616 19552 9632 19616
rect 9696 19552 9702 19616
rect 9386 19551 9702 19552
rect 17827 19616 18143 19617
rect 17827 19552 17833 19616
rect 17897 19552 17913 19616
rect 17977 19552 17993 19616
rect 18057 19552 18073 19616
rect 18137 19552 18143 19616
rect 17827 19551 18143 19552
rect 26268 19616 26584 19617
rect 26268 19552 26274 19616
rect 26338 19552 26354 19616
rect 26418 19552 26434 19616
rect 26498 19552 26514 19616
rect 26578 19552 26584 19616
rect 26268 19551 26584 19552
rect 34709 19616 35025 19617
rect 34709 19552 34715 19616
rect 34779 19552 34795 19616
rect 34859 19552 34875 19616
rect 34939 19552 34955 19616
rect 35019 19552 35025 19616
rect 34709 19551 35025 19552
rect 5166 19072 5482 19073
rect 5166 19008 5172 19072
rect 5236 19008 5252 19072
rect 5316 19008 5332 19072
rect 5396 19008 5412 19072
rect 5476 19008 5482 19072
rect 5166 19007 5482 19008
rect 13607 19072 13923 19073
rect 13607 19008 13613 19072
rect 13677 19008 13693 19072
rect 13757 19008 13773 19072
rect 13837 19008 13853 19072
rect 13917 19008 13923 19072
rect 13607 19007 13923 19008
rect 22048 19072 22364 19073
rect 22048 19008 22054 19072
rect 22118 19008 22134 19072
rect 22198 19008 22214 19072
rect 22278 19008 22294 19072
rect 22358 19008 22364 19072
rect 22048 19007 22364 19008
rect 30489 19072 30805 19073
rect 30489 19008 30495 19072
rect 30559 19008 30575 19072
rect 30639 19008 30655 19072
rect 30719 19008 30735 19072
rect 30799 19008 30805 19072
rect 30489 19007 30805 19008
rect 9386 18528 9702 18529
rect 9386 18464 9392 18528
rect 9456 18464 9472 18528
rect 9536 18464 9552 18528
rect 9616 18464 9632 18528
rect 9696 18464 9702 18528
rect 9386 18463 9702 18464
rect 17827 18528 18143 18529
rect 17827 18464 17833 18528
rect 17897 18464 17913 18528
rect 17977 18464 17993 18528
rect 18057 18464 18073 18528
rect 18137 18464 18143 18528
rect 17827 18463 18143 18464
rect 26268 18528 26584 18529
rect 26268 18464 26274 18528
rect 26338 18464 26354 18528
rect 26418 18464 26434 18528
rect 26498 18464 26514 18528
rect 26578 18464 26584 18528
rect 26268 18463 26584 18464
rect 34709 18528 35025 18529
rect 34709 18464 34715 18528
rect 34779 18464 34795 18528
rect 34859 18464 34875 18528
rect 34939 18464 34955 18528
rect 35019 18464 35025 18528
rect 34709 18463 35025 18464
rect 5166 17984 5482 17985
rect 5166 17920 5172 17984
rect 5236 17920 5252 17984
rect 5316 17920 5332 17984
rect 5396 17920 5412 17984
rect 5476 17920 5482 17984
rect 5166 17919 5482 17920
rect 13607 17984 13923 17985
rect 13607 17920 13613 17984
rect 13677 17920 13693 17984
rect 13757 17920 13773 17984
rect 13837 17920 13853 17984
rect 13917 17920 13923 17984
rect 13607 17919 13923 17920
rect 22048 17984 22364 17985
rect 22048 17920 22054 17984
rect 22118 17920 22134 17984
rect 22198 17920 22214 17984
rect 22278 17920 22294 17984
rect 22358 17920 22364 17984
rect 22048 17919 22364 17920
rect 30489 17984 30805 17985
rect 30489 17920 30495 17984
rect 30559 17920 30575 17984
rect 30639 17920 30655 17984
rect 30719 17920 30735 17984
rect 30799 17920 30805 17984
rect 30489 17919 30805 17920
rect 9386 17440 9702 17441
rect 9386 17376 9392 17440
rect 9456 17376 9472 17440
rect 9536 17376 9552 17440
rect 9616 17376 9632 17440
rect 9696 17376 9702 17440
rect 9386 17375 9702 17376
rect 17827 17440 18143 17441
rect 17827 17376 17833 17440
rect 17897 17376 17913 17440
rect 17977 17376 17993 17440
rect 18057 17376 18073 17440
rect 18137 17376 18143 17440
rect 17827 17375 18143 17376
rect 26268 17440 26584 17441
rect 26268 17376 26274 17440
rect 26338 17376 26354 17440
rect 26418 17376 26434 17440
rect 26498 17376 26514 17440
rect 26578 17376 26584 17440
rect 26268 17375 26584 17376
rect 34709 17440 35025 17441
rect 34709 17376 34715 17440
rect 34779 17376 34795 17440
rect 34859 17376 34875 17440
rect 34939 17376 34955 17440
rect 35019 17376 35025 17440
rect 34709 17375 35025 17376
rect 5166 16896 5482 16897
rect 5166 16832 5172 16896
rect 5236 16832 5252 16896
rect 5316 16832 5332 16896
rect 5396 16832 5412 16896
rect 5476 16832 5482 16896
rect 5166 16831 5482 16832
rect 13607 16896 13923 16897
rect 13607 16832 13613 16896
rect 13677 16832 13693 16896
rect 13757 16832 13773 16896
rect 13837 16832 13853 16896
rect 13917 16832 13923 16896
rect 13607 16831 13923 16832
rect 22048 16896 22364 16897
rect 22048 16832 22054 16896
rect 22118 16832 22134 16896
rect 22198 16832 22214 16896
rect 22278 16832 22294 16896
rect 22358 16832 22364 16896
rect 22048 16831 22364 16832
rect 30489 16896 30805 16897
rect 30489 16832 30495 16896
rect 30559 16832 30575 16896
rect 30639 16832 30655 16896
rect 30719 16832 30735 16896
rect 30799 16832 30805 16896
rect 30489 16831 30805 16832
rect 9386 16352 9702 16353
rect 9386 16288 9392 16352
rect 9456 16288 9472 16352
rect 9536 16288 9552 16352
rect 9616 16288 9632 16352
rect 9696 16288 9702 16352
rect 9386 16287 9702 16288
rect 17827 16352 18143 16353
rect 17827 16288 17833 16352
rect 17897 16288 17913 16352
rect 17977 16288 17993 16352
rect 18057 16288 18073 16352
rect 18137 16288 18143 16352
rect 17827 16287 18143 16288
rect 26268 16352 26584 16353
rect 26268 16288 26274 16352
rect 26338 16288 26354 16352
rect 26418 16288 26434 16352
rect 26498 16288 26514 16352
rect 26578 16288 26584 16352
rect 26268 16287 26584 16288
rect 34709 16352 35025 16353
rect 34709 16288 34715 16352
rect 34779 16288 34795 16352
rect 34859 16288 34875 16352
rect 34939 16288 34955 16352
rect 35019 16288 35025 16352
rect 34709 16287 35025 16288
rect 5166 15808 5482 15809
rect 5166 15744 5172 15808
rect 5236 15744 5252 15808
rect 5316 15744 5332 15808
rect 5396 15744 5412 15808
rect 5476 15744 5482 15808
rect 5166 15743 5482 15744
rect 13607 15808 13923 15809
rect 13607 15744 13613 15808
rect 13677 15744 13693 15808
rect 13757 15744 13773 15808
rect 13837 15744 13853 15808
rect 13917 15744 13923 15808
rect 13607 15743 13923 15744
rect 22048 15808 22364 15809
rect 22048 15744 22054 15808
rect 22118 15744 22134 15808
rect 22198 15744 22214 15808
rect 22278 15744 22294 15808
rect 22358 15744 22364 15808
rect 22048 15743 22364 15744
rect 30489 15808 30805 15809
rect 30489 15744 30495 15808
rect 30559 15744 30575 15808
rect 30639 15744 30655 15808
rect 30719 15744 30735 15808
rect 30799 15744 30805 15808
rect 30489 15743 30805 15744
rect 9386 15264 9702 15265
rect 9386 15200 9392 15264
rect 9456 15200 9472 15264
rect 9536 15200 9552 15264
rect 9616 15200 9632 15264
rect 9696 15200 9702 15264
rect 9386 15199 9702 15200
rect 17827 15264 18143 15265
rect 17827 15200 17833 15264
rect 17897 15200 17913 15264
rect 17977 15200 17993 15264
rect 18057 15200 18073 15264
rect 18137 15200 18143 15264
rect 17827 15199 18143 15200
rect 26268 15264 26584 15265
rect 26268 15200 26274 15264
rect 26338 15200 26354 15264
rect 26418 15200 26434 15264
rect 26498 15200 26514 15264
rect 26578 15200 26584 15264
rect 26268 15199 26584 15200
rect 34709 15264 35025 15265
rect 34709 15200 34715 15264
rect 34779 15200 34795 15264
rect 34859 15200 34875 15264
rect 34939 15200 34955 15264
rect 35019 15200 35025 15264
rect 34709 15199 35025 15200
rect 5166 14720 5482 14721
rect 5166 14656 5172 14720
rect 5236 14656 5252 14720
rect 5316 14656 5332 14720
rect 5396 14656 5412 14720
rect 5476 14656 5482 14720
rect 5166 14655 5482 14656
rect 13607 14720 13923 14721
rect 13607 14656 13613 14720
rect 13677 14656 13693 14720
rect 13757 14656 13773 14720
rect 13837 14656 13853 14720
rect 13917 14656 13923 14720
rect 13607 14655 13923 14656
rect 22048 14720 22364 14721
rect 22048 14656 22054 14720
rect 22118 14656 22134 14720
rect 22198 14656 22214 14720
rect 22278 14656 22294 14720
rect 22358 14656 22364 14720
rect 22048 14655 22364 14656
rect 30489 14720 30805 14721
rect 30489 14656 30495 14720
rect 30559 14656 30575 14720
rect 30639 14656 30655 14720
rect 30719 14656 30735 14720
rect 30799 14656 30805 14720
rect 30489 14655 30805 14656
rect 0 14378 800 14468
rect 933 14378 999 14381
rect 0 14376 999 14378
rect 0 14320 938 14376
rect 994 14320 999 14376
rect 0 14318 999 14320
rect 0 14228 800 14318
rect 933 14315 999 14318
rect 9386 14176 9702 14177
rect 9386 14112 9392 14176
rect 9456 14112 9472 14176
rect 9536 14112 9552 14176
rect 9616 14112 9632 14176
rect 9696 14112 9702 14176
rect 9386 14111 9702 14112
rect 17827 14176 18143 14177
rect 17827 14112 17833 14176
rect 17897 14112 17913 14176
rect 17977 14112 17993 14176
rect 18057 14112 18073 14176
rect 18137 14112 18143 14176
rect 17827 14111 18143 14112
rect 26268 14176 26584 14177
rect 26268 14112 26274 14176
rect 26338 14112 26354 14176
rect 26418 14112 26434 14176
rect 26498 14112 26514 14176
rect 26578 14112 26584 14176
rect 26268 14111 26584 14112
rect 34709 14176 35025 14177
rect 34709 14112 34715 14176
rect 34779 14112 34795 14176
rect 34859 14112 34875 14176
rect 34939 14112 34955 14176
rect 35019 14112 35025 14176
rect 34709 14111 35025 14112
rect 5166 13632 5482 13633
rect 5166 13568 5172 13632
rect 5236 13568 5252 13632
rect 5316 13568 5332 13632
rect 5396 13568 5412 13632
rect 5476 13568 5482 13632
rect 5166 13567 5482 13568
rect 13607 13632 13923 13633
rect 13607 13568 13613 13632
rect 13677 13568 13693 13632
rect 13757 13568 13773 13632
rect 13837 13568 13853 13632
rect 13917 13568 13923 13632
rect 13607 13567 13923 13568
rect 22048 13632 22364 13633
rect 22048 13568 22054 13632
rect 22118 13568 22134 13632
rect 22198 13568 22214 13632
rect 22278 13568 22294 13632
rect 22358 13568 22364 13632
rect 22048 13567 22364 13568
rect 30489 13632 30805 13633
rect 30489 13568 30495 13632
rect 30559 13568 30575 13632
rect 30639 13568 30655 13632
rect 30719 13568 30735 13632
rect 30799 13568 30805 13632
rect 30489 13567 30805 13568
rect 9386 13088 9702 13089
rect 9386 13024 9392 13088
rect 9456 13024 9472 13088
rect 9536 13024 9552 13088
rect 9616 13024 9632 13088
rect 9696 13024 9702 13088
rect 9386 13023 9702 13024
rect 17827 13088 18143 13089
rect 17827 13024 17833 13088
rect 17897 13024 17913 13088
rect 17977 13024 17993 13088
rect 18057 13024 18073 13088
rect 18137 13024 18143 13088
rect 17827 13023 18143 13024
rect 26268 13088 26584 13089
rect 26268 13024 26274 13088
rect 26338 13024 26354 13088
rect 26418 13024 26434 13088
rect 26498 13024 26514 13088
rect 26578 13024 26584 13088
rect 26268 13023 26584 13024
rect 34709 13088 35025 13089
rect 34709 13024 34715 13088
rect 34779 13024 34795 13088
rect 34859 13024 34875 13088
rect 34939 13024 34955 13088
rect 35019 13024 35025 13088
rect 34709 13023 35025 13024
rect 35200 13021 36000 13108
rect 35157 13016 36000 13021
rect 35157 12960 35162 13016
rect 35218 12960 36000 13016
rect 35157 12955 36000 12960
rect 35200 12868 36000 12955
rect 5166 12544 5482 12545
rect 5166 12480 5172 12544
rect 5236 12480 5252 12544
rect 5316 12480 5332 12544
rect 5396 12480 5412 12544
rect 5476 12480 5482 12544
rect 5166 12479 5482 12480
rect 13607 12544 13923 12545
rect 13607 12480 13613 12544
rect 13677 12480 13693 12544
rect 13757 12480 13773 12544
rect 13837 12480 13853 12544
rect 13917 12480 13923 12544
rect 13607 12479 13923 12480
rect 22048 12544 22364 12545
rect 22048 12480 22054 12544
rect 22118 12480 22134 12544
rect 22198 12480 22214 12544
rect 22278 12480 22294 12544
rect 22358 12480 22364 12544
rect 22048 12479 22364 12480
rect 30489 12544 30805 12545
rect 30489 12480 30495 12544
rect 30559 12480 30575 12544
rect 30639 12480 30655 12544
rect 30719 12480 30735 12544
rect 30799 12480 30805 12544
rect 30489 12479 30805 12480
rect 9386 12000 9702 12001
rect 9386 11936 9392 12000
rect 9456 11936 9472 12000
rect 9536 11936 9552 12000
rect 9616 11936 9632 12000
rect 9696 11936 9702 12000
rect 9386 11935 9702 11936
rect 17827 12000 18143 12001
rect 17827 11936 17833 12000
rect 17897 11936 17913 12000
rect 17977 11936 17993 12000
rect 18057 11936 18073 12000
rect 18137 11936 18143 12000
rect 17827 11935 18143 11936
rect 26268 12000 26584 12001
rect 26268 11936 26274 12000
rect 26338 11936 26354 12000
rect 26418 11936 26434 12000
rect 26498 11936 26514 12000
rect 26578 11936 26584 12000
rect 26268 11935 26584 11936
rect 34709 12000 35025 12001
rect 34709 11936 34715 12000
rect 34779 11936 34795 12000
rect 34859 11936 34875 12000
rect 34939 11936 34955 12000
rect 35019 11936 35025 12000
rect 34709 11935 35025 11936
rect 5166 11456 5482 11457
rect 5166 11392 5172 11456
rect 5236 11392 5252 11456
rect 5316 11392 5332 11456
rect 5396 11392 5412 11456
rect 5476 11392 5482 11456
rect 5166 11391 5482 11392
rect 13607 11456 13923 11457
rect 13607 11392 13613 11456
rect 13677 11392 13693 11456
rect 13757 11392 13773 11456
rect 13837 11392 13853 11456
rect 13917 11392 13923 11456
rect 13607 11391 13923 11392
rect 22048 11456 22364 11457
rect 22048 11392 22054 11456
rect 22118 11392 22134 11456
rect 22198 11392 22214 11456
rect 22278 11392 22294 11456
rect 22358 11392 22364 11456
rect 22048 11391 22364 11392
rect 30489 11456 30805 11457
rect 30489 11392 30495 11456
rect 30559 11392 30575 11456
rect 30639 11392 30655 11456
rect 30719 11392 30735 11456
rect 30799 11392 30805 11456
rect 30489 11391 30805 11392
rect 9386 10912 9702 10913
rect 9386 10848 9392 10912
rect 9456 10848 9472 10912
rect 9536 10848 9552 10912
rect 9616 10848 9632 10912
rect 9696 10848 9702 10912
rect 9386 10847 9702 10848
rect 17827 10912 18143 10913
rect 17827 10848 17833 10912
rect 17897 10848 17913 10912
rect 17977 10848 17993 10912
rect 18057 10848 18073 10912
rect 18137 10848 18143 10912
rect 17827 10847 18143 10848
rect 26268 10912 26584 10913
rect 26268 10848 26274 10912
rect 26338 10848 26354 10912
rect 26418 10848 26434 10912
rect 26498 10848 26514 10912
rect 26578 10848 26584 10912
rect 26268 10847 26584 10848
rect 34709 10912 35025 10913
rect 34709 10848 34715 10912
rect 34779 10848 34795 10912
rect 34859 10848 34875 10912
rect 34939 10848 34955 10912
rect 35019 10848 35025 10912
rect 34709 10847 35025 10848
rect 5166 10368 5482 10369
rect 5166 10304 5172 10368
rect 5236 10304 5252 10368
rect 5316 10304 5332 10368
rect 5396 10304 5412 10368
rect 5476 10304 5482 10368
rect 5166 10303 5482 10304
rect 13607 10368 13923 10369
rect 13607 10304 13613 10368
rect 13677 10304 13693 10368
rect 13757 10304 13773 10368
rect 13837 10304 13853 10368
rect 13917 10304 13923 10368
rect 13607 10303 13923 10304
rect 22048 10368 22364 10369
rect 22048 10304 22054 10368
rect 22118 10304 22134 10368
rect 22198 10304 22214 10368
rect 22278 10304 22294 10368
rect 22358 10304 22364 10368
rect 22048 10303 22364 10304
rect 30489 10368 30805 10369
rect 30489 10304 30495 10368
rect 30559 10304 30575 10368
rect 30639 10304 30655 10368
rect 30719 10304 30735 10368
rect 30799 10304 30805 10368
rect 30489 10303 30805 10304
rect 9386 9824 9702 9825
rect 9386 9760 9392 9824
rect 9456 9760 9472 9824
rect 9536 9760 9552 9824
rect 9616 9760 9632 9824
rect 9696 9760 9702 9824
rect 9386 9759 9702 9760
rect 17827 9824 18143 9825
rect 17827 9760 17833 9824
rect 17897 9760 17913 9824
rect 17977 9760 17993 9824
rect 18057 9760 18073 9824
rect 18137 9760 18143 9824
rect 17827 9759 18143 9760
rect 26268 9824 26584 9825
rect 26268 9760 26274 9824
rect 26338 9760 26354 9824
rect 26418 9760 26434 9824
rect 26498 9760 26514 9824
rect 26578 9760 26584 9824
rect 26268 9759 26584 9760
rect 34709 9824 35025 9825
rect 34709 9760 34715 9824
rect 34779 9760 34795 9824
rect 34859 9760 34875 9824
rect 34939 9760 34955 9824
rect 35019 9760 35025 9824
rect 34709 9759 35025 9760
rect 5166 9280 5482 9281
rect 5166 9216 5172 9280
rect 5236 9216 5252 9280
rect 5316 9216 5332 9280
rect 5396 9216 5412 9280
rect 5476 9216 5482 9280
rect 5166 9215 5482 9216
rect 13607 9280 13923 9281
rect 13607 9216 13613 9280
rect 13677 9216 13693 9280
rect 13757 9216 13773 9280
rect 13837 9216 13853 9280
rect 13917 9216 13923 9280
rect 13607 9215 13923 9216
rect 22048 9280 22364 9281
rect 22048 9216 22054 9280
rect 22118 9216 22134 9280
rect 22198 9216 22214 9280
rect 22278 9216 22294 9280
rect 22358 9216 22364 9280
rect 22048 9215 22364 9216
rect 30489 9280 30805 9281
rect 30489 9216 30495 9280
rect 30559 9216 30575 9280
rect 30639 9216 30655 9280
rect 30719 9216 30735 9280
rect 30799 9216 30805 9280
rect 30489 9215 30805 9216
rect 9386 8736 9702 8737
rect 9386 8672 9392 8736
rect 9456 8672 9472 8736
rect 9536 8672 9552 8736
rect 9616 8672 9632 8736
rect 9696 8672 9702 8736
rect 9386 8671 9702 8672
rect 17827 8736 18143 8737
rect 17827 8672 17833 8736
rect 17897 8672 17913 8736
rect 17977 8672 17993 8736
rect 18057 8672 18073 8736
rect 18137 8672 18143 8736
rect 17827 8671 18143 8672
rect 26268 8736 26584 8737
rect 26268 8672 26274 8736
rect 26338 8672 26354 8736
rect 26418 8672 26434 8736
rect 26498 8672 26514 8736
rect 26578 8672 26584 8736
rect 26268 8671 26584 8672
rect 34709 8736 35025 8737
rect 34709 8672 34715 8736
rect 34779 8672 34795 8736
rect 34859 8672 34875 8736
rect 34939 8672 34955 8736
rect 35019 8672 35025 8736
rect 34709 8671 35025 8672
rect 5166 8192 5482 8193
rect 5166 8128 5172 8192
rect 5236 8128 5252 8192
rect 5316 8128 5332 8192
rect 5396 8128 5412 8192
rect 5476 8128 5482 8192
rect 5166 8127 5482 8128
rect 13607 8192 13923 8193
rect 13607 8128 13613 8192
rect 13677 8128 13693 8192
rect 13757 8128 13773 8192
rect 13837 8128 13853 8192
rect 13917 8128 13923 8192
rect 13607 8127 13923 8128
rect 22048 8192 22364 8193
rect 22048 8128 22054 8192
rect 22118 8128 22134 8192
rect 22198 8128 22214 8192
rect 22278 8128 22294 8192
rect 22358 8128 22364 8192
rect 22048 8127 22364 8128
rect 30489 8192 30805 8193
rect 30489 8128 30495 8192
rect 30559 8128 30575 8192
rect 30639 8128 30655 8192
rect 30719 8128 30735 8192
rect 30799 8128 30805 8192
rect 30489 8127 30805 8128
rect 9386 7648 9702 7649
rect 9386 7584 9392 7648
rect 9456 7584 9472 7648
rect 9536 7584 9552 7648
rect 9616 7584 9632 7648
rect 9696 7584 9702 7648
rect 9386 7583 9702 7584
rect 17827 7648 18143 7649
rect 17827 7584 17833 7648
rect 17897 7584 17913 7648
rect 17977 7584 17993 7648
rect 18057 7584 18073 7648
rect 18137 7584 18143 7648
rect 17827 7583 18143 7584
rect 26268 7648 26584 7649
rect 26268 7584 26274 7648
rect 26338 7584 26354 7648
rect 26418 7584 26434 7648
rect 26498 7584 26514 7648
rect 26578 7584 26584 7648
rect 26268 7583 26584 7584
rect 34709 7648 35025 7649
rect 34709 7584 34715 7648
rect 34779 7584 34795 7648
rect 34859 7584 34875 7648
rect 34939 7584 34955 7648
rect 35019 7584 35025 7648
rect 34709 7583 35025 7584
rect 5166 7104 5482 7105
rect 5166 7040 5172 7104
rect 5236 7040 5252 7104
rect 5316 7040 5332 7104
rect 5396 7040 5412 7104
rect 5476 7040 5482 7104
rect 5166 7039 5482 7040
rect 13607 7104 13923 7105
rect 13607 7040 13613 7104
rect 13677 7040 13693 7104
rect 13757 7040 13773 7104
rect 13837 7040 13853 7104
rect 13917 7040 13923 7104
rect 13607 7039 13923 7040
rect 22048 7104 22364 7105
rect 22048 7040 22054 7104
rect 22118 7040 22134 7104
rect 22198 7040 22214 7104
rect 22278 7040 22294 7104
rect 22358 7040 22364 7104
rect 22048 7039 22364 7040
rect 30489 7104 30805 7105
rect 30489 7040 30495 7104
rect 30559 7040 30575 7104
rect 30639 7040 30655 7104
rect 30719 7040 30735 7104
rect 30799 7040 30805 7104
rect 30489 7039 30805 7040
rect 0 6898 800 6988
rect 1393 6898 1459 6901
rect 0 6896 1459 6898
rect 0 6840 1398 6896
rect 1454 6840 1459 6896
rect 0 6838 1459 6840
rect 0 6748 800 6838
rect 1393 6835 1459 6838
rect 9386 6560 9702 6561
rect 9386 6496 9392 6560
rect 9456 6496 9472 6560
rect 9536 6496 9552 6560
rect 9616 6496 9632 6560
rect 9696 6496 9702 6560
rect 9386 6495 9702 6496
rect 17827 6560 18143 6561
rect 17827 6496 17833 6560
rect 17897 6496 17913 6560
rect 17977 6496 17993 6560
rect 18057 6496 18073 6560
rect 18137 6496 18143 6560
rect 17827 6495 18143 6496
rect 26268 6560 26584 6561
rect 26268 6496 26274 6560
rect 26338 6496 26354 6560
rect 26418 6496 26434 6560
rect 26498 6496 26514 6560
rect 26578 6496 26584 6560
rect 26268 6495 26584 6496
rect 34709 6560 35025 6561
rect 34709 6496 34715 6560
rect 34779 6496 34795 6560
rect 34859 6496 34875 6560
rect 34939 6496 34955 6560
rect 35019 6496 35025 6560
rect 34709 6495 35025 6496
rect 5166 6016 5482 6017
rect 5166 5952 5172 6016
rect 5236 5952 5252 6016
rect 5316 5952 5332 6016
rect 5396 5952 5412 6016
rect 5476 5952 5482 6016
rect 5166 5951 5482 5952
rect 13607 6016 13923 6017
rect 13607 5952 13613 6016
rect 13677 5952 13693 6016
rect 13757 5952 13773 6016
rect 13837 5952 13853 6016
rect 13917 5952 13923 6016
rect 13607 5951 13923 5952
rect 22048 6016 22364 6017
rect 22048 5952 22054 6016
rect 22118 5952 22134 6016
rect 22198 5952 22214 6016
rect 22278 5952 22294 6016
rect 22358 5952 22364 6016
rect 22048 5951 22364 5952
rect 30489 6016 30805 6017
rect 30489 5952 30495 6016
rect 30559 5952 30575 6016
rect 30639 5952 30655 6016
rect 30719 5952 30735 6016
rect 30799 5952 30805 6016
rect 30489 5951 30805 5952
rect 34513 5674 34579 5677
rect 34513 5672 35220 5674
rect 34513 5616 34518 5672
rect 34574 5628 35220 5672
rect 34574 5616 36000 5628
rect 34513 5614 36000 5616
rect 34513 5611 34579 5614
rect 35160 5478 36000 5614
rect 9386 5472 9702 5473
rect 9386 5408 9392 5472
rect 9456 5408 9472 5472
rect 9536 5408 9552 5472
rect 9616 5408 9632 5472
rect 9696 5408 9702 5472
rect 9386 5407 9702 5408
rect 17827 5472 18143 5473
rect 17827 5408 17833 5472
rect 17897 5408 17913 5472
rect 17977 5408 17993 5472
rect 18057 5408 18073 5472
rect 18137 5408 18143 5472
rect 17827 5407 18143 5408
rect 26268 5472 26584 5473
rect 26268 5408 26274 5472
rect 26338 5408 26354 5472
rect 26418 5408 26434 5472
rect 26498 5408 26514 5472
rect 26578 5408 26584 5472
rect 26268 5407 26584 5408
rect 34709 5472 35025 5473
rect 34709 5408 34715 5472
rect 34779 5408 34795 5472
rect 34859 5408 34875 5472
rect 34939 5408 34955 5472
rect 35019 5408 35025 5472
rect 34709 5407 35025 5408
rect 35200 5388 36000 5478
rect 5166 4928 5482 4929
rect 5166 4864 5172 4928
rect 5236 4864 5252 4928
rect 5316 4864 5332 4928
rect 5396 4864 5412 4928
rect 5476 4864 5482 4928
rect 5166 4863 5482 4864
rect 13607 4928 13923 4929
rect 13607 4864 13613 4928
rect 13677 4864 13693 4928
rect 13757 4864 13773 4928
rect 13837 4864 13853 4928
rect 13917 4864 13923 4928
rect 13607 4863 13923 4864
rect 22048 4928 22364 4929
rect 22048 4864 22054 4928
rect 22118 4864 22134 4928
rect 22198 4864 22214 4928
rect 22278 4864 22294 4928
rect 22358 4864 22364 4928
rect 22048 4863 22364 4864
rect 30489 4928 30805 4929
rect 30489 4864 30495 4928
rect 30559 4864 30575 4928
rect 30639 4864 30655 4928
rect 30719 4864 30735 4928
rect 30799 4864 30805 4928
rect 30489 4863 30805 4864
rect 9386 4384 9702 4385
rect 9386 4320 9392 4384
rect 9456 4320 9472 4384
rect 9536 4320 9552 4384
rect 9616 4320 9632 4384
rect 9696 4320 9702 4384
rect 9386 4319 9702 4320
rect 17827 4384 18143 4385
rect 17827 4320 17833 4384
rect 17897 4320 17913 4384
rect 17977 4320 17993 4384
rect 18057 4320 18073 4384
rect 18137 4320 18143 4384
rect 17827 4319 18143 4320
rect 26268 4384 26584 4385
rect 26268 4320 26274 4384
rect 26338 4320 26354 4384
rect 26418 4320 26434 4384
rect 26498 4320 26514 4384
rect 26578 4320 26584 4384
rect 26268 4319 26584 4320
rect 34709 4384 35025 4385
rect 34709 4320 34715 4384
rect 34779 4320 34795 4384
rect 34859 4320 34875 4384
rect 34939 4320 34955 4384
rect 35019 4320 35025 4384
rect 34709 4319 35025 4320
rect 5166 3840 5482 3841
rect 5166 3776 5172 3840
rect 5236 3776 5252 3840
rect 5316 3776 5332 3840
rect 5396 3776 5412 3840
rect 5476 3776 5482 3840
rect 5166 3775 5482 3776
rect 13607 3840 13923 3841
rect 13607 3776 13613 3840
rect 13677 3776 13693 3840
rect 13757 3776 13773 3840
rect 13837 3776 13853 3840
rect 13917 3776 13923 3840
rect 13607 3775 13923 3776
rect 22048 3840 22364 3841
rect 22048 3776 22054 3840
rect 22118 3776 22134 3840
rect 22198 3776 22214 3840
rect 22278 3776 22294 3840
rect 22358 3776 22364 3840
rect 22048 3775 22364 3776
rect 30489 3840 30805 3841
rect 30489 3776 30495 3840
rect 30559 3776 30575 3840
rect 30639 3776 30655 3840
rect 30719 3776 30735 3840
rect 30799 3776 30805 3840
rect 30489 3775 30805 3776
rect 9386 3296 9702 3297
rect 9386 3232 9392 3296
rect 9456 3232 9472 3296
rect 9536 3232 9552 3296
rect 9616 3232 9632 3296
rect 9696 3232 9702 3296
rect 9386 3231 9702 3232
rect 17827 3296 18143 3297
rect 17827 3232 17833 3296
rect 17897 3232 17913 3296
rect 17977 3232 17993 3296
rect 18057 3232 18073 3296
rect 18137 3232 18143 3296
rect 17827 3231 18143 3232
rect 26268 3296 26584 3297
rect 26268 3232 26274 3296
rect 26338 3232 26354 3296
rect 26418 3232 26434 3296
rect 26498 3232 26514 3296
rect 26578 3232 26584 3296
rect 26268 3231 26584 3232
rect 34709 3296 35025 3297
rect 34709 3232 34715 3296
rect 34779 3232 34795 3296
rect 34859 3232 34875 3296
rect 34939 3232 34955 3296
rect 35019 3232 35025 3296
rect 34709 3231 35025 3232
rect 5166 2752 5482 2753
rect 5166 2688 5172 2752
rect 5236 2688 5252 2752
rect 5316 2688 5332 2752
rect 5396 2688 5412 2752
rect 5476 2688 5482 2752
rect 5166 2687 5482 2688
rect 13607 2752 13923 2753
rect 13607 2688 13613 2752
rect 13677 2688 13693 2752
rect 13757 2688 13773 2752
rect 13837 2688 13853 2752
rect 13917 2688 13923 2752
rect 13607 2687 13923 2688
rect 22048 2752 22364 2753
rect 22048 2688 22054 2752
rect 22118 2688 22134 2752
rect 22198 2688 22214 2752
rect 22278 2688 22294 2752
rect 22358 2688 22364 2752
rect 22048 2687 22364 2688
rect 30489 2752 30805 2753
rect 30489 2688 30495 2752
rect 30559 2688 30575 2752
rect 30639 2688 30655 2752
rect 30719 2688 30735 2752
rect 30799 2688 30805 2752
rect 30489 2687 30805 2688
rect 9386 2208 9702 2209
rect 9386 2144 9392 2208
rect 9456 2144 9472 2208
rect 9536 2144 9552 2208
rect 9616 2144 9632 2208
rect 9696 2144 9702 2208
rect 9386 2143 9702 2144
rect 17827 2208 18143 2209
rect 17827 2144 17833 2208
rect 17897 2144 17913 2208
rect 17977 2144 17993 2208
rect 18057 2144 18073 2208
rect 18137 2144 18143 2208
rect 17827 2143 18143 2144
rect 26268 2208 26584 2209
rect 26268 2144 26274 2208
rect 26338 2144 26354 2208
rect 26418 2144 26434 2208
rect 26498 2144 26514 2208
rect 26578 2144 26584 2208
rect 26268 2143 26584 2144
rect 34709 2208 35025 2209
rect 34709 2144 34715 2208
rect 34779 2144 34795 2208
rect 34859 2144 34875 2208
rect 34939 2144 34955 2208
rect 35019 2144 35025 2208
rect 34709 2143 35025 2144
<< via3 >>
rect 5172 39740 5236 39744
rect 5172 39684 5176 39740
rect 5176 39684 5232 39740
rect 5232 39684 5236 39740
rect 5172 39680 5236 39684
rect 5252 39740 5316 39744
rect 5252 39684 5256 39740
rect 5256 39684 5312 39740
rect 5312 39684 5316 39740
rect 5252 39680 5316 39684
rect 5332 39740 5396 39744
rect 5332 39684 5336 39740
rect 5336 39684 5392 39740
rect 5392 39684 5396 39740
rect 5332 39680 5396 39684
rect 5412 39740 5476 39744
rect 5412 39684 5416 39740
rect 5416 39684 5472 39740
rect 5472 39684 5476 39740
rect 5412 39680 5476 39684
rect 13613 39740 13677 39744
rect 13613 39684 13617 39740
rect 13617 39684 13673 39740
rect 13673 39684 13677 39740
rect 13613 39680 13677 39684
rect 13693 39740 13757 39744
rect 13693 39684 13697 39740
rect 13697 39684 13753 39740
rect 13753 39684 13757 39740
rect 13693 39680 13757 39684
rect 13773 39740 13837 39744
rect 13773 39684 13777 39740
rect 13777 39684 13833 39740
rect 13833 39684 13837 39740
rect 13773 39680 13837 39684
rect 13853 39740 13917 39744
rect 13853 39684 13857 39740
rect 13857 39684 13913 39740
rect 13913 39684 13917 39740
rect 13853 39680 13917 39684
rect 22054 39740 22118 39744
rect 22054 39684 22058 39740
rect 22058 39684 22114 39740
rect 22114 39684 22118 39740
rect 22054 39680 22118 39684
rect 22134 39740 22198 39744
rect 22134 39684 22138 39740
rect 22138 39684 22194 39740
rect 22194 39684 22198 39740
rect 22134 39680 22198 39684
rect 22214 39740 22278 39744
rect 22214 39684 22218 39740
rect 22218 39684 22274 39740
rect 22274 39684 22278 39740
rect 22214 39680 22278 39684
rect 22294 39740 22358 39744
rect 22294 39684 22298 39740
rect 22298 39684 22354 39740
rect 22354 39684 22358 39740
rect 22294 39680 22358 39684
rect 30495 39740 30559 39744
rect 30495 39684 30499 39740
rect 30499 39684 30555 39740
rect 30555 39684 30559 39740
rect 30495 39680 30559 39684
rect 30575 39740 30639 39744
rect 30575 39684 30579 39740
rect 30579 39684 30635 39740
rect 30635 39684 30639 39740
rect 30575 39680 30639 39684
rect 30655 39740 30719 39744
rect 30655 39684 30659 39740
rect 30659 39684 30715 39740
rect 30715 39684 30719 39740
rect 30655 39680 30719 39684
rect 30735 39740 30799 39744
rect 30735 39684 30739 39740
rect 30739 39684 30795 39740
rect 30795 39684 30799 39740
rect 30735 39680 30799 39684
rect 9392 39196 9456 39200
rect 9392 39140 9396 39196
rect 9396 39140 9452 39196
rect 9452 39140 9456 39196
rect 9392 39136 9456 39140
rect 9472 39196 9536 39200
rect 9472 39140 9476 39196
rect 9476 39140 9532 39196
rect 9532 39140 9536 39196
rect 9472 39136 9536 39140
rect 9552 39196 9616 39200
rect 9552 39140 9556 39196
rect 9556 39140 9612 39196
rect 9612 39140 9616 39196
rect 9552 39136 9616 39140
rect 9632 39196 9696 39200
rect 9632 39140 9636 39196
rect 9636 39140 9692 39196
rect 9692 39140 9696 39196
rect 9632 39136 9696 39140
rect 17833 39196 17897 39200
rect 17833 39140 17837 39196
rect 17837 39140 17893 39196
rect 17893 39140 17897 39196
rect 17833 39136 17897 39140
rect 17913 39196 17977 39200
rect 17913 39140 17917 39196
rect 17917 39140 17973 39196
rect 17973 39140 17977 39196
rect 17913 39136 17977 39140
rect 17993 39196 18057 39200
rect 17993 39140 17997 39196
rect 17997 39140 18053 39196
rect 18053 39140 18057 39196
rect 17993 39136 18057 39140
rect 18073 39196 18137 39200
rect 18073 39140 18077 39196
rect 18077 39140 18133 39196
rect 18133 39140 18137 39196
rect 18073 39136 18137 39140
rect 26274 39196 26338 39200
rect 26274 39140 26278 39196
rect 26278 39140 26334 39196
rect 26334 39140 26338 39196
rect 26274 39136 26338 39140
rect 26354 39196 26418 39200
rect 26354 39140 26358 39196
rect 26358 39140 26414 39196
rect 26414 39140 26418 39196
rect 26354 39136 26418 39140
rect 26434 39196 26498 39200
rect 26434 39140 26438 39196
rect 26438 39140 26494 39196
rect 26494 39140 26498 39196
rect 26434 39136 26498 39140
rect 26514 39196 26578 39200
rect 26514 39140 26518 39196
rect 26518 39140 26574 39196
rect 26574 39140 26578 39196
rect 26514 39136 26578 39140
rect 34715 39196 34779 39200
rect 34715 39140 34719 39196
rect 34719 39140 34775 39196
rect 34775 39140 34779 39196
rect 34715 39136 34779 39140
rect 34795 39196 34859 39200
rect 34795 39140 34799 39196
rect 34799 39140 34855 39196
rect 34855 39140 34859 39196
rect 34795 39136 34859 39140
rect 34875 39196 34939 39200
rect 34875 39140 34879 39196
rect 34879 39140 34935 39196
rect 34935 39140 34939 39196
rect 34875 39136 34939 39140
rect 34955 39196 35019 39200
rect 34955 39140 34959 39196
rect 34959 39140 35015 39196
rect 35015 39140 35019 39196
rect 34955 39136 35019 39140
rect 5172 38652 5236 38656
rect 5172 38596 5176 38652
rect 5176 38596 5232 38652
rect 5232 38596 5236 38652
rect 5172 38592 5236 38596
rect 5252 38652 5316 38656
rect 5252 38596 5256 38652
rect 5256 38596 5312 38652
rect 5312 38596 5316 38652
rect 5252 38592 5316 38596
rect 5332 38652 5396 38656
rect 5332 38596 5336 38652
rect 5336 38596 5392 38652
rect 5392 38596 5396 38652
rect 5332 38592 5396 38596
rect 5412 38652 5476 38656
rect 5412 38596 5416 38652
rect 5416 38596 5472 38652
rect 5472 38596 5476 38652
rect 5412 38592 5476 38596
rect 13613 38652 13677 38656
rect 13613 38596 13617 38652
rect 13617 38596 13673 38652
rect 13673 38596 13677 38652
rect 13613 38592 13677 38596
rect 13693 38652 13757 38656
rect 13693 38596 13697 38652
rect 13697 38596 13753 38652
rect 13753 38596 13757 38652
rect 13693 38592 13757 38596
rect 13773 38652 13837 38656
rect 13773 38596 13777 38652
rect 13777 38596 13833 38652
rect 13833 38596 13837 38652
rect 13773 38592 13837 38596
rect 13853 38652 13917 38656
rect 13853 38596 13857 38652
rect 13857 38596 13913 38652
rect 13913 38596 13917 38652
rect 13853 38592 13917 38596
rect 22054 38652 22118 38656
rect 22054 38596 22058 38652
rect 22058 38596 22114 38652
rect 22114 38596 22118 38652
rect 22054 38592 22118 38596
rect 22134 38652 22198 38656
rect 22134 38596 22138 38652
rect 22138 38596 22194 38652
rect 22194 38596 22198 38652
rect 22134 38592 22198 38596
rect 22214 38652 22278 38656
rect 22214 38596 22218 38652
rect 22218 38596 22274 38652
rect 22274 38596 22278 38652
rect 22214 38592 22278 38596
rect 22294 38652 22358 38656
rect 22294 38596 22298 38652
rect 22298 38596 22354 38652
rect 22354 38596 22358 38652
rect 22294 38592 22358 38596
rect 30495 38652 30559 38656
rect 30495 38596 30499 38652
rect 30499 38596 30555 38652
rect 30555 38596 30559 38652
rect 30495 38592 30559 38596
rect 30575 38652 30639 38656
rect 30575 38596 30579 38652
rect 30579 38596 30635 38652
rect 30635 38596 30639 38652
rect 30575 38592 30639 38596
rect 30655 38652 30719 38656
rect 30655 38596 30659 38652
rect 30659 38596 30715 38652
rect 30715 38596 30719 38652
rect 30655 38592 30719 38596
rect 30735 38652 30799 38656
rect 30735 38596 30739 38652
rect 30739 38596 30795 38652
rect 30795 38596 30799 38652
rect 30735 38592 30799 38596
rect 9392 38108 9456 38112
rect 9392 38052 9396 38108
rect 9396 38052 9452 38108
rect 9452 38052 9456 38108
rect 9392 38048 9456 38052
rect 9472 38108 9536 38112
rect 9472 38052 9476 38108
rect 9476 38052 9532 38108
rect 9532 38052 9536 38108
rect 9472 38048 9536 38052
rect 9552 38108 9616 38112
rect 9552 38052 9556 38108
rect 9556 38052 9612 38108
rect 9612 38052 9616 38108
rect 9552 38048 9616 38052
rect 9632 38108 9696 38112
rect 9632 38052 9636 38108
rect 9636 38052 9692 38108
rect 9692 38052 9696 38108
rect 9632 38048 9696 38052
rect 17833 38108 17897 38112
rect 17833 38052 17837 38108
rect 17837 38052 17893 38108
rect 17893 38052 17897 38108
rect 17833 38048 17897 38052
rect 17913 38108 17977 38112
rect 17913 38052 17917 38108
rect 17917 38052 17973 38108
rect 17973 38052 17977 38108
rect 17913 38048 17977 38052
rect 17993 38108 18057 38112
rect 17993 38052 17997 38108
rect 17997 38052 18053 38108
rect 18053 38052 18057 38108
rect 17993 38048 18057 38052
rect 18073 38108 18137 38112
rect 18073 38052 18077 38108
rect 18077 38052 18133 38108
rect 18133 38052 18137 38108
rect 18073 38048 18137 38052
rect 26274 38108 26338 38112
rect 26274 38052 26278 38108
rect 26278 38052 26334 38108
rect 26334 38052 26338 38108
rect 26274 38048 26338 38052
rect 26354 38108 26418 38112
rect 26354 38052 26358 38108
rect 26358 38052 26414 38108
rect 26414 38052 26418 38108
rect 26354 38048 26418 38052
rect 26434 38108 26498 38112
rect 26434 38052 26438 38108
rect 26438 38052 26494 38108
rect 26494 38052 26498 38108
rect 26434 38048 26498 38052
rect 26514 38108 26578 38112
rect 26514 38052 26518 38108
rect 26518 38052 26574 38108
rect 26574 38052 26578 38108
rect 26514 38048 26578 38052
rect 34715 38108 34779 38112
rect 34715 38052 34719 38108
rect 34719 38052 34775 38108
rect 34775 38052 34779 38108
rect 34715 38048 34779 38052
rect 34795 38108 34859 38112
rect 34795 38052 34799 38108
rect 34799 38052 34855 38108
rect 34855 38052 34859 38108
rect 34795 38048 34859 38052
rect 34875 38108 34939 38112
rect 34875 38052 34879 38108
rect 34879 38052 34935 38108
rect 34935 38052 34939 38108
rect 34875 38048 34939 38052
rect 34955 38108 35019 38112
rect 34955 38052 34959 38108
rect 34959 38052 35015 38108
rect 35015 38052 35019 38108
rect 34955 38048 35019 38052
rect 5172 37564 5236 37568
rect 5172 37508 5176 37564
rect 5176 37508 5232 37564
rect 5232 37508 5236 37564
rect 5172 37504 5236 37508
rect 5252 37564 5316 37568
rect 5252 37508 5256 37564
rect 5256 37508 5312 37564
rect 5312 37508 5316 37564
rect 5252 37504 5316 37508
rect 5332 37564 5396 37568
rect 5332 37508 5336 37564
rect 5336 37508 5392 37564
rect 5392 37508 5396 37564
rect 5332 37504 5396 37508
rect 5412 37564 5476 37568
rect 5412 37508 5416 37564
rect 5416 37508 5472 37564
rect 5472 37508 5476 37564
rect 5412 37504 5476 37508
rect 13613 37564 13677 37568
rect 13613 37508 13617 37564
rect 13617 37508 13673 37564
rect 13673 37508 13677 37564
rect 13613 37504 13677 37508
rect 13693 37564 13757 37568
rect 13693 37508 13697 37564
rect 13697 37508 13753 37564
rect 13753 37508 13757 37564
rect 13693 37504 13757 37508
rect 13773 37564 13837 37568
rect 13773 37508 13777 37564
rect 13777 37508 13833 37564
rect 13833 37508 13837 37564
rect 13773 37504 13837 37508
rect 13853 37564 13917 37568
rect 13853 37508 13857 37564
rect 13857 37508 13913 37564
rect 13913 37508 13917 37564
rect 13853 37504 13917 37508
rect 22054 37564 22118 37568
rect 22054 37508 22058 37564
rect 22058 37508 22114 37564
rect 22114 37508 22118 37564
rect 22054 37504 22118 37508
rect 22134 37564 22198 37568
rect 22134 37508 22138 37564
rect 22138 37508 22194 37564
rect 22194 37508 22198 37564
rect 22134 37504 22198 37508
rect 22214 37564 22278 37568
rect 22214 37508 22218 37564
rect 22218 37508 22274 37564
rect 22274 37508 22278 37564
rect 22214 37504 22278 37508
rect 22294 37564 22358 37568
rect 22294 37508 22298 37564
rect 22298 37508 22354 37564
rect 22354 37508 22358 37564
rect 22294 37504 22358 37508
rect 30495 37564 30559 37568
rect 30495 37508 30499 37564
rect 30499 37508 30555 37564
rect 30555 37508 30559 37564
rect 30495 37504 30559 37508
rect 30575 37564 30639 37568
rect 30575 37508 30579 37564
rect 30579 37508 30635 37564
rect 30635 37508 30639 37564
rect 30575 37504 30639 37508
rect 30655 37564 30719 37568
rect 30655 37508 30659 37564
rect 30659 37508 30715 37564
rect 30715 37508 30719 37564
rect 30655 37504 30719 37508
rect 30735 37564 30799 37568
rect 30735 37508 30739 37564
rect 30739 37508 30795 37564
rect 30795 37508 30799 37564
rect 30735 37504 30799 37508
rect 9392 37020 9456 37024
rect 9392 36964 9396 37020
rect 9396 36964 9452 37020
rect 9452 36964 9456 37020
rect 9392 36960 9456 36964
rect 9472 37020 9536 37024
rect 9472 36964 9476 37020
rect 9476 36964 9532 37020
rect 9532 36964 9536 37020
rect 9472 36960 9536 36964
rect 9552 37020 9616 37024
rect 9552 36964 9556 37020
rect 9556 36964 9612 37020
rect 9612 36964 9616 37020
rect 9552 36960 9616 36964
rect 9632 37020 9696 37024
rect 9632 36964 9636 37020
rect 9636 36964 9692 37020
rect 9692 36964 9696 37020
rect 9632 36960 9696 36964
rect 17833 37020 17897 37024
rect 17833 36964 17837 37020
rect 17837 36964 17893 37020
rect 17893 36964 17897 37020
rect 17833 36960 17897 36964
rect 17913 37020 17977 37024
rect 17913 36964 17917 37020
rect 17917 36964 17973 37020
rect 17973 36964 17977 37020
rect 17913 36960 17977 36964
rect 17993 37020 18057 37024
rect 17993 36964 17997 37020
rect 17997 36964 18053 37020
rect 18053 36964 18057 37020
rect 17993 36960 18057 36964
rect 18073 37020 18137 37024
rect 18073 36964 18077 37020
rect 18077 36964 18133 37020
rect 18133 36964 18137 37020
rect 18073 36960 18137 36964
rect 26274 37020 26338 37024
rect 26274 36964 26278 37020
rect 26278 36964 26334 37020
rect 26334 36964 26338 37020
rect 26274 36960 26338 36964
rect 26354 37020 26418 37024
rect 26354 36964 26358 37020
rect 26358 36964 26414 37020
rect 26414 36964 26418 37020
rect 26354 36960 26418 36964
rect 26434 37020 26498 37024
rect 26434 36964 26438 37020
rect 26438 36964 26494 37020
rect 26494 36964 26498 37020
rect 26434 36960 26498 36964
rect 26514 37020 26578 37024
rect 26514 36964 26518 37020
rect 26518 36964 26574 37020
rect 26574 36964 26578 37020
rect 26514 36960 26578 36964
rect 34715 37020 34779 37024
rect 34715 36964 34719 37020
rect 34719 36964 34775 37020
rect 34775 36964 34779 37020
rect 34715 36960 34779 36964
rect 34795 37020 34859 37024
rect 34795 36964 34799 37020
rect 34799 36964 34855 37020
rect 34855 36964 34859 37020
rect 34795 36960 34859 36964
rect 34875 37020 34939 37024
rect 34875 36964 34879 37020
rect 34879 36964 34935 37020
rect 34935 36964 34939 37020
rect 34875 36960 34939 36964
rect 34955 37020 35019 37024
rect 34955 36964 34959 37020
rect 34959 36964 35015 37020
rect 35015 36964 35019 37020
rect 34955 36960 35019 36964
rect 5172 36476 5236 36480
rect 5172 36420 5176 36476
rect 5176 36420 5232 36476
rect 5232 36420 5236 36476
rect 5172 36416 5236 36420
rect 5252 36476 5316 36480
rect 5252 36420 5256 36476
rect 5256 36420 5312 36476
rect 5312 36420 5316 36476
rect 5252 36416 5316 36420
rect 5332 36476 5396 36480
rect 5332 36420 5336 36476
rect 5336 36420 5392 36476
rect 5392 36420 5396 36476
rect 5332 36416 5396 36420
rect 5412 36476 5476 36480
rect 5412 36420 5416 36476
rect 5416 36420 5472 36476
rect 5472 36420 5476 36476
rect 5412 36416 5476 36420
rect 13613 36476 13677 36480
rect 13613 36420 13617 36476
rect 13617 36420 13673 36476
rect 13673 36420 13677 36476
rect 13613 36416 13677 36420
rect 13693 36476 13757 36480
rect 13693 36420 13697 36476
rect 13697 36420 13753 36476
rect 13753 36420 13757 36476
rect 13693 36416 13757 36420
rect 13773 36476 13837 36480
rect 13773 36420 13777 36476
rect 13777 36420 13833 36476
rect 13833 36420 13837 36476
rect 13773 36416 13837 36420
rect 13853 36476 13917 36480
rect 13853 36420 13857 36476
rect 13857 36420 13913 36476
rect 13913 36420 13917 36476
rect 13853 36416 13917 36420
rect 22054 36476 22118 36480
rect 22054 36420 22058 36476
rect 22058 36420 22114 36476
rect 22114 36420 22118 36476
rect 22054 36416 22118 36420
rect 22134 36476 22198 36480
rect 22134 36420 22138 36476
rect 22138 36420 22194 36476
rect 22194 36420 22198 36476
rect 22134 36416 22198 36420
rect 22214 36476 22278 36480
rect 22214 36420 22218 36476
rect 22218 36420 22274 36476
rect 22274 36420 22278 36476
rect 22214 36416 22278 36420
rect 22294 36476 22358 36480
rect 22294 36420 22298 36476
rect 22298 36420 22354 36476
rect 22354 36420 22358 36476
rect 22294 36416 22358 36420
rect 30495 36476 30559 36480
rect 30495 36420 30499 36476
rect 30499 36420 30555 36476
rect 30555 36420 30559 36476
rect 30495 36416 30559 36420
rect 30575 36476 30639 36480
rect 30575 36420 30579 36476
rect 30579 36420 30635 36476
rect 30635 36420 30639 36476
rect 30575 36416 30639 36420
rect 30655 36476 30719 36480
rect 30655 36420 30659 36476
rect 30659 36420 30715 36476
rect 30715 36420 30719 36476
rect 30655 36416 30719 36420
rect 30735 36476 30799 36480
rect 30735 36420 30739 36476
rect 30739 36420 30795 36476
rect 30795 36420 30799 36476
rect 30735 36416 30799 36420
rect 9392 35932 9456 35936
rect 9392 35876 9396 35932
rect 9396 35876 9452 35932
rect 9452 35876 9456 35932
rect 9392 35872 9456 35876
rect 9472 35932 9536 35936
rect 9472 35876 9476 35932
rect 9476 35876 9532 35932
rect 9532 35876 9536 35932
rect 9472 35872 9536 35876
rect 9552 35932 9616 35936
rect 9552 35876 9556 35932
rect 9556 35876 9612 35932
rect 9612 35876 9616 35932
rect 9552 35872 9616 35876
rect 9632 35932 9696 35936
rect 9632 35876 9636 35932
rect 9636 35876 9692 35932
rect 9692 35876 9696 35932
rect 9632 35872 9696 35876
rect 17833 35932 17897 35936
rect 17833 35876 17837 35932
rect 17837 35876 17893 35932
rect 17893 35876 17897 35932
rect 17833 35872 17897 35876
rect 17913 35932 17977 35936
rect 17913 35876 17917 35932
rect 17917 35876 17973 35932
rect 17973 35876 17977 35932
rect 17913 35872 17977 35876
rect 17993 35932 18057 35936
rect 17993 35876 17997 35932
rect 17997 35876 18053 35932
rect 18053 35876 18057 35932
rect 17993 35872 18057 35876
rect 18073 35932 18137 35936
rect 18073 35876 18077 35932
rect 18077 35876 18133 35932
rect 18133 35876 18137 35932
rect 18073 35872 18137 35876
rect 26274 35932 26338 35936
rect 26274 35876 26278 35932
rect 26278 35876 26334 35932
rect 26334 35876 26338 35932
rect 26274 35872 26338 35876
rect 26354 35932 26418 35936
rect 26354 35876 26358 35932
rect 26358 35876 26414 35932
rect 26414 35876 26418 35932
rect 26354 35872 26418 35876
rect 26434 35932 26498 35936
rect 26434 35876 26438 35932
rect 26438 35876 26494 35932
rect 26494 35876 26498 35932
rect 26434 35872 26498 35876
rect 26514 35932 26578 35936
rect 26514 35876 26518 35932
rect 26518 35876 26574 35932
rect 26574 35876 26578 35932
rect 26514 35872 26578 35876
rect 34715 35932 34779 35936
rect 34715 35876 34719 35932
rect 34719 35876 34775 35932
rect 34775 35876 34779 35932
rect 34715 35872 34779 35876
rect 34795 35932 34859 35936
rect 34795 35876 34799 35932
rect 34799 35876 34855 35932
rect 34855 35876 34859 35932
rect 34795 35872 34859 35876
rect 34875 35932 34939 35936
rect 34875 35876 34879 35932
rect 34879 35876 34935 35932
rect 34935 35876 34939 35932
rect 34875 35872 34939 35876
rect 34955 35932 35019 35936
rect 34955 35876 34959 35932
rect 34959 35876 35015 35932
rect 35015 35876 35019 35932
rect 34955 35872 35019 35876
rect 5172 35388 5236 35392
rect 5172 35332 5176 35388
rect 5176 35332 5232 35388
rect 5232 35332 5236 35388
rect 5172 35328 5236 35332
rect 5252 35388 5316 35392
rect 5252 35332 5256 35388
rect 5256 35332 5312 35388
rect 5312 35332 5316 35388
rect 5252 35328 5316 35332
rect 5332 35388 5396 35392
rect 5332 35332 5336 35388
rect 5336 35332 5392 35388
rect 5392 35332 5396 35388
rect 5332 35328 5396 35332
rect 5412 35388 5476 35392
rect 5412 35332 5416 35388
rect 5416 35332 5472 35388
rect 5472 35332 5476 35388
rect 5412 35328 5476 35332
rect 13613 35388 13677 35392
rect 13613 35332 13617 35388
rect 13617 35332 13673 35388
rect 13673 35332 13677 35388
rect 13613 35328 13677 35332
rect 13693 35388 13757 35392
rect 13693 35332 13697 35388
rect 13697 35332 13753 35388
rect 13753 35332 13757 35388
rect 13693 35328 13757 35332
rect 13773 35388 13837 35392
rect 13773 35332 13777 35388
rect 13777 35332 13833 35388
rect 13833 35332 13837 35388
rect 13773 35328 13837 35332
rect 13853 35388 13917 35392
rect 13853 35332 13857 35388
rect 13857 35332 13913 35388
rect 13913 35332 13917 35388
rect 13853 35328 13917 35332
rect 22054 35388 22118 35392
rect 22054 35332 22058 35388
rect 22058 35332 22114 35388
rect 22114 35332 22118 35388
rect 22054 35328 22118 35332
rect 22134 35388 22198 35392
rect 22134 35332 22138 35388
rect 22138 35332 22194 35388
rect 22194 35332 22198 35388
rect 22134 35328 22198 35332
rect 22214 35388 22278 35392
rect 22214 35332 22218 35388
rect 22218 35332 22274 35388
rect 22274 35332 22278 35388
rect 22214 35328 22278 35332
rect 22294 35388 22358 35392
rect 22294 35332 22298 35388
rect 22298 35332 22354 35388
rect 22354 35332 22358 35388
rect 22294 35328 22358 35332
rect 30495 35388 30559 35392
rect 30495 35332 30499 35388
rect 30499 35332 30555 35388
rect 30555 35332 30559 35388
rect 30495 35328 30559 35332
rect 30575 35388 30639 35392
rect 30575 35332 30579 35388
rect 30579 35332 30635 35388
rect 30635 35332 30639 35388
rect 30575 35328 30639 35332
rect 30655 35388 30719 35392
rect 30655 35332 30659 35388
rect 30659 35332 30715 35388
rect 30715 35332 30719 35388
rect 30655 35328 30719 35332
rect 30735 35388 30799 35392
rect 30735 35332 30739 35388
rect 30739 35332 30795 35388
rect 30795 35332 30799 35388
rect 30735 35328 30799 35332
rect 9392 34844 9456 34848
rect 9392 34788 9396 34844
rect 9396 34788 9452 34844
rect 9452 34788 9456 34844
rect 9392 34784 9456 34788
rect 9472 34844 9536 34848
rect 9472 34788 9476 34844
rect 9476 34788 9532 34844
rect 9532 34788 9536 34844
rect 9472 34784 9536 34788
rect 9552 34844 9616 34848
rect 9552 34788 9556 34844
rect 9556 34788 9612 34844
rect 9612 34788 9616 34844
rect 9552 34784 9616 34788
rect 9632 34844 9696 34848
rect 9632 34788 9636 34844
rect 9636 34788 9692 34844
rect 9692 34788 9696 34844
rect 9632 34784 9696 34788
rect 17833 34844 17897 34848
rect 17833 34788 17837 34844
rect 17837 34788 17893 34844
rect 17893 34788 17897 34844
rect 17833 34784 17897 34788
rect 17913 34844 17977 34848
rect 17913 34788 17917 34844
rect 17917 34788 17973 34844
rect 17973 34788 17977 34844
rect 17913 34784 17977 34788
rect 17993 34844 18057 34848
rect 17993 34788 17997 34844
rect 17997 34788 18053 34844
rect 18053 34788 18057 34844
rect 17993 34784 18057 34788
rect 18073 34844 18137 34848
rect 18073 34788 18077 34844
rect 18077 34788 18133 34844
rect 18133 34788 18137 34844
rect 18073 34784 18137 34788
rect 26274 34844 26338 34848
rect 26274 34788 26278 34844
rect 26278 34788 26334 34844
rect 26334 34788 26338 34844
rect 26274 34784 26338 34788
rect 26354 34844 26418 34848
rect 26354 34788 26358 34844
rect 26358 34788 26414 34844
rect 26414 34788 26418 34844
rect 26354 34784 26418 34788
rect 26434 34844 26498 34848
rect 26434 34788 26438 34844
rect 26438 34788 26494 34844
rect 26494 34788 26498 34844
rect 26434 34784 26498 34788
rect 26514 34844 26578 34848
rect 26514 34788 26518 34844
rect 26518 34788 26574 34844
rect 26574 34788 26578 34844
rect 26514 34784 26578 34788
rect 34715 34844 34779 34848
rect 34715 34788 34719 34844
rect 34719 34788 34775 34844
rect 34775 34788 34779 34844
rect 34715 34784 34779 34788
rect 34795 34844 34859 34848
rect 34795 34788 34799 34844
rect 34799 34788 34855 34844
rect 34855 34788 34859 34844
rect 34795 34784 34859 34788
rect 34875 34844 34939 34848
rect 34875 34788 34879 34844
rect 34879 34788 34935 34844
rect 34935 34788 34939 34844
rect 34875 34784 34939 34788
rect 34955 34844 35019 34848
rect 34955 34788 34959 34844
rect 34959 34788 35015 34844
rect 35015 34788 35019 34844
rect 34955 34784 35019 34788
rect 5172 34300 5236 34304
rect 5172 34244 5176 34300
rect 5176 34244 5232 34300
rect 5232 34244 5236 34300
rect 5172 34240 5236 34244
rect 5252 34300 5316 34304
rect 5252 34244 5256 34300
rect 5256 34244 5312 34300
rect 5312 34244 5316 34300
rect 5252 34240 5316 34244
rect 5332 34300 5396 34304
rect 5332 34244 5336 34300
rect 5336 34244 5392 34300
rect 5392 34244 5396 34300
rect 5332 34240 5396 34244
rect 5412 34300 5476 34304
rect 5412 34244 5416 34300
rect 5416 34244 5472 34300
rect 5472 34244 5476 34300
rect 5412 34240 5476 34244
rect 13613 34300 13677 34304
rect 13613 34244 13617 34300
rect 13617 34244 13673 34300
rect 13673 34244 13677 34300
rect 13613 34240 13677 34244
rect 13693 34300 13757 34304
rect 13693 34244 13697 34300
rect 13697 34244 13753 34300
rect 13753 34244 13757 34300
rect 13693 34240 13757 34244
rect 13773 34300 13837 34304
rect 13773 34244 13777 34300
rect 13777 34244 13833 34300
rect 13833 34244 13837 34300
rect 13773 34240 13837 34244
rect 13853 34300 13917 34304
rect 13853 34244 13857 34300
rect 13857 34244 13913 34300
rect 13913 34244 13917 34300
rect 13853 34240 13917 34244
rect 22054 34300 22118 34304
rect 22054 34244 22058 34300
rect 22058 34244 22114 34300
rect 22114 34244 22118 34300
rect 22054 34240 22118 34244
rect 22134 34300 22198 34304
rect 22134 34244 22138 34300
rect 22138 34244 22194 34300
rect 22194 34244 22198 34300
rect 22134 34240 22198 34244
rect 22214 34300 22278 34304
rect 22214 34244 22218 34300
rect 22218 34244 22274 34300
rect 22274 34244 22278 34300
rect 22214 34240 22278 34244
rect 22294 34300 22358 34304
rect 22294 34244 22298 34300
rect 22298 34244 22354 34300
rect 22354 34244 22358 34300
rect 22294 34240 22358 34244
rect 30495 34300 30559 34304
rect 30495 34244 30499 34300
rect 30499 34244 30555 34300
rect 30555 34244 30559 34300
rect 30495 34240 30559 34244
rect 30575 34300 30639 34304
rect 30575 34244 30579 34300
rect 30579 34244 30635 34300
rect 30635 34244 30639 34300
rect 30575 34240 30639 34244
rect 30655 34300 30719 34304
rect 30655 34244 30659 34300
rect 30659 34244 30715 34300
rect 30715 34244 30719 34300
rect 30655 34240 30719 34244
rect 30735 34300 30799 34304
rect 30735 34244 30739 34300
rect 30739 34244 30795 34300
rect 30795 34244 30799 34300
rect 30735 34240 30799 34244
rect 9392 33756 9456 33760
rect 9392 33700 9396 33756
rect 9396 33700 9452 33756
rect 9452 33700 9456 33756
rect 9392 33696 9456 33700
rect 9472 33756 9536 33760
rect 9472 33700 9476 33756
rect 9476 33700 9532 33756
rect 9532 33700 9536 33756
rect 9472 33696 9536 33700
rect 9552 33756 9616 33760
rect 9552 33700 9556 33756
rect 9556 33700 9612 33756
rect 9612 33700 9616 33756
rect 9552 33696 9616 33700
rect 9632 33756 9696 33760
rect 9632 33700 9636 33756
rect 9636 33700 9692 33756
rect 9692 33700 9696 33756
rect 9632 33696 9696 33700
rect 17833 33756 17897 33760
rect 17833 33700 17837 33756
rect 17837 33700 17893 33756
rect 17893 33700 17897 33756
rect 17833 33696 17897 33700
rect 17913 33756 17977 33760
rect 17913 33700 17917 33756
rect 17917 33700 17973 33756
rect 17973 33700 17977 33756
rect 17913 33696 17977 33700
rect 17993 33756 18057 33760
rect 17993 33700 17997 33756
rect 17997 33700 18053 33756
rect 18053 33700 18057 33756
rect 17993 33696 18057 33700
rect 18073 33756 18137 33760
rect 18073 33700 18077 33756
rect 18077 33700 18133 33756
rect 18133 33700 18137 33756
rect 18073 33696 18137 33700
rect 26274 33756 26338 33760
rect 26274 33700 26278 33756
rect 26278 33700 26334 33756
rect 26334 33700 26338 33756
rect 26274 33696 26338 33700
rect 26354 33756 26418 33760
rect 26354 33700 26358 33756
rect 26358 33700 26414 33756
rect 26414 33700 26418 33756
rect 26354 33696 26418 33700
rect 26434 33756 26498 33760
rect 26434 33700 26438 33756
rect 26438 33700 26494 33756
rect 26494 33700 26498 33756
rect 26434 33696 26498 33700
rect 26514 33756 26578 33760
rect 26514 33700 26518 33756
rect 26518 33700 26574 33756
rect 26574 33700 26578 33756
rect 26514 33696 26578 33700
rect 34715 33756 34779 33760
rect 34715 33700 34719 33756
rect 34719 33700 34775 33756
rect 34775 33700 34779 33756
rect 34715 33696 34779 33700
rect 34795 33756 34859 33760
rect 34795 33700 34799 33756
rect 34799 33700 34855 33756
rect 34855 33700 34859 33756
rect 34795 33696 34859 33700
rect 34875 33756 34939 33760
rect 34875 33700 34879 33756
rect 34879 33700 34935 33756
rect 34935 33700 34939 33756
rect 34875 33696 34939 33700
rect 34955 33756 35019 33760
rect 34955 33700 34959 33756
rect 34959 33700 35015 33756
rect 35015 33700 35019 33756
rect 34955 33696 35019 33700
rect 5172 33212 5236 33216
rect 5172 33156 5176 33212
rect 5176 33156 5232 33212
rect 5232 33156 5236 33212
rect 5172 33152 5236 33156
rect 5252 33212 5316 33216
rect 5252 33156 5256 33212
rect 5256 33156 5312 33212
rect 5312 33156 5316 33212
rect 5252 33152 5316 33156
rect 5332 33212 5396 33216
rect 5332 33156 5336 33212
rect 5336 33156 5392 33212
rect 5392 33156 5396 33212
rect 5332 33152 5396 33156
rect 5412 33212 5476 33216
rect 5412 33156 5416 33212
rect 5416 33156 5472 33212
rect 5472 33156 5476 33212
rect 5412 33152 5476 33156
rect 13613 33212 13677 33216
rect 13613 33156 13617 33212
rect 13617 33156 13673 33212
rect 13673 33156 13677 33212
rect 13613 33152 13677 33156
rect 13693 33212 13757 33216
rect 13693 33156 13697 33212
rect 13697 33156 13753 33212
rect 13753 33156 13757 33212
rect 13693 33152 13757 33156
rect 13773 33212 13837 33216
rect 13773 33156 13777 33212
rect 13777 33156 13833 33212
rect 13833 33156 13837 33212
rect 13773 33152 13837 33156
rect 13853 33212 13917 33216
rect 13853 33156 13857 33212
rect 13857 33156 13913 33212
rect 13913 33156 13917 33212
rect 13853 33152 13917 33156
rect 22054 33212 22118 33216
rect 22054 33156 22058 33212
rect 22058 33156 22114 33212
rect 22114 33156 22118 33212
rect 22054 33152 22118 33156
rect 22134 33212 22198 33216
rect 22134 33156 22138 33212
rect 22138 33156 22194 33212
rect 22194 33156 22198 33212
rect 22134 33152 22198 33156
rect 22214 33212 22278 33216
rect 22214 33156 22218 33212
rect 22218 33156 22274 33212
rect 22274 33156 22278 33212
rect 22214 33152 22278 33156
rect 22294 33212 22358 33216
rect 22294 33156 22298 33212
rect 22298 33156 22354 33212
rect 22354 33156 22358 33212
rect 22294 33152 22358 33156
rect 30495 33212 30559 33216
rect 30495 33156 30499 33212
rect 30499 33156 30555 33212
rect 30555 33156 30559 33212
rect 30495 33152 30559 33156
rect 30575 33212 30639 33216
rect 30575 33156 30579 33212
rect 30579 33156 30635 33212
rect 30635 33156 30639 33212
rect 30575 33152 30639 33156
rect 30655 33212 30719 33216
rect 30655 33156 30659 33212
rect 30659 33156 30715 33212
rect 30715 33156 30719 33212
rect 30655 33152 30719 33156
rect 30735 33212 30799 33216
rect 30735 33156 30739 33212
rect 30739 33156 30795 33212
rect 30795 33156 30799 33212
rect 30735 33152 30799 33156
rect 9392 32668 9456 32672
rect 9392 32612 9396 32668
rect 9396 32612 9452 32668
rect 9452 32612 9456 32668
rect 9392 32608 9456 32612
rect 9472 32668 9536 32672
rect 9472 32612 9476 32668
rect 9476 32612 9532 32668
rect 9532 32612 9536 32668
rect 9472 32608 9536 32612
rect 9552 32668 9616 32672
rect 9552 32612 9556 32668
rect 9556 32612 9612 32668
rect 9612 32612 9616 32668
rect 9552 32608 9616 32612
rect 9632 32668 9696 32672
rect 9632 32612 9636 32668
rect 9636 32612 9692 32668
rect 9692 32612 9696 32668
rect 9632 32608 9696 32612
rect 17833 32668 17897 32672
rect 17833 32612 17837 32668
rect 17837 32612 17893 32668
rect 17893 32612 17897 32668
rect 17833 32608 17897 32612
rect 17913 32668 17977 32672
rect 17913 32612 17917 32668
rect 17917 32612 17973 32668
rect 17973 32612 17977 32668
rect 17913 32608 17977 32612
rect 17993 32668 18057 32672
rect 17993 32612 17997 32668
rect 17997 32612 18053 32668
rect 18053 32612 18057 32668
rect 17993 32608 18057 32612
rect 18073 32668 18137 32672
rect 18073 32612 18077 32668
rect 18077 32612 18133 32668
rect 18133 32612 18137 32668
rect 18073 32608 18137 32612
rect 26274 32668 26338 32672
rect 26274 32612 26278 32668
rect 26278 32612 26334 32668
rect 26334 32612 26338 32668
rect 26274 32608 26338 32612
rect 26354 32668 26418 32672
rect 26354 32612 26358 32668
rect 26358 32612 26414 32668
rect 26414 32612 26418 32668
rect 26354 32608 26418 32612
rect 26434 32668 26498 32672
rect 26434 32612 26438 32668
rect 26438 32612 26494 32668
rect 26494 32612 26498 32668
rect 26434 32608 26498 32612
rect 26514 32668 26578 32672
rect 26514 32612 26518 32668
rect 26518 32612 26574 32668
rect 26574 32612 26578 32668
rect 26514 32608 26578 32612
rect 34715 32668 34779 32672
rect 34715 32612 34719 32668
rect 34719 32612 34775 32668
rect 34775 32612 34779 32668
rect 34715 32608 34779 32612
rect 34795 32668 34859 32672
rect 34795 32612 34799 32668
rect 34799 32612 34855 32668
rect 34855 32612 34859 32668
rect 34795 32608 34859 32612
rect 34875 32668 34939 32672
rect 34875 32612 34879 32668
rect 34879 32612 34935 32668
rect 34935 32612 34939 32668
rect 34875 32608 34939 32612
rect 34955 32668 35019 32672
rect 34955 32612 34959 32668
rect 34959 32612 35015 32668
rect 35015 32612 35019 32668
rect 34955 32608 35019 32612
rect 5172 32124 5236 32128
rect 5172 32068 5176 32124
rect 5176 32068 5232 32124
rect 5232 32068 5236 32124
rect 5172 32064 5236 32068
rect 5252 32124 5316 32128
rect 5252 32068 5256 32124
rect 5256 32068 5312 32124
rect 5312 32068 5316 32124
rect 5252 32064 5316 32068
rect 5332 32124 5396 32128
rect 5332 32068 5336 32124
rect 5336 32068 5392 32124
rect 5392 32068 5396 32124
rect 5332 32064 5396 32068
rect 5412 32124 5476 32128
rect 5412 32068 5416 32124
rect 5416 32068 5472 32124
rect 5472 32068 5476 32124
rect 5412 32064 5476 32068
rect 13613 32124 13677 32128
rect 13613 32068 13617 32124
rect 13617 32068 13673 32124
rect 13673 32068 13677 32124
rect 13613 32064 13677 32068
rect 13693 32124 13757 32128
rect 13693 32068 13697 32124
rect 13697 32068 13753 32124
rect 13753 32068 13757 32124
rect 13693 32064 13757 32068
rect 13773 32124 13837 32128
rect 13773 32068 13777 32124
rect 13777 32068 13833 32124
rect 13833 32068 13837 32124
rect 13773 32064 13837 32068
rect 13853 32124 13917 32128
rect 13853 32068 13857 32124
rect 13857 32068 13913 32124
rect 13913 32068 13917 32124
rect 13853 32064 13917 32068
rect 22054 32124 22118 32128
rect 22054 32068 22058 32124
rect 22058 32068 22114 32124
rect 22114 32068 22118 32124
rect 22054 32064 22118 32068
rect 22134 32124 22198 32128
rect 22134 32068 22138 32124
rect 22138 32068 22194 32124
rect 22194 32068 22198 32124
rect 22134 32064 22198 32068
rect 22214 32124 22278 32128
rect 22214 32068 22218 32124
rect 22218 32068 22274 32124
rect 22274 32068 22278 32124
rect 22214 32064 22278 32068
rect 22294 32124 22358 32128
rect 22294 32068 22298 32124
rect 22298 32068 22354 32124
rect 22354 32068 22358 32124
rect 22294 32064 22358 32068
rect 30495 32124 30559 32128
rect 30495 32068 30499 32124
rect 30499 32068 30555 32124
rect 30555 32068 30559 32124
rect 30495 32064 30559 32068
rect 30575 32124 30639 32128
rect 30575 32068 30579 32124
rect 30579 32068 30635 32124
rect 30635 32068 30639 32124
rect 30575 32064 30639 32068
rect 30655 32124 30719 32128
rect 30655 32068 30659 32124
rect 30659 32068 30715 32124
rect 30715 32068 30719 32124
rect 30655 32064 30719 32068
rect 30735 32124 30799 32128
rect 30735 32068 30739 32124
rect 30739 32068 30795 32124
rect 30795 32068 30799 32124
rect 30735 32064 30799 32068
rect 9392 31580 9456 31584
rect 9392 31524 9396 31580
rect 9396 31524 9452 31580
rect 9452 31524 9456 31580
rect 9392 31520 9456 31524
rect 9472 31580 9536 31584
rect 9472 31524 9476 31580
rect 9476 31524 9532 31580
rect 9532 31524 9536 31580
rect 9472 31520 9536 31524
rect 9552 31580 9616 31584
rect 9552 31524 9556 31580
rect 9556 31524 9612 31580
rect 9612 31524 9616 31580
rect 9552 31520 9616 31524
rect 9632 31580 9696 31584
rect 9632 31524 9636 31580
rect 9636 31524 9692 31580
rect 9692 31524 9696 31580
rect 9632 31520 9696 31524
rect 17833 31580 17897 31584
rect 17833 31524 17837 31580
rect 17837 31524 17893 31580
rect 17893 31524 17897 31580
rect 17833 31520 17897 31524
rect 17913 31580 17977 31584
rect 17913 31524 17917 31580
rect 17917 31524 17973 31580
rect 17973 31524 17977 31580
rect 17913 31520 17977 31524
rect 17993 31580 18057 31584
rect 17993 31524 17997 31580
rect 17997 31524 18053 31580
rect 18053 31524 18057 31580
rect 17993 31520 18057 31524
rect 18073 31580 18137 31584
rect 18073 31524 18077 31580
rect 18077 31524 18133 31580
rect 18133 31524 18137 31580
rect 18073 31520 18137 31524
rect 26274 31580 26338 31584
rect 26274 31524 26278 31580
rect 26278 31524 26334 31580
rect 26334 31524 26338 31580
rect 26274 31520 26338 31524
rect 26354 31580 26418 31584
rect 26354 31524 26358 31580
rect 26358 31524 26414 31580
rect 26414 31524 26418 31580
rect 26354 31520 26418 31524
rect 26434 31580 26498 31584
rect 26434 31524 26438 31580
rect 26438 31524 26494 31580
rect 26494 31524 26498 31580
rect 26434 31520 26498 31524
rect 26514 31580 26578 31584
rect 26514 31524 26518 31580
rect 26518 31524 26574 31580
rect 26574 31524 26578 31580
rect 26514 31520 26578 31524
rect 34715 31580 34779 31584
rect 34715 31524 34719 31580
rect 34719 31524 34775 31580
rect 34775 31524 34779 31580
rect 34715 31520 34779 31524
rect 34795 31580 34859 31584
rect 34795 31524 34799 31580
rect 34799 31524 34855 31580
rect 34855 31524 34859 31580
rect 34795 31520 34859 31524
rect 34875 31580 34939 31584
rect 34875 31524 34879 31580
rect 34879 31524 34935 31580
rect 34935 31524 34939 31580
rect 34875 31520 34939 31524
rect 34955 31580 35019 31584
rect 34955 31524 34959 31580
rect 34959 31524 35015 31580
rect 35015 31524 35019 31580
rect 34955 31520 35019 31524
rect 5172 31036 5236 31040
rect 5172 30980 5176 31036
rect 5176 30980 5232 31036
rect 5232 30980 5236 31036
rect 5172 30976 5236 30980
rect 5252 31036 5316 31040
rect 5252 30980 5256 31036
rect 5256 30980 5312 31036
rect 5312 30980 5316 31036
rect 5252 30976 5316 30980
rect 5332 31036 5396 31040
rect 5332 30980 5336 31036
rect 5336 30980 5392 31036
rect 5392 30980 5396 31036
rect 5332 30976 5396 30980
rect 5412 31036 5476 31040
rect 5412 30980 5416 31036
rect 5416 30980 5472 31036
rect 5472 30980 5476 31036
rect 5412 30976 5476 30980
rect 13613 31036 13677 31040
rect 13613 30980 13617 31036
rect 13617 30980 13673 31036
rect 13673 30980 13677 31036
rect 13613 30976 13677 30980
rect 13693 31036 13757 31040
rect 13693 30980 13697 31036
rect 13697 30980 13753 31036
rect 13753 30980 13757 31036
rect 13693 30976 13757 30980
rect 13773 31036 13837 31040
rect 13773 30980 13777 31036
rect 13777 30980 13833 31036
rect 13833 30980 13837 31036
rect 13773 30976 13837 30980
rect 13853 31036 13917 31040
rect 13853 30980 13857 31036
rect 13857 30980 13913 31036
rect 13913 30980 13917 31036
rect 13853 30976 13917 30980
rect 22054 31036 22118 31040
rect 22054 30980 22058 31036
rect 22058 30980 22114 31036
rect 22114 30980 22118 31036
rect 22054 30976 22118 30980
rect 22134 31036 22198 31040
rect 22134 30980 22138 31036
rect 22138 30980 22194 31036
rect 22194 30980 22198 31036
rect 22134 30976 22198 30980
rect 22214 31036 22278 31040
rect 22214 30980 22218 31036
rect 22218 30980 22274 31036
rect 22274 30980 22278 31036
rect 22214 30976 22278 30980
rect 22294 31036 22358 31040
rect 22294 30980 22298 31036
rect 22298 30980 22354 31036
rect 22354 30980 22358 31036
rect 22294 30976 22358 30980
rect 30495 31036 30559 31040
rect 30495 30980 30499 31036
rect 30499 30980 30555 31036
rect 30555 30980 30559 31036
rect 30495 30976 30559 30980
rect 30575 31036 30639 31040
rect 30575 30980 30579 31036
rect 30579 30980 30635 31036
rect 30635 30980 30639 31036
rect 30575 30976 30639 30980
rect 30655 31036 30719 31040
rect 30655 30980 30659 31036
rect 30659 30980 30715 31036
rect 30715 30980 30719 31036
rect 30655 30976 30719 30980
rect 30735 31036 30799 31040
rect 30735 30980 30739 31036
rect 30739 30980 30795 31036
rect 30795 30980 30799 31036
rect 30735 30976 30799 30980
rect 9392 30492 9456 30496
rect 9392 30436 9396 30492
rect 9396 30436 9452 30492
rect 9452 30436 9456 30492
rect 9392 30432 9456 30436
rect 9472 30492 9536 30496
rect 9472 30436 9476 30492
rect 9476 30436 9532 30492
rect 9532 30436 9536 30492
rect 9472 30432 9536 30436
rect 9552 30492 9616 30496
rect 9552 30436 9556 30492
rect 9556 30436 9612 30492
rect 9612 30436 9616 30492
rect 9552 30432 9616 30436
rect 9632 30492 9696 30496
rect 9632 30436 9636 30492
rect 9636 30436 9692 30492
rect 9692 30436 9696 30492
rect 9632 30432 9696 30436
rect 17833 30492 17897 30496
rect 17833 30436 17837 30492
rect 17837 30436 17893 30492
rect 17893 30436 17897 30492
rect 17833 30432 17897 30436
rect 17913 30492 17977 30496
rect 17913 30436 17917 30492
rect 17917 30436 17973 30492
rect 17973 30436 17977 30492
rect 17913 30432 17977 30436
rect 17993 30492 18057 30496
rect 17993 30436 17997 30492
rect 17997 30436 18053 30492
rect 18053 30436 18057 30492
rect 17993 30432 18057 30436
rect 18073 30492 18137 30496
rect 18073 30436 18077 30492
rect 18077 30436 18133 30492
rect 18133 30436 18137 30492
rect 18073 30432 18137 30436
rect 26274 30492 26338 30496
rect 26274 30436 26278 30492
rect 26278 30436 26334 30492
rect 26334 30436 26338 30492
rect 26274 30432 26338 30436
rect 26354 30492 26418 30496
rect 26354 30436 26358 30492
rect 26358 30436 26414 30492
rect 26414 30436 26418 30492
rect 26354 30432 26418 30436
rect 26434 30492 26498 30496
rect 26434 30436 26438 30492
rect 26438 30436 26494 30492
rect 26494 30436 26498 30492
rect 26434 30432 26498 30436
rect 26514 30492 26578 30496
rect 26514 30436 26518 30492
rect 26518 30436 26574 30492
rect 26574 30436 26578 30492
rect 26514 30432 26578 30436
rect 34715 30492 34779 30496
rect 34715 30436 34719 30492
rect 34719 30436 34775 30492
rect 34775 30436 34779 30492
rect 34715 30432 34779 30436
rect 34795 30492 34859 30496
rect 34795 30436 34799 30492
rect 34799 30436 34855 30492
rect 34855 30436 34859 30492
rect 34795 30432 34859 30436
rect 34875 30492 34939 30496
rect 34875 30436 34879 30492
rect 34879 30436 34935 30492
rect 34935 30436 34939 30492
rect 34875 30432 34939 30436
rect 34955 30492 35019 30496
rect 34955 30436 34959 30492
rect 34959 30436 35015 30492
rect 35015 30436 35019 30492
rect 34955 30432 35019 30436
rect 5172 29948 5236 29952
rect 5172 29892 5176 29948
rect 5176 29892 5232 29948
rect 5232 29892 5236 29948
rect 5172 29888 5236 29892
rect 5252 29948 5316 29952
rect 5252 29892 5256 29948
rect 5256 29892 5312 29948
rect 5312 29892 5316 29948
rect 5252 29888 5316 29892
rect 5332 29948 5396 29952
rect 5332 29892 5336 29948
rect 5336 29892 5392 29948
rect 5392 29892 5396 29948
rect 5332 29888 5396 29892
rect 5412 29948 5476 29952
rect 5412 29892 5416 29948
rect 5416 29892 5472 29948
rect 5472 29892 5476 29948
rect 5412 29888 5476 29892
rect 13613 29948 13677 29952
rect 13613 29892 13617 29948
rect 13617 29892 13673 29948
rect 13673 29892 13677 29948
rect 13613 29888 13677 29892
rect 13693 29948 13757 29952
rect 13693 29892 13697 29948
rect 13697 29892 13753 29948
rect 13753 29892 13757 29948
rect 13693 29888 13757 29892
rect 13773 29948 13837 29952
rect 13773 29892 13777 29948
rect 13777 29892 13833 29948
rect 13833 29892 13837 29948
rect 13773 29888 13837 29892
rect 13853 29948 13917 29952
rect 13853 29892 13857 29948
rect 13857 29892 13913 29948
rect 13913 29892 13917 29948
rect 13853 29888 13917 29892
rect 22054 29948 22118 29952
rect 22054 29892 22058 29948
rect 22058 29892 22114 29948
rect 22114 29892 22118 29948
rect 22054 29888 22118 29892
rect 22134 29948 22198 29952
rect 22134 29892 22138 29948
rect 22138 29892 22194 29948
rect 22194 29892 22198 29948
rect 22134 29888 22198 29892
rect 22214 29948 22278 29952
rect 22214 29892 22218 29948
rect 22218 29892 22274 29948
rect 22274 29892 22278 29948
rect 22214 29888 22278 29892
rect 22294 29948 22358 29952
rect 22294 29892 22298 29948
rect 22298 29892 22354 29948
rect 22354 29892 22358 29948
rect 22294 29888 22358 29892
rect 30495 29948 30559 29952
rect 30495 29892 30499 29948
rect 30499 29892 30555 29948
rect 30555 29892 30559 29948
rect 30495 29888 30559 29892
rect 30575 29948 30639 29952
rect 30575 29892 30579 29948
rect 30579 29892 30635 29948
rect 30635 29892 30639 29948
rect 30575 29888 30639 29892
rect 30655 29948 30719 29952
rect 30655 29892 30659 29948
rect 30659 29892 30715 29948
rect 30715 29892 30719 29948
rect 30655 29888 30719 29892
rect 30735 29948 30799 29952
rect 30735 29892 30739 29948
rect 30739 29892 30795 29948
rect 30795 29892 30799 29948
rect 30735 29888 30799 29892
rect 9392 29404 9456 29408
rect 9392 29348 9396 29404
rect 9396 29348 9452 29404
rect 9452 29348 9456 29404
rect 9392 29344 9456 29348
rect 9472 29404 9536 29408
rect 9472 29348 9476 29404
rect 9476 29348 9532 29404
rect 9532 29348 9536 29404
rect 9472 29344 9536 29348
rect 9552 29404 9616 29408
rect 9552 29348 9556 29404
rect 9556 29348 9612 29404
rect 9612 29348 9616 29404
rect 9552 29344 9616 29348
rect 9632 29404 9696 29408
rect 9632 29348 9636 29404
rect 9636 29348 9692 29404
rect 9692 29348 9696 29404
rect 9632 29344 9696 29348
rect 17833 29404 17897 29408
rect 17833 29348 17837 29404
rect 17837 29348 17893 29404
rect 17893 29348 17897 29404
rect 17833 29344 17897 29348
rect 17913 29404 17977 29408
rect 17913 29348 17917 29404
rect 17917 29348 17973 29404
rect 17973 29348 17977 29404
rect 17913 29344 17977 29348
rect 17993 29404 18057 29408
rect 17993 29348 17997 29404
rect 17997 29348 18053 29404
rect 18053 29348 18057 29404
rect 17993 29344 18057 29348
rect 18073 29404 18137 29408
rect 18073 29348 18077 29404
rect 18077 29348 18133 29404
rect 18133 29348 18137 29404
rect 18073 29344 18137 29348
rect 26274 29404 26338 29408
rect 26274 29348 26278 29404
rect 26278 29348 26334 29404
rect 26334 29348 26338 29404
rect 26274 29344 26338 29348
rect 26354 29404 26418 29408
rect 26354 29348 26358 29404
rect 26358 29348 26414 29404
rect 26414 29348 26418 29404
rect 26354 29344 26418 29348
rect 26434 29404 26498 29408
rect 26434 29348 26438 29404
rect 26438 29348 26494 29404
rect 26494 29348 26498 29404
rect 26434 29344 26498 29348
rect 26514 29404 26578 29408
rect 26514 29348 26518 29404
rect 26518 29348 26574 29404
rect 26574 29348 26578 29404
rect 26514 29344 26578 29348
rect 34715 29404 34779 29408
rect 34715 29348 34719 29404
rect 34719 29348 34775 29404
rect 34775 29348 34779 29404
rect 34715 29344 34779 29348
rect 34795 29404 34859 29408
rect 34795 29348 34799 29404
rect 34799 29348 34855 29404
rect 34855 29348 34859 29404
rect 34795 29344 34859 29348
rect 34875 29404 34939 29408
rect 34875 29348 34879 29404
rect 34879 29348 34935 29404
rect 34935 29348 34939 29404
rect 34875 29344 34939 29348
rect 34955 29404 35019 29408
rect 34955 29348 34959 29404
rect 34959 29348 35015 29404
rect 35015 29348 35019 29404
rect 34955 29344 35019 29348
rect 5172 28860 5236 28864
rect 5172 28804 5176 28860
rect 5176 28804 5232 28860
rect 5232 28804 5236 28860
rect 5172 28800 5236 28804
rect 5252 28860 5316 28864
rect 5252 28804 5256 28860
rect 5256 28804 5312 28860
rect 5312 28804 5316 28860
rect 5252 28800 5316 28804
rect 5332 28860 5396 28864
rect 5332 28804 5336 28860
rect 5336 28804 5392 28860
rect 5392 28804 5396 28860
rect 5332 28800 5396 28804
rect 5412 28860 5476 28864
rect 5412 28804 5416 28860
rect 5416 28804 5472 28860
rect 5472 28804 5476 28860
rect 5412 28800 5476 28804
rect 13613 28860 13677 28864
rect 13613 28804 13617 28860
rect 13617 28804 13673 28860
rect 13673 28804 13677 28860
rect 13613 28800 13677 28804
rect 13693 28860 13757 28864
rect 13693 28804 13697 28860
rect 13697 28804 13753 28860
rect 13753 28804 13757 28860
rect 13693 28800 13757 28804
rect 13773 28860 13837 28864
rect 13773 28804 13777 28860
rect 13777 28804 13833 28860
rect 13833 28804 13837 28860
rect 13773 28800 13837 28804
rect 13853 28860 13917 28864
rect 13853 28804 13857 28860
rect 13857 28804 13913 28860
rect 13913 28804 13917 28860
rect 13853 28800 13917 28804
rect 22054 28860 22118 28864
rect 22054 28804 22058 28860
rect 22058 28804 22114 28860
rect 22114 28804 22118 28860
rect 22054 28800 22118 28804
rect 22134 28860 22198 28864
rect 22134 28804 22138 28860
rect 22138 28804 22194 28860
rect 22194 28804 22198 28860
rect 22134 28800 22198 28804
rect 22214 28860 22278 28864
rect 22214 28804 22218 28860
rect 22218 28804 22274 28860
rect 22274 28804 22278 28860
rect 22214 28800 22278 28804
rect 22294 28860 22358 28864
rect 22294 28804 22298 28860
rect 22298 28804 22354 28860
rect 22354 28804 22358 28860
rect 22294 28800 22358 28804
rect 30495 28860 30559 28864
rect 30495 28804 30499 28860
rect 30499 28804 30555 28860
rect 30555 28804 30559 28860
rect 30495 28800 30559 28804
rect 30575 28860 30639 28864
rect 30575 28804 30579 28860
rect 30579 28804 30635 28860
rect 30635 28804 30639 28860
rect 30575 28800 30639 28804
rect 30655 28860 30719 28864
rect 30655 28804 30659 28860
rect 30659 28804 30715 28860
rect 30715 28804 30719 28860
rect 30655 28800 30719 28804
rect 30735 28860 30799 28864
rect 30735 28804 30739 28860
rect 30739 28804 30795 28860
rect 30795 28804 30799 28860
rect 30735 28800 30799 28804
rect 9392 28316 9456 28320
rect 9392 28260 9396 28316
rect 9396 28260 9452 28316
rect 9452 28260 9456 28316
rect 9392 28256 9456 28260
rect 9472 28316 9536 28320
rect 9472 28260 9476 28316
rect 9476 28260 9532 28316
rect 9532 28260 9536 28316
rect 9472 28256 9536 28260
rect 9552 28316 9616 28320
rect 9552 28260 9556 28316
rect 9556 28260 9612 28316
rect 9612 28260 9616 28316
rect 9552 28256 9616 28260
rect 9632 28316 9696 28320
rect 9632 28260 9636 28316
rect 9636 28260 9692 28316
rect 9692 28260 9696 28316
rect 9632 28256 9696 28260
rect 17833 28316 17897 28320
rect 17833 28260 17837 28316
rect 17837 28260 17893 28316
rect 17893 28260 17897 28316
rect 17833 28256 17897 28260
rect 17913 28316 17977 28320
rect 17913 28260 17917 28316
rect 17917 28260 17973 28316
rect 17973 28260 17977 28316
rect 17913 28256 17977 28260
rect 17993 28316 18057 28320
rect 17993 28260 17997 28316
rect 17997 28260 18053 28316
rect 18053 28260 18057 28316
rect 17993 28256 18057 28260
rect 18073 28316 18137 28320
rect 18073 28260 18077 28316
rect 18077 28260 18133 28316
rect 18133 28260 18137 28316
rect 18073 28256 18137 28260
rect 26274 28316 26338 28320
rect 26274 28260 26278 28316
rect 26278 28260 26334 28316
rect 26334 28260 26338 28316
rect 26274 28256 26338 28260
rect 26354 28316 26418 28320
rect 26354 28260 26358 28316
rect 26358 28260 26414 28316
rect 26414 28260 26418 28316
rect 26354 28256 26418 28260
rect 26434 28316 26498 28320
rect 26434 28260 26438 28316
rect 26438 28260 26494 28316
rect 26494 28260 26498 28316
rect 26434 28256 26498 28260
rect 26514 28316 26578 28320
rect 26514 28260 26518 28316
rect 26518 28260 26574 28316
rect 26574 28260 26578 28316
rect 26514 28256 26578 28260
rect 34715 28316 34779 28320
rect 34715 28260 34719 28316
rect 34719 28260 34775 28316
rect 34775 28260 34779 28316
rect 34715 28256 34779 28260
rect 34795 28316 34859 28320
rect 34795 28260 34799 28316
rect 34799 28260 34855 28316
rect 34855 28260 34859 28316
rect 34795 28256 34859 28260
rect 34875 28316 34939 28320
rect 34875 28260 34879 28316
rect 34879 28260 34935 28316
rect 34935 28260 34939 28316
rect 34875 28256 34939 28260
rect 34955 28316 35019 28320
rect 34955 28260 34959 28316
rect 34959 28260 35015 28316
rect 35015 28260 35019 28316
rect 34955 28256 35019 28260
rect 5172 27772 5236 27776
rect 5172 27716 5176 27772
rect 5176 27716 5232 27772
rect 5232 27716 5236 27772
rect 5172 27712 5236 27716
rect 5252 27772 5316 27776
rect 5252 27716 5256 27772
rect 5256 27716 5312 27772
rect 5312 27716 5316 27772
rect 5252 27712 5316 27716
rect 5332 27772 5396 27776
rect 5332 27716 5336 27772
rect 5336 27716 5392 27772
rect 5392 27716 5396 27772
rect 5332 27712 5396 27716
rect 5412 27772 5476 27776
rect 5412 27716 5416 27772
rect 5416 27716 5472 27772
rect 5472 27716 5476 27772
rect 5412 27712 5476 27716
rect 13613 27772 13677 27776
rect 13613 27716 13617 27772
rect 13617 27716 13673 27772
rect 13673 27716 13677 27772
rect 13613 27712 13677 27716
rect 13693 27772 13757 27776
rect 13693 27716 13697 27772
rect 13697 27716 13753 27772
rect 13753 27716 13757 27772
rect 13693 27712 13757 27716
rect 13773 27772 13837 27776
rect 13773 27716 13777 27772
rect 13777 27716 13833 27772
rect 13833 27716 13837 27772
rect 13773 27712 13837 27716
rect 13853 27772 13917 27776
rect 13853 27716 13857 27772
rect 13857 27716 13913 27772
rect 13913 27716 13917 27772
rect 13853 27712 13917 27716
rect 22054 27772 22118 27776
rect 22054 27716 22058 27772
rect 22058 27716 22114 27772
rect 22114 27716 22118 27772
rect 22054 27712 22118 27716
rect 22134 27772 22198 27776
rect 22134 27716 22138 27772
rect 22138 27716 22194 27772
rect 22194 27716 22198 27772
rect 22134 27712 22198 27716
rect 22214 27772 22278 27776
rect 22214 27716 22218 27772
rect 22218 27716 22274 27772
rect 22274 27716 22278 27772
rect 22214 27712 22278 27716
rect 22294 27772 22358 27776
rect 22294 27716 22298 27772
rect 22298 27716 22354 27772
rect 22354 27716 22358 27772
rect 22294 27712 22358 27716
rect 30495 27772 30559 27776
rect 30495 27716 30499 27772
rect 30499 27716 30555 27772
rect 30555 27716 30559 27772
rect 30495 27712 30559 27716
rect 30575 27772 30639 27776
rect 30575 27716 30579 27772
rect 30579 27716 30635 27772
rect 30635 27716 30639 27772
rect 30575 27712 30639 27716
rect 30655 27772 30719 27776
rect 30655 27716 30659 27772
rect 30659 27716 30715 27772
rect 30715 27716 30719 27772
rect 30655 27712 30719 27716
rect 30735 27772 30799 27776
rect 30735 27716 30739 27772
rect 30739 27716 30795 27772
rect 30795 27716 30799 27772
rect 30735 27712 30799 27716
rect 9392 27228 9456 27232
rect 9392 27172 9396 27228
rect 9396 27172 9452 27228
rect 9452 27172 9456 27228
rect 9392 27168 9456 27172
rect 9472 27228 9536 27232
rect 9472 27172 9476 27228
rect 9476 27172 9532 27228
rect 9532 27172 9536 27228
rect 9472 27168 9536 27172
rect 9552 27228 9616 27232
rect 9552 27172 9556 27228
rect 9556 27172 9612 27228
rect 9612 27172 9616 27228
rect 9552 27168 9616 27172
rect 9632 27228 9696 27232
rect 9632 27172 9636 27228
rect 9636 27172 9692 27228
rect 9692 27172 9696 27228
rect 9632 27168 9696 27172
rect 17833 27228 17897 27232
rect 17833 27172 17837 27228
rect 17837 27172 17893 27228
rect 17893 27172 17897 27228
rect 17833 27168 17897 27172
rect 17913 27228 17977 27232
rect 17913 27172 17917 27228
rect 17917 27172 17973 27228
rect 17973 27172 17977 27228
rect 17913 27168 17977 27172
rect 17993 27228 18057 27232
rect 17993 27172 17997 27228
rect 17997 27172 18053 27228
rect 18053 27172 18057 27228
rect 17993 27168 18057 27172
rect 18073 27228 18137 27232
rect 18073 27172 18077 27228
rect 18077 27172 18133 27228
rect 18133 27172 18137 27228
rect 18073 27168 18137 27172
rect 26274 27228 26338 27232
rect 26274 27172 26278 27228
rect 26278 27172 26334 27228
rect 26334 27172 26338 27228
rect 26274 27168 26338 27172
rect 26354 27228 26418 27232
rect 26354 27172 26358 27228
rect 26358 27172 26414 27228
rect 26414 27172 26418 27228
rect 26354 27168 26418 27172
rect 26434 27228 26498 27232
rect 26434 27172 26438 27228
rect 26438 27172 26494 27228
rect 26494 27172 26498 27228
rect 26434 27168 26498 27172
rect 26514 27228 26578 27232
rect 26514 27172 26518 27228
rect 26518 27172 26574 27228
rect 26574 27172 26578 27228
rect 26514 27168 26578 27172
rect 34715 27228 34779 27232
rect 34715 27172 34719 27228
rect 34719 27172 34775 27228
rect 34775 27172 34779 27228
rect 34715 27168 34779 27172
rect 34795 27228 34859 27232
rect 34795 27172 34799 27228
rect 34799 27172 34855 27228
rect 34855 27172 34859 27228
rect 34795 27168 34859 27172
rect 34875 27228 34939 27232
rect 34875 27172 34879 27228
rect 34879 27172 34935 27228
rect 34935 27172 34939 27228
rect 34875 27168 34939 27172
rect 34955 27228 35019 27232
rect 34955 27172 34959 27228
rect 34959 27172 35015 27228
rect 35015 27172 35019 27228
rect 34955 27168 35019 27172
rect 5172 26684 5236 26688
rect 5172 26628 5176 26684
rect 5176 26628 5232 26684
rect 5232 26628 5236 26684
rect 5172 26624 5236 26628
rect 5252 26684 5316 26688
rect 5252 26628 5256 26684
rect 5256 26628 5312 26684
rect 5312 26628 5316 26684
rect 5252 26624 5316 26628
rect 5332 26684 5396 26688
rect 5332 26628 5336 26684
rect 5336 26628 5392 26684
rect 5392 26628 5396 26684
rect 5332 26624 5396 26628
rect 5412 26684 5476 26688
rect 5412 26628 5416 26684
rect 5416 26628 5472 26684
rect 5472 26628 5476 26684
rect 5412 26624 5476 26628
rect 13613 26684 13677 26688
rect 13613 26628 13617 26684
rect 13617 26628 13673 26684
rect 13673 26628 13677 26684
rect 13613 26624 13677 26628
rect 13693 26684 13757 26688
rect 13693 26628 13697 26684
rect 13697 26628 13753 26684
rect 13753 26628 13757 26684
rect 13693 26624 13757 26628
rect 13773 26684 13837 26688
rect 13773 26628 13777 26684
rect 13777 26628 13833 26684
rect 13833 26628 13837 26684
rect 13773 26624 13837 26628
rect 13853 26684 13917 26688
rect 13853 26628 13857 26684
rect 13857 26628 13913 26684
rect 13913 26628 13917 26684
rect 13853 26624 13917 26628
rect 22054 26684 22118 26688
rect 22054 26628 22058 26684
rect 22058 26628 22114 26684
rect 22114 26628 22118 26684
rect 22054 26624 22118 26628
rect 22134 26684 22198 26688
rect 22134 26628 22138 26684
rect 22138 26628 22194 26684
rect 22194 26628 22198 26684
rect 22134 26624 22198 26628
rect 22214 26684 22278 26688
rect 22214 26628 22218 26684
rect 22218 26628 22274 26684
rect 22274 26628 22278 26684
rect 22214 26624 22278 26628
rect 22294 26684 22358 26688
rect 22294 26628 22298 26684
rect 22298 26628 22354 26684
rect 22354 26628 22358 26684
rect 22294 26624 22358 26628
rect 30495 26684 30559 26688
rect 30495 26628 30499 26684
rect 30499 26628 30555 26684
rect 30555 26628 30559 26684
rect 30495 26624 30559 26628
rect 30575 26684 30639 26688
rect 30575 26628 30579 26684
rect 30579 26628 30635 26684
rect 30635 26628 30639 26684
rect 30575 26624 30639 26628
rect 30655 26684 30719 26688
rect 30655 26628 30659 26684
rect 30659 26628 30715 26684
rect 30715 26628 30719 26684
rect 30655 26624 30719 26628
rect 30735 26684 30799 26688
rect 30735 26628 30739 26684
rect 30739 26628 30795 26684
rect 30795 26628 30799 26684
rect 30735 26624 30799 26628
rect 9392 26140 9456 26144
rect 9392 26084 9396 26140
rect 9396 26084 9452 26140
rect 9452 26084 9456 26140
rect 9392 26080 9456 26084
rect 9472 26140 9536 26144
rect 9472 26084 9476 26140
rect 9476 26084 9532 26140
rect 9532 26084 9536 26140
rect 9472 26080 9536 26084
rect 9552 26140 9616 26144
rect 9552 26084 9556 26140
rect 9556 26084 9612 26140
rect 9612 26084 9616 26140
rect 9552 26080 9616 26084
rect 9632 26140 9696 26144
rect 9632 26084 9636 26140
rect 9636 26084 9692 26140
rect 9692 26084 9696 26140
rect 9632 26080 9696 26084
rect 17833 26140 17897 26144
rect 17833 26084 17837 26140
rect 17837 26084 17893 26140
rect 17893 26084 17897 26140
rect 17833 26080 17897 26084
rect 17913 26140 17977 26144
rect 17913 26084 17917 26140
rect 17917 26084 17973 26140
rect 17973 26084 17977 26140
rect 17913 26080 17977 26084
rect 17993 26140 18057 26144
rect 17993 26084 17997 26140
rect 17997 26084 18053 26140
rect 18053 26084 18057 26140
rect 17993 26080 18057 26084
rect 18073 26140 18137 26144
rect 18073 26084 18077 26140
rect 18077 26084 18133 26140
rect 18133 26084 18137 26140
rect 18073 26080 18137 26084
rect 26274 26140 26338 26144
rect 26274 26084 26278 26140
rect 26278 26084 26334 26140
rect 26334 26084 26338 26140
rect 26274 26080 26338 26084
rect 26354 26140 26418 26144
rect 26354 26084 26358 26140
rect 26358 26084 26414 26140
rect 26414 26084 26418 26140
rect 26354 26080 26418 26084
rect 26434 26140 26498 26144
rect 26434 26084 26438 26140
rect 26438 26084 26494 26140
rect 26494 26084 26498 26140
rect 26434 26080 26498 26084
rect 26514 26140 26578 26144
rect 26514 26084 26518 26140
rect 26518 26084 26574 26140
rect 26574 26084 26578 26140
rect 26514 26080 26578 26084
rect 34715 26140 34779 26144
rect 34715 26084 34719 26140
rect 34719 26084 34775 26140
rect 34775 26084 34779 26140
rect 34715 26080 34779 26084
rect 34795 26140 34859 26144
rect 34795 26084 34799 26140
rect 34799 26084 34855 26140
rect 34855 26084 34859 26140
rect 34795 26080 34859 26084
rect 34875 26140 34939 26144
rect 34875 26084 34879 26140
rect 34879 26084 34935 26140
rect 34935 26084 34939 26140
rect 34875 26080 34939 26084
rect 34955 26140 35019 26144
rect 34955 26084 34959 26140
rect 34959 26084 35015 26140
rect 35015 26084 35019 26140
rect 34955 26080 35019 26084
rect 5172 25596 5236 25600
rect 5172 25540 5176 25596
rect 5176 25540 5232 25596
rect 5232 25540 5236 25596
rect 5172 25536 5236 25540
rect 5252 25596 5316 25600
rect 5252 25540 5256 25596
rect 5256 25540 5312 25596
rect 5312 25540 5316 25596
rect 5252 25536 5316 25540
rect 5332 25596 5396 25600
rect 5332 25540 5336 25596
rect 5336 25540 5392 25596
rect 5392 25540 5396 25596
rect 5332 25536 5396 25540
rect 5412 25596 5476 25600
rect 5412 25540 5416 25596
rect 5416 25540 5472 25596
rect 5472 25540 5476 25596
rect 5412 25536 5476 25540
rect 13613 25596 13677 25600
rect 13613 25540 13617 25596
rect 13617 25540 13673 25596
rect 13673 25540 13677 25596
rect 13613 25536 13677 25540
rect 13693 25596 13757 25600
rect 13693 25540 13697 25596
rect 13697 25540 13753 25596
rect 13753 25540 13757 25596
rect 13693 25536 13757 25540
rect 13773 25596 13837 25600
rect 13773 25540 13777 25596
rect 13777 25540 13833 25596
rect 13833 25540 13837 25596
rect 13773 25536 13837 25540
rect 13853 25596 13917 25600
rect 13853 25540 13857 25596
rect 13857 25540 13913 25596
rect 13913 25540 13917 25596
rect 13853 25536 13917 25540
rect 22054 25596 22118 25600
rect 22054 25540 22058 25596
rect 22058 25540 22114 25596
rect 22114 25540 22118 25596
rect 22054 25536 22118 25540
rect 22134 25596 22198 25600
rect 22134 25540 22138 25596
rect 22138 25540 22194 25596
rect 22194 25540 22198 25596
rect 22134 25536 22198 25540
rect 22214 25596 22278 25600
rect 22214 25540 22218 25596
rect 22218 25540 22274 25596
rect 22274 25540 22278 25596
rect 22214 25536 22278 25540
rect 22294 25596 22358 25600
rect 22294 25540 22298 25596
rect 22298 25540 22354 25596
rect 22354 25540 22358 25596
rect 22294 25536 22358 25540
rect 30495 25596 30559 25600
rect 30495 25540 30499 25596
rect 30499 25540 30555 25596
rect 30555 25540 30559 25596
rect 30495 25536 30559 25540
rect 30575 25596 30639 25600
rect 30575 25540 30579 25596
rect 30579 25540 30635 25596
rect 30635 25540 30639 25596
rect 30575 25536 30639 25540
rect 30655 25596 30719 25600
rect 30655 25540 30659 25596
rect 30659 25540 30715 25596
rect 30715 25540 30719 25596
rect 30655 25536 30719 25540
rect 30735 25596 30799 25600
rect 30735 25540 30739 25596
rect 30739 25540 30795 25596
rect 30795 25540 30799 25596
rect 30735 25536 30799 25540
rect 9392 25052 9456 25056
rect 9392 24996 9396 25052
rect 9396 24996 9452 25052
rect 9452 24996 9456 25052
rect 9392 24992 9456 24996
rect 9472 25052 9536 25056
rect 9472 24996 9476 25052
rect 9476 24996 9532 25052
rect 9532 24996 9536 25052
rect 9472 24992 9536 24996
rect 9552 25052 9616 25056
rect 9552 24996 9556 25052
rect 9556 24996 9612 25052
rect 9612 24996 9616 25052
rect 9552 24992 9616 24996
rect 9632 25052 9696 25056
rect 9632 24996 9636 25052
rect 9636 24996 9692 25052
rect 9692 24996 9696 25052
rect 9632 24992 9696 24996
rect 17833 25052 17897 25056
rect 17833 24996 17837 25052
rect 17837 24996 17893 25052
rect 17893 24996 17897 25052
rect 17833 24992 17897 24996
rect 17913 25052 17977 25056
rect 17913 24996 17917 25052
rect 17917 24996 17973 25052
rect 17973 24996 17977 25052
rect 17913 24992 17977 24996
rect 17993 25052 18057 25056
rect 17993 24996 17997 25052
rect 17997 24996 18053 25052
rect 18053 24996 18057 25052
rect 17993 24992 18057 24996
rect 18073 25052 18137 25056
rect 18073 24996 18077 25052
rect 18077 24996 18133 25052
rect 18133 24996 18137 25052
rect 18073 24992 18137 24996
rect 26274 25052 26338 25056
rect 26274 24996 26278 25052
rect 26278 24996 26334 25052
rect 26334 24996 26338 25052
rect 26274 24992 26338 24996
rect 26354 25052 26418 25056
rect 26354 24996 26358 25052
rect 26358 24996 26414 25052
rect 26414 24996 26418 25052
rect 26354 24992 26418 24996
rect 26434 25052 26498 25056
rect 26434 24996 26438 25052
rect 26438 24996 26494 25052
rect 26494 24996 26498 25052
rect 26434 24992 26498 24996
rect 26514 25052 26578 25056
rect 26514 24996 26518 25052
rect 26518 24996 26574 25052
rect 26574 24996 26578 25052
rect 26514 24992 26578 24996
rect 34715 25052 34779 25056
rect 34715 24996 34719 25052
rect 34719 24996 34775 25052
rect 34775 24996 34779 25052
rect 34715 24992 34779 24996
rect 34795 25052 34859 25056
rect 34795 24996 34799 25052
rect 34799 24996 34855 25052
rect 34855 24996 34859 25052
rect 34795 24992 34859 24996
rect 34875 25052 34939 25056
rect 34875 24996 34879 25052
rect 34879 24996 34935 25052
rect 34935 24996 34939 25052
rect 34875 24992 34939 24996
rect 34955 25052 35019 25056
rect 34955 24996 34959 25052
rect 34959 24996 35015 25052
rect 35015 24996 35019 25052
rect 34955 24992 35019 24996
rect 5172 24508 5236 24512
rect 5172 24452 5176 24508
rect 5176 24452 5232 24508
rect 5232 24452 5236 24508
rect 5172 24448 5236 24452
rect 5252 24508 5316 24512
rect 5252 24452 5256 24508
rect 5256 24452 5312 24508
rect 5312 24452 5316 24508
rect 5252 24448 5316 24452
rect 5332 24508 5396 24512
rect 5332 24452 5336 24508
rect 5336 24452 5392 24508
rect 5392 24452 5396 24508
rect 5332 24448 5396 24452
rect 5412 24508 5476 24512
rect 5412 24452 5416 24508
rect 5416 24452 5472 24508
rect 5472 24452 5476 24508
rect 5412 24448 5476 24452
rect 13613 24508 13677 24512
rect 13613 24452 13617 24508
rect 13617 24452 13673 24508
rect 13673 24452 13677 24508
rect 13613 24448 13677 24452
rect 13693 24508 13757 24512
rect 13693 24452 13697 24508
rect 13697 24452 13753 24508
rect 13753 24452 13757 24508
rect 13693 24448 13757 24452
rect 13773 24508 13837 24512
rect 13773 24452 13777 24508
rect 13777 24452 13833 24508
rect 13833 24452 13837 24508
rect 13773 24448 13837 24452
rect 13853 24508 13917 24512
rect 13853 24452 13857 24508
rect 13857 24452 13913 24508
rect 13913 24452 13917 24508
rect 13853 24448 13917 24452
rect 22054 24508 22118 24512
rect 22054 24452 22058 24508
rect 22058 24452 22114 24508
rect 22114 24452 22118 24508
rect 22054 24448 22118 24452
rect 22134 24508 22198 24512
rect 22134 24452 22138 24508
rect 22138 24452 22194 24508
rect 22194 24452 22198 24508
rect 22134 24448 22198 24452
rect 22214 24508 22278 24512
rect 22214 24452 22218 24508
rect 22218 24452 22274 24508
rect 22274 24452 22278 24508
rect 22214 24448 22278 24452
rect 22294 24508 22358 24512
rect 22294 24452 22298 24508
rect 22298 24452 22354 24508
rect 22354 24452 22358 24508
rect 22294 24448 22358 24452
rect 30495 24508 30559 24512
rect 30495 24452 30499 24508
rect 30499 24452 30555 24508
rect 30555 24452 30559 24508
rect 30495 24448 30559 24452
rect 30575 24508 30639 24512
rect 30575 24452 30579 24508
rect 30579 24452 30635 24508
rect 30635 24452 30639 24508
rect 30575 24448 30639 24452
rect 30655 24508 30719 24512
rect 30655 24452 30659 24508
rect 30659 24452 30715 24508
rect 30715 24452 30719 24508
rect 30655 24448 30719 24452
rect 30735 24508 30799 24512
rect 30735 24452 30739 24508
rect 30739 24452 30795 24508
rect 30795 24452 30799 24508
rect 30735 24448 30799 24452
rect 9392 23964 9456 23968
rect 9392 23908 9396 23964
rect 9396 23908 9452 23964
rect 9452 23908 9456 23964
rect 9392 23904 9456 23908
rect 9472 23964 9536 23968
rect 9472 23908 9476 23964
rect 9476 23908 9532 23964
rect 9532 23908 9536 23964
rect 9472 23904 9536 23908
rect 9552 23964 9616 23968
rect 9552 23908 9556 23964
rect 9556 23908 9612 23964
rect 9612 23908 9616 23964
rect 9552 23904 9616 23908
rect 9632 23964 9696 23968
rect 9632 23908 9636 23964
rect 9636 23908 9692 23964
rect 9692 23908 9696 23964
rect 9632 23904 9696 23908
rect 17833 23964 17897 23968
rect 17833 23908 17837 23964
rect 17837 23908 17893 23964
rect 17893 23908 17897 23964
rect 17833 23904 17897 23908
rect 17913 23964 17977 23968
rect 17913 23908 17917 23964
rect 17917 23908 17973 23964
rect 17973 23908 17977 23964
rect 17913 23904 17977 23908
rect 17993 23964 18057 23968
rect 17993 23908 17997 23964
rect 17997 23908 18053 23964
rect 18053 23908 18057 23964
rect 17993 23904 18057 23908
rect 18073 23964 18137 23968
rect 18073 23908 18077 23964
rect 18077 23908 18133 23964
rect 18133 23908 18137 23964
rect 18073 23904 18137 23908
rect 26274 23964 26338 23968
rect 26274 23908 26278 23964
rect 26278 23908 26334 23964
rect 26334 23908 26338 23964
rect 26274 23904 26338 23908
rect 26354 23964 26418 23968
rect 26354 23908 26358 23964
rect 26358 23908 26414 23964
rect 26414 23908 26418 23964
rect 26354 23904 26418 23908
rect 26434 23964 26498 23968
rect 26434 23908 26438 23964
rect 26438 23908 26494 23964
rect 26494 23908 26498 23964
rect 26434 23904 26498 23908
rect 26514 23964 26578 23968
rect 26514 23908 26518 23964
rect 26518 23908 26574 23964
rect 26574 23908 26578 23964
rect 26514 23904 26578 23908
rect 34715 23964 34779 23968
rect 34715 23908 34719 23964
rect 34719 23908 34775 23964
rect 34775 23908 34779 23964
rect 34715 23904 34779 23908
rect 34795 23964 34859 23968
rect 34795 23908 34799 23964
rect 34799 23908 34855 23964
rect 34855 23908 34859 23964
rect 34795 23904 34859 23908
rect 34875 23964 34939 23968
rect 34875 23908 34879 23964
rect 34879 23908 34935 23964
rect 34935 23908 34939 23964
rect 34875 23904 34939 23908
rect 34955 23964 35019 23968
rect 34955 23908 34959 23964
rect 34959 23908 35015 23964
rect 35015 23908 35019 23964
rect 34955 23904 35019 23908
rect 5172 23420 5236 23424
rect 5172 23364 5176 23420
rect 5176 23364 5232 23420
rect 5232 23364 5236 23420
rect 5172 23360 5236 23364
rect 5252 23420 5316 23424
rect 5252 23364 5256 23420
rect 5256 23364 5312 23420
rect 5312 23364 5316 23420
rect 5252 23360 5316 23364
rect 5332 23420 5396 23424
rect 5332 23364 5336 23420
rect 5336 23364 5392 23420
rect 5392 23364 5396 23420
rect 5332 23360 5396 23364
rect 5412 23420 5476 23424
rect 5412 23364 5416 23420
rect 5416 23364 5472 23420
rect 5472 23364 5476 23420
rect 5412 23360 5476 23364
rect 13613 23420 13677 23424
rect 13613 23364 13617 23420
rect 13617 23364 13673 23420
rect 13673 23364 13677 23420
rect 13613 23360 13677 23364
rect 13693 23420 13757 23424
rect 13693 23364 13697 23420
rect 13697 23364 13753 23420
rect 13753 23364 13757 23420
rect 13693 23360 13757 23364
rect 13773 23420 13837 23424
rect 13773 23364 13777 23420
rect 13777 23364 13833 23420
rect 13833 23364 13837 23420
rect 13773 23360 13837 23364
rect 13853 23420 13917 23424
rect 13853 23364 13857 23420
rect 13857 23364 13913 23420
rect 13913 23364 13917 23420
rect 13853 23360 13917 23364
rect 22054 23420 22118 23424
rect 22054 23364 22058 23420
rect 22058 23364 22114 23420
rect 22114 23364 22118 23420
rect 22054 23360 22118 23364
rect 22134 23420 22198 23424
rect 22134 23364 22138 23420
rect 22138 23364 22194 23420
rect 22194 23364 22198 23420
rect 22134 23360 22198 23364
rect 22214 23420 22278 23424
rect 22214 23364 22218 23420
rect 22218 23364 22274 23420
rect 22274 23364 22278 23420
rect 22214 23360 22278 23364
rect 22294 23420 22358 23424
rect 22294 23364 22298 23420
rect 22298 23364 22354 23420
rect 22354 23364 22358 23420
rect 22294 23360 22358 23364
rect 30495 23420 30559 23424
rect 30495 23364 30499 23420
rect 30499 23364 30555 23420
rect 30555 23364 30559 23420
rect 30495 23360 30559 23364
rect 30575 23420 30639 23424
rect 30575 23364 30579 23420
rect 30579 23364 30635 23420
rect 30635 23364 30639 23420
rect 30575 23360 30639 23364
rect 30655 23420 30719 23424
rect 30655 23364 30659 23420
rect 30659 23364 30715 23420
rect 30715 23364 30719 23420
rect 30655 23360 30719 23364
rect 30735 23420 30799 23424
rect 30735 23364 30739 23420
rect 30739 23364 30795 23420
rect 30795 23364 30799 23420
rect 30735 23360 30799 23364
rect 9392 22876 9456 22880
rect 9392 22820 9396 22876
rect 9396 22820 9452 22876
rect 9452 22820 9456 22876
rect 9392 22816 9456 22820
rect 9472 22876 9536 22880
rect 9472 22820 9476 22876
rect 9476 22820 9532 22876
rect 9532 22820 9536 22876
rect 9472 22816 9536 22820
rect 9552 22876 9616 22880
rect 9552 22820 9556 22876
rect 9556 22820 9612 22876
rect 9612 22820 9616 22876
rect 9552 22816 9616 22820
rect 9632 22876 9696 22880
rect 9632 22820 9636 22876
rect 9636 22820 9692 22876
rect 9692 22820 9696 22876
rect 9632 22816 9696 22820
rect 17833 22876 17897 22880
rect 17833 22820 17837 22876
rect 17837 22820 17893 22876
rect 17893 22820 17897 22876
rect 17833 22816 17897 22820
rect 17913 22876 17977 22880
rect 17913 22820 17917 22876
rect 17917 22820 17973 22876
rect 17973 22820 17977 22876
rect 17913 22816 17977 22820
rect 17993 22876 18057 22880
rect 17993 22820 17997 22876
rect 17997 22820 18053 22876
rect 18053 22820 18057 22876
rect 17993 22816 18057 22820
rect 18073 22876 18137 22880
rect 18073 22820 18077 22876
rect 18077 22820 18133 22876
rect 18133 22820 18137 22876
rect 18073 22816 18137 22820
rect 26274 22876 26338 22880
rect 26274 22820 26278 22876
rect 26278 22820 26334 22876
rect 26334 22820 26338 22876
rect 26274 22816 26338 22820
rect 26354 22876 26418 22880
rect 26354 22820 26358 22876
rect 26358 22820 26414 22876
rect 26414 22820 26418 22876
rect 26354 22816 26418 22820
rect 26434 22876 26498 22880
rect 26434 22820 26438 22876
rect 26438 22820 26494 22876
rect 26494 22820 26498 22876
rect 26434 22816 26498 22820
rect 26514 22876 26578 22880
rect 26514 22820 26518 22876
rect 26518 22820 26574 22876
rect 26574 22820 26578 22876
rect 26514 22816 26578 22820
rect 34715 22876 34779 22880
rect 34715 22820 34719 22876
rect 34719 22820 34775 22876
rect 34775 22820 34779 22876
rect 34715 22816 34779 22820
rect 34795 22876 34859 22880
rect 34795 22820 34799 22876
rect 34799 22820 34855 22876
rect 34855 22820 34859 22876
rect 34795 22816 34859 22820
rect 34875 22876 34939 22880
rect 34875 22820 34879 22876
rect 34879 22820 34935 22876
rect 34935 22820 34939 22876
rect 34875 22816 34939 22820
rect 34955 22876 35019 22880
rect 34955 22820 34959 22876
rect 34959 22820 35015 22876
rect 35015 22820 35019 22876
rect 34955 22816 35019 22820
rect 5172 22332 5236 22336
rect 5172 22276 5176 22332
rect 5176 22276 5232 22332
rect 5232 22276 5236 22332
rect 5172 22272 5236 22276
rect 5252 22332 5316 22336
rect 5252 22276 5256 22332
rect 5256 22276 5312 22332
rect 5312 22276 5316 22332
rect 5252 22272 5316 22276
rect 5332 22332 5396 22336
rect 5332 22276 5336 22332
rect 5336 22276 5392 22332
rect 5392 22276 5396 22332
rect 5332 22272 5396 22276
rect 5412 22332 5476 22336
rect 5412 22276 5416 22332
rect 5416 22276 5472 22332
rect 5472 22276 5476 22332
rect 5412 22272 5476 22276
rect 13613 22332 13677 22336
rect 13613 22276 13617 22332
rect 13617 22276 13673 22332
rect 13673 22276 13677 22332
rect 13613 22272 13677 22276
rect 13693 22332 13757 22336
rect 13693 22276 13697 22332
rect 13697 22276 13753 22332
rect 13753 22276 13757 22332
rect 13693 22272 13757 22276
rect 13773 22332 13837 22336
rect 13773 22276 13777 22332
rect 13777 22276 13833 22332
rect 13833 22276 13837 22332
rect 13773 22272 13837 22276
rect 13853 22332 13917 22336
rect 13853 22276 13857 22332
rect 13857 22276 13913 22332
rect 13913 22276 13917 22332
rect 13853 22272 13917 22276
rect 22054 22332 22118 22336
rect 22054 22276 22058 22332
rect 22058 22276 22114 22332
rect 22114 22276 22118 22332
rect 22054 22272 22118 22276
rect 22134 22332 22198 22336
rect 22134 22276 22138 22332
rect 22138 22276 22194 22332
rect 22194 22276 22198 22332
rect 22134 22272 22198 22276
rect 22214 22332 22278 22336
rect 22214 22276 22218 22332
rect 22218 22276 22274 22332
rect 22274 22276 22278 22332
rect 22214 22272 22278 22276
rect 22294 22332 22358 22336
rect 22294 22276 22298 22332
rect 22298 22276 22354 22332
rect 22354 22276 22358 22332
rect 22294 22272 22358 22276
rect 30495 22332 30559 22336
rect 30495 22276 30499 22332
rect 30499 22276 30555 22332
rect 30555 22276 30559 22332
rect 30495 22272 30559 22276
rect 30575 22332 30639 22336
rect 30575 22276 30579 22332
rect 30579 22276 30635 22332
rect 30635 22276 30639 22332
rect 30575 22272 30639 22276
rect 30655 22332 30719 22336
rect 30655 22276 30659 22332
rect 30659 22276 30715 22332
rect 30715 22276 30719 22332
rect 30655 22272 30719 22276
rect 30735 22332 30799 22336
rect 30735 22276 30739 22332
rect 30739 22276 30795 22332
rect 30795 22276 30799 22332
rect 30735 22272 30799 22276
rect 9392 21788 9456 21792
rect 9392 21732 9396 21788
rect 9396 21732 9452 21788
rect 9452 21732 9456 21788
rect 9392 21728 9456 21732
rect 9472 21788 9536 21792
rect 9472 21732 9476 21788
rect 9476 21732 9532 21788
rect 9532 21732 9536 21788
rect 9472 21728 9536 21732
rect 9552 21788 9616 21792
rect 9552 21732 9556 21788
rect 9556 21732 9612 21788
rect 9612 21732 9616 21788
rect 9552 21728 9616 21732
rect 9632 21788 9696 21792
rect 9632 21732 9636 21788
rect 9636 21732 9692 21788
rect 9692 21732 9696 21788
rect 9632 21728 9696 21732
rect 17833 21788 17897 21792
rect 17833 21732 17837 21788
rect 17837 21732 17893 21788
rect 17893 21732 17897 21788
rect 17833 21728 17897 21732
rect 17913 21788 17977 21792
rect 17913 21732 17917 21788
rect 17917 21732 17973 21788
rect 17973 21732 17977 21788
rect 17913 21728 17977 21732
rect 17993 21788 18057 21792
rect 17993 21732 17997 21788
rect 17997 21732 18053 21788
rect 18053 21732 18057 21788
rect 17993 21728 18057 21732
rect 18073 21788 18137 21792
rect 18073 21732 18077 21788
rect 18077 21732 18133 21788
rect 18133 21732 18137 21788
rect 18073 21728 18137 21732
rect 26274 21788 26338 21792
rect 26274 21732 26278 21788
rect 26278 21732 26334 21788
rect 26334 21732 26338 21788
rect 26274 21728 26338 21732
rect 26354 21788 26418 21792
rect 26354 21732 26358 21788
rect 26358 21732 26414 21788
rect 26414 21732 26418 21788
rect 26354 21728 26418 21732
rect 26434 21788 26498 21792
rect 26434 21732 26438 21788
rect 26438 21732 26494 21788
rect 26494 21732 26498 21788
rect 26434 21728 26498 21732
rect 26514 21788 26578 21792
rect 26514 21732 26518 21788
rect 26518 21732 26574 21788
rect 26574 21732 26578 21788
rect 26514 21728 26578 21732
rect 34715 21788 34779 21792
rect 34715 21732 34719 21788
rect 34719 21732 34775 21788
rect 34775 21732 34779 21788
rect 34715 21728 34779 21732
rect 34795 21788 34859 21792
rect 34795 21732 34799 21788
rect 34799 21732 34855 21788
rect 34855 21732 34859 21788
rect 34795 21728 34859 21732
rect 34875 21788 34939 21792
rect 34875 21732 34879 21788
rect 34879 21732 34935 21788
rect 34935 21732 34939 21788
rect 34875 21728 34939 21732
rect 34955 21788 35019 21792
rect 34955 21732 34959 21788
rect 34959 21732 35015 21788
rect 35015 21732 35019 21788
rect 34955 21728 35019 21732
rect 5172 21244 5236 21248
rect 5172 21188 5176 21244
rect 5176 21188 5232 21244
rect 5232 21188 5236 21244
rect 5172 21184 5236 21188
rect 5252 21244 5316 21248
rect 5252 21188 5256 21244
rect 5256 21188 5312 21244
rect 5312 21188 5316 21244
rect 5252 21184 5316 21188
rect 5332 21244 5396 21248
rect 5332 21188 5336 21244
rect 5336 21188 5392 21244
rect 5392 21188 5396 21244
rect 5332 21184 5396 21188
rect 5412 21244 5476 21248
rect 5412 21188 5416 21244
rect 5416 21188 5472 21244
rect 5472 21188 5476 21244
rect 5412 21184 5476 21188
rect 13613 21244 13677 21248
rect 13613 21188 13617 21244
rect 13617 21188 13673 21244
rect 13673 21188 13677 21244
rect 13613 21184 13677 21188
rect 13693 21244 13757 21248
rect 13693 21188 13697 21244
rect 13697 21188 13753 21244
rect 13753 21188 13757 21244
rect 13693 21184 13757 21188
rect 13773 21244 13837 21248
rect 13773 21188 13777 21244
rect 13777 21188 13833 21244
rect 13833 21188 13837 21244
rect 13773 21184 13837 21188
rect 13853 21244 13917 21248
rect 13853 21188 13857 21244
rect 13857 21188 13913 21244
rect 13913 21188 13917 21244
rect 13853 21184 13917 21188
rect 22054 21244 22118 21248
rect 22054 21188 22058 21244
rect 22058 21188 22114 21244
rect 22114 21188 22118 21244
rect 22054 21184 22118 21188
rect 22134 21244 22198 21248
rect 22134 21188 22138 21244
rect 22138 21188 22194 21244
rect 22194 21188 22198 21244
rect 22134 21184 22198 21188
rect 22214 21244 22278 21248
rect 22214 21188 22218 21244
rect 22218 21188 22274 21244
rect 22274 21188 22278 21244
rect 22214 21184 22278 21188
rect 22294 21244 22358 21248
rect 22294 21188 22298 21244
rect 22298 21188 22354 21244
rect 22354 21188 22358 21244
rect 22294 21184 22358 21188
rect 30495 21244 30559 21248
rect 30495 21188 30499 21244
rect 30499 21188 30555 21244
rect 30555 21188 30559 21244
rect 30495 21184 30559 21188
rect 30575 21244 30639 21248
rect 30575 21188 30579 21244
rect 30579 21188 30635 21244
rect 30635 21188 30639 21244
rect 30575 21184 30639 21188
rect 30655 21244 30719 21248
rect 30655 21188 30659 21244
rect 30659 21188 30715 21244
rect 30715 21188 30719 21244
rect 30655 21184 30719 21188
rect 30735 21244 30799 21248
rect 30735 21188 30739 21244
rect 30739 21188 30795 21244
rect 30795 21188 30799 21244
rect 30735 21184 30799 21188
rect 9392 20700 9456 20704
rect 9392 20644 9396 20700
rect 9396 20644 9452 20700
rect 9452 20644 9456 20700
rect 9392 20640 9456 20644
rect 9472 20700 9536 20704
rect 9472 20644 9476 20700
rect 9476 20644 9532 20700
rect 9532 20644 9536 20700
rect 9472 20640 9536 20644
rect 9552 20700 9616 20704
rect 9552 20644 9556 20700
rect 9556 20644 9612 20700
rect 9612 20644 9616 20700
rect 9552 20640 9616 20644
rect 9632 20700 9696 20704
rect 9632 20644 9636 20700
rect 9636 20644 9692 20700
rect 9692 20644 9696 20700
rect 9632 20640 9696 20644
rect 17833 20700 17897 20704
rect 17833 20644 17837 20700
rect 17837 20644 17893 20700
rect 17893 20644 17897 20700
rect 17833 20640 17897 20644
rect 17913 20700 17977 20704
rect 17913 20644 17917 20700
rect 17917 20644 17973 20700
rect 17973 20644 17977 20700
rect 17913 20640 17977 20644
rect 17993 20700 18057 20704
rect 17993 20644 17997 20700
rect 17997 20644 18053 20700
rect 18053 20644 18057 20700
rect 17993 20640 18057 20644
rect 18073 20700 18137 20704
rect 18073 20644 18077 20700
rect 18077 20644 18133 20700
rect 18133 20644 18137 20700
rect 18073 20640 18137 20644
rect 26274 20700 26338 20704
rect 26274 20644 26278 20700
rect 26278 20644 26334 20700
rect 26334 20644 26338 20700
rect 26274 20640 26338 20644
rect 26354 20700 26418 20704
rect 26354 20644 26358 20700
rect 26358 20644 26414 20700
rect 26414 20644 26418 20700
rect 26354 20640 26418 20644
rect 26434 20700 26498 20704
rect 26434 20644 26438 20700
rect 26438 20644 26494 20700
rect 26494 20644 26498 20700
rect 26434 20640 26498 20644
rect 26514 20700 26578 20704
rect 26514 20644 26518 20700
rect 26518 20644 26574 20700
rect 26574 20644 26578 20700
rect 26514 20640 26578 20644
rect 34715 20700 34779 20704
rect 34715 20644 34719 20700
rect 34719 20644 34775 20700
rect 34775 20644 34779 20700
rect 34715 20640 34779 20644
rect 34795 20700 34859 20704
rect 34795 20644 34799 20700
rect 34799 20644 34855 20700
rect 34855 20644 34859 20700
rect 34795 20640 34859 20644
rect 34875 20700 34939 20704
rect 34875 20644 34879 20700
rect 34879 20644 34935 20700
rect 34935 20644 34939 20700
rect 34875 20640 34939 20644
rect 34955 20700 35019 20704
rect 34955 20644 34959 20700
rect 34959 20644 35015 20700
rect 35015 20644 35019 20700
rect 34955 20640 35019 20644
rect 5172 20156 5236 20160
rect 5172 20100 5176 20156
rect 5176 20100 5232 20156
rect 5232 20100 5236 20156
rect 5172 20096 5236 20100
rect 5252 20156 5316 20160
rect 5252 20100 5256 20156
rect 5256 20100 5312 20156
rect 5312 20100 5316 20156
rect 5252 20096 5316 20100
rect 5332 20156 5396 20160
rect 5332 20100 5336 20156
rect 5336 20100 5392 20156
rect 5392 20100 5396 20156
rect 5332 20096 5396 20100
rect 5412 20156 5476 20160
rect 5412 20100 5416 20156
rect 5416 20100 5472 20156
rect 5472 20100 5476 20156
rect 5412 20096 5476 20100
rect 13613 20156 13677 20160
rect 13613 20100 13617 20156
rect 13617 20100 13673 20156
rect 13673 20100 13677 20156
rect 13613 20096 13677 20100
rect 13693 20156 13757 20160
rect 13693 20100 13697 20156
rect 13697 20100 13753 20156
rect 13753 20100 13757 20156
rect 13693 20096 13757 20100
rect 13773 20156 13837 20160
rect 13773 20100 13777 20156
rect 13777 20100 13833 20156
rect 13833 20100 13837 20156
rect 13773 20096 13837 20100
rect 13853 20156 13917 20160
rect 13853 20100 13857 20156
rect 13857 20100 13913 20156
rect 13913 20100 13917 20156
rect 13853 20096 13917 20100
rect 22054 20156 22118 20160
rect 22054 20100 22058 20156
rect 22058 20100 22114 20156
rect 22114 20100 22118 20156
rect 22054 20096 22118 20100
rect 22134 20156 22198 20160
rect 22134 20100 22138 20156
rect 22138 20100 22194 20156
rect 22194 20100 22198 20156
rect 22134 20096 22198 20100
rect 22214 20156 22278 20160
rect 22214 20100 22218 20156
rect 22218 20100 22274 20156
rect 22274 20100 22278 20156
rect 22214 20096 22278 20100
rect 22294 20156 22358 20160
rect 22294 20100 22298 20156
rect 22298 20100 22354 20156
rect 22354 20100 22358 20156
rect 22294 20096 22358 20100
rect 30495 20156 30559 20160
rect 30495 20100 30499 20156
rect 30499 20100 30555 20156
rect 30555 20100 30559 20156
rect 30495 20096 30559 20100
rect 30575 20156 30639 20160
rect 30575 20100 30579 20156
rect 30579 20100 30635 20156
rect 30635 20100 30639 20156
rect 30575 20096 30639 20100
rect 30655 20156 30719 20160
rect 30655 20100 30659 20156
rect 30659 20100 30715 20156
rect 30715 20100 30719 20156
rect 30655 20096 30719 20100
rect 30735 20156 30799 20160
rect 30735 20100 30739 20156
rect 30739 20100 30795 20156
rect 30795 20100 30799 20156
rect 30735 20096 30799 20100
rect 9392 19612 9456 19616
rect 9392 19556 9396 19612
rect 9396 19556 9452 19612
rect 9452 19556 9456 19612
rect 9392 19552 9456 19556
rect 9472 19612 9536 19616
rect 9472 19556 9476 19612
rect 9476 19556 9532 19612
rect 9532 19556 9536 19612
rect 9472 19552 9536 19556
rect 9552 19612 9616 19616
rect 9552 19556 9556 19612
rect 9556 19556 9612 19612
rect 9612 19556 9616 19612
rect 9552 19552 9616 19556
rect 9632 19612 9696 19616
rect 9632 19556 9636 19612
rect 9636 19556 9692 19612
rect 9692 19556 9696 19612
rect 9632 19552 9696 19556
rect 17833 19612 17897 19616
rect 17833 19556 17837 19612
rect 17837 19556 17893 19612
rect 17893 19556 17897 19612
rect 17833 19552 17897 19556
rect 17913 19612 17977 19616
rect 17913 19556 17917 19612
rect 17917 19556 17973 19612
rect 17973 19556 17977 19612
rect 17913 19552 17977 19556
rect 17993 19612 18057 19616
rect 17993 19556 17997 19612
rect 17997 19556 18053 19612
rect 18053 19556 18057 19612
rect 17993 19552 18057 19556
rect 18073 19612 18137 19616
rect 18073 19556 18077 19612
rect 18077 19556 18133 19612
rect 18133 19556 18137 19612
rect 18073 19552 18137 19556
rect 26274 19612 26338 19616
rect 26274 19556 26278 19612
rect 26278 19556 26334 19612
rect 26334 19556 26338 19612
rect 26274 19552 26338 19556
rect 26354 19612 26418 19616
rect 26354 19556 26358 19612
rect 26358 19556 26414 19612
rect 26414 19556 26418 19612
rect 26354 19552 26418 19556
rect 26434 19612 26498 19616
rect 26434 19556 26438 19612
rect 26438 19556 26494 19612
rect 26494 19556 26498 19612
rect 26434 19552 26498 19556
rect 26514 19612 26578 19616
rect 26514 19556 26518 19612
rect 26518 19556 26574 19612
rect 26574 19556 26578 19612
rect 26514 19552 26578 19556
rect 34715 19612 34779 19616
rect 34715 19556 34719 19612
rect 34719 19556 34775 19612
rect 34775 19556 34779 19612
rect 34715 19552 34779 19556
rect 34795 19612 34859 19616
rect 34795 19556 34799 19612
rect 34799 19556 34855 19612
rect 34855 19556 34859 19612
rect 34795 19552 34859 19556
rect 34875 19612 34939 19616
rect 34875 19556 34879 19612
rect 34879 19556 34935 19612
rect 34935 19556 34939 19612
rect 34875 19552 34939 19556
rect 34955 19612 35019 19616
rect 34955 19556 34959 19612
rect 34959 19556 35015 19612
rect 35015 19556 35019 19612
rect 34955 19552 35019 19556
rect 5172 19068 5236 19072
rect 5172 19012 5176 19068
rect 5176 19012 5232 19068
rect 5232 19012 5236 19068
rect 5172 19008 5236 19012
rect 5252 19068 5316 19072
rect 5252 19012 5256 19068
rect 5256 19012 5312 19068
rect 5312 19012 5316 19068
rect 5252 19008 5316 19012
rect 5332 19068 5396 19072
rect 5332 19012 5336 19068
rect 5336 19012 5392 19068
rect 5392 19012 5396 19068
rect 5332 19008 5396 19012
rect 5412 19068 5476 19072
rect 5412 19012 5416 19068
rect 5416 19012 5472 19068
rect 5472 19012 5476 19068
rect 5412 19008 5476 19012
rect 13613 19068 13677 19072
rect 13613 19012 13617 19068
rect 13617 19012 13673 19068
rect 13673 19012 13677 19068
rect 13613 19008 13677 19012
rect 13693 19068 13757 19072
rect 13693 19012 13697 19068
rect 13697 19012 13753 19068
rect 13753 19012 13757 19068
rect 13693 19008 13757 19012
rect 13773 19068 13837 19072
rect 13773 19012 13777 19068
rect 13777 19012 13833 19068
rect 13833 19012 13837 19068
rect 13773 19008 13837 19012
rect 13853 19068 13917 19072
rect 13853 19012 13857 19068
rect 13857 19012 13913 19068
rect 13913 19012 13917 19068
rect 13853 19008 13917 19012
rect 22054 19068 22118 19072
rect 22054 19012 22058 19068
rect 22058 19012 22114 19068
rect 22114 19012 22118 19068
rect 22054 19008 22118 19012
rect 22134 19068 22198 19072
rect 22134 19012 22138 19068
rect 22138 19012 22194 19068
rect 22194 19012 22198 19068
rect 22134 19008 22198 19012
rect 22214 19068 22278 19072
rect 22214 19012 22218 19068
rect 22218 19012 22274 19068
rect 22274 19012 22278 19068
rect 22214 19008 22278 19012
rect 22294 19068 22358 19072
rect 22294 19012 22298 19068
rect 22298 19012 22354 19068
rect 22354 19012 22358 19068
rect 22294 19008 22358 19012
rect 30495 19068 30559 19072
rect 30495 19012 30499 19068
rect 30499 19012 30555 19068
rect 30555 19012 30559 19068
rect 30495 19008 30559 19012
rect 30575 19068 30639 19072
rect 30575 19012 30579 19068
rect 30579 19012 30635 19068
rect 30635 19012 30639 19068
rect 30575 19008 30639 19012
rect 30655 19068 30719 19072
rect 30655 19012 30659 19068
rect 30659 19012 30715 19068
rect 30715 19012 30719 19068
rect 30655 19008 30719 19012
rect 30735 19068 30799 19072
rect 30735 19012 30739 19068
rect 30739 19012 30795 19068
rect 30795 19012 30799 19068
rect 30735 19008 30799 19012
rect 9392 18524 9456 18528
rect 9392 18468 9396 18524
rect 9396 18468 9452 18524
rect 9452 18468 9456 18524
rect 9392 18464 9456 18468
rect 9472 18524 9536 18528
rect 9472 18468 9476 18524
rect 9476 18468 9532 18524
rect 9532 18468 9536 18524
rect 9472 18464 9536 18468
rect 9552 18524 9616 18528
rect 9552 18468 9556 18524
rect 9556 18468 9612 18524
rect 9612 18468 9616 18524
rect 9552 18464 9616 18468
rect 9632 18524 9696 18528
rect 9632 18468 9636 18524
rect 9636 18468 9692 18524
rect 9692 18468 9696 18524
rect 9632 18464 9696 18468
rect 17833 18524 17897 18528
rect 17833 18468 17837 18524
rect 17837 18468 17893 18524
rect 17893 18468 17897 18524
rect 17833 18464 17897 18468
rect 17913 18524 17977 18528
rect 17913 18468 17917 18524
rect 17917 18468 17973 18524
rect 17973 18468 17977 18524
rect 17913 18464 17977 18468
rect 17993 18524 18057 18528
rect 17993 18468 17997 18524
rect 17997 18468 18053 18524
rect 18053 18468 18057 18524
rect 17993 18464 18057 18468
rect 18073 18524 18137 18528
rect 18073 18468 18077 18524
rect 18077 18468 18133 18524
rect 18133 18468 18137 18524
rect 18073 18464 18137 18468
rect 26274 18524 26338 18528
rect 26274 18468 26278 18524
rect 26278 18468 26334 18524
rect 26334 18468 26338 18524
rect 26274 18464 26338 18468
rect 26354 18524 26418 18528
rect 26354 18468 26358 18524
rect 26358 18468 26414 18524
rect 26414 18468 26418 18524
rect 26354 18464 26418 18468
rect 26434 18524 26498 18528
rect 26434 18468 26438 18524
rect 26438 18468 26494 18524
rect 26494 18468 26498 18524
rect 26434 18464 26498 18468
rect 26514 18524 26578 18528
rect 26514 18468 26518 18524
rect 26518 18468 26574 18524
rect 26574 18468 26578 18524
rect 26514 18464 26578 18468
rect 34715 18524 34779 18528
rect 34715 18468 34719 18524
rect 34719 18468 34775 18524
rect 34775 18468 34779 18524
rect 34715 18464 34779 18468
rect 34795 18524 34859 18528
rect 34795 18468 34799 18524
rect 34799 18468 34855 18524
rect 34855 18468 34859 18524
rect 34795 18464 34859 18468
rect 34875 18524 34939 18528
rect 34875 18468 34879 18524
rect 34879 18468 34935 18524
rect 34935 18468 34939 18524
rect 34875 18464 34939 18468
rect 34955 18524 35019 18528
rect 34955 18468 34959 18524
rect 34959 18468 35015 18524
rect 35015 18468 35019 18524
rect 34955 18464 35019 18468
rect 5172 17980 5236 17984
rect 5172 17924 5176 17980
rect 5176 17924 5232 17980
rect 5232 17924 5236 17980
rect 5172 17920 5236 17924
rect 5252 17980 5316 17984
rect 5252 17924 5256 17980
rect 5256 17924 5312 17980
rect 5312 17924 5316 17980
rect 5252 17920 5316 17924
rect 5332 17980 5396 17984
rect 5332 17924 5336 17980
rect 5336 17924 5392 17980
rect 5392 17924 5396 17980
rect 5332 17920 5396 17924
rect 5412 17980 5476 17984
rect 5412 17924 5416 17980
rect 5416 17924 5472 17980
rect 5472 17924 5476 17980
rect 5412 17920 5476 17924
rect 13613 17980 13677 17984
rect 13613 17924 13617 17980
rect 13617 17924 13673 17980
rect 13673 17924 13677 17980
rect 13613 17920 13677 17924
rect 13693 17980 13757 17984
rect 13693 17924 13697 17980
rect 13697 17924 13753 17980
rect 13753 17924 13757 17980
rect 13693 17920 13757 17924
rect 13773 17980 13837 17984
rect 13773 17924 13777 17980
rect 13777 17924 13833 17980
rect 13833 17924 13837 17980
rect 13773 17920 13837 17924
rect 13853 17980 13917 17984
rect 13853 17924 13857 17980
rect 13857 17924 13913 17980
rect 13913 17924 13917 17980
rect 13853 17920 13917 17924
rect 22054 17980 22118 17984
rect 22054 17924 22058 17980
rect 22058 17924 22114 17980
rect 22114 17924 22118 17980
rect 22054 17920 22118 17924
rect 22134 17980 22198 17984
rect 22134 17924 22138 17980
rect 22138 17924 22194 17980
rect 22194 17924 22198 17980
rect 22134 17920 22198 17924
rect 22214 17980 22278 17984
rect 22214 17924 22218 17980
rect 22218 17924 22274 17980
rect 22274 17924 22278 17980
rect 22214 17920 22278 17924
rect 22294 17980 22358 17984
rect 22294 17924 22298 17980
rect 22298 17924 22354 17980
rect 22354 17924 22358 17980
rect 22294 17920 22358 17924
rect 30495 17980 30559 17984
rect 30495 17924 30499 17980
rect 30499 17924 30555 17980
rect 30555 17924 30559 17980
rect 30495 17920 30559 17924
rect 30575 17980 30639 17984
rect 30575 17924 30579 17980
rect 30579 17924 30635 17980
rect 30635 17924 30639 17980
rect 30575 17920 30639 17924
rect 30655 17980 30719 17984
rect 30655 17924 30659 17980
rect 30659 17924 30715 17980
rect 30715 17924 30719 17980
rect 30655 17920 30719 17924
rect 30735 17980 30799 17984
rect 30735 17924 30739 17980
rect 30739 17924 30795 17980
rect 30795 17924 30799 17980
rect 30735 17920 30799 17924
rect 9392 17436 9456 17440
rect 9392 17380 9396 17436
rect 9396 17380 9452 17436
rect 9452 17380 9456 17436
rect 9392 17376 9456 17380
rect 9472 17436 9536 17440
rect 9472 17380 9476 17436
rect 9476 17380 9532 17436
rect 9532 17380 9536 17436
rect 9472 17376 9536 17380
rect 9552 17436 9616 17440
rect 9552 17380 9556 17436
rect 9556 17380 9612 17436
rect 9612 17380 9616 17436
rect 9552 17376 9616 17380
rect 9632 17436 9696 17440
rect 9632 17380 9636 17436
rect 9636 17380 9692 17436
rect 9692 17380 9696 17436
rect 9632 17376 9696 17380
rect 17833 17436 17897 17440
rect 17833 17380 17837 17436
rect 17837 17380 17893 17436
rect 17893 17380 17897 17436
rect 17833 17376 17897 17380
rect 17913 17436 17977 17440
rect 17913 17380 17917 17436
rect 17917 17380 17973 17436
rect 17973 17380 17977 17436
rect 17913 17376 17977 17380
rect 17993 17436 18057 17440
rect 17993 17380 17997 17436
rect 17997 17380 18053 17436
rect 18053 17380 18057 17436
rect 17993 17376 18057 17380
rect 18073 17436 18137 17440
rect 18073 17380 18077 17436
rect 18077 17380 18133 17436
rect 18133 17380 18137 17436
rect 18073 17376 18137 17380
rect 26274 17436 26338 17440
rect 26274 17380 26278 17436
rect 26278 17380 26334 17436
rect 26334 17380 26338 17436
rect 26274 17376 26338 17380
rect 26354 17436 26418 17440
rect 26354 17380 26358 17436
rect 26358 17380 26414 17436
rect 26414 17380 26418 17436
rect 26354 17376 26418 17380
rect 26434 17436 26498 17440
rect 26434 17380 26438 17436
rect 26438 17380 26494 17436
rect 26494 17380 26498 17436
rect 26434 17376 26498 17380
rect 26514 17436 26578 17440
rect 26514 17380 26518 17436
rect 26518 17380 26574 17436
rect 26574 17380 26578 17436
rect 26514 17376 26578 17380
rect 34715 17436 34779 17440
rect 34715 17380 34719 17436
rect 34719 17380 34775 17436
rect 34775 17380 34779 17436
rect 34715 17376 34779 17380
rect 34795 17436 34859 17440
rect 34795 17380 34799 17436
rect 34799 17380 34855 17436
rect 34855 17380 34859 17436
rect 34795 17376 34859 17380
rect 34875 17436 34939 17440
rect 34875 17380 34879 17436
rect 34879 17380 34935 17436
rect 34935 17380 34939 17436
rect 34875 17376 34939 17380
rect 34955 17436 35019 17440
rect 34955 17380 34959 17436
rect 34959 17380 35015 17436
rect 35015 17380 35019 17436
rect 34955 17376 35019 17380
rect 5172 16892 5236 16896
rect 5172 16836 5176 16892
rect 5176 16836 5232 16892
rect 5232 16836 5236 16892
rect 5172 16832 5236 16836
rect 5252 16892 5316 16896
rect 5252 16836 5256 16892
rect 5256 16836 5312 16892
rect 5312 16836 5316 16892
rect 5252 16832 5316 16836
rect 5332 16892 5396 16896
rect 5332 16836 5336 16892
rect 5336 16836 5392 16892
rect 5392 16836 5396 16892
rect 5332 16832 5396 16836
rect 5412 16892 5476 16896
rect 5412 16836 5416 16892
rect 5416 16836 5472 16892
rect 5472 16836 5476 16892
rect 5412 16832 5476 16836
rect 13613 16892 13677 16896
rect 13613 16836 13617 16892
rect 13617 16836 13673 16892
rect 13673 16836 13677 16892
rect 13613 16832 13677 16836
rect 13693 16892 13757 16896
rect 13693 16836 13697 16892
rect 13697 16836 13753 16892
rect 13753 16836 13757 16892
rect 13693 16832 13757 16836
rect 13773 16892 13837 16896
rect 13773 16836 13777 16892
rect 13777 16836 13833 16892
rect 13833 16836 13837 16892
rect 13773 16832 13837 16836
rect 13853 16892 13917 16896
rect 13853 16836 13857 16892
rect 13857 16836 13913 16892
rect 13913 16836 13917 16892
rect 13853 16832 13917 16836
rect 22054 16892 22118 16896
rect 22054 16836 22058 16892
rect 22058 16836 22114 16892
rect 22114 16836 22118 16892
rect 22054 16832 22118 16836
rect 22134 16892 22198 16896
rect 22134 16836 22138 16892
rect 22138 16836 22194 16892
rect 22194 16836 22198 16892
rect 22134 16832 22198 16836
rect 22214 16892 22278 16896
rect 22214 16836 22218 16892
rect 22218 16836 22274 16892
rect 22274 16836 22278 16892
rect 22214 16832 22278 16836
rect 22294 16892 22358 16896
rect 22294 16836 22298 16892
rect 22298 16836 22354 16892
rect 22354 16836 22358 16892
rect 22294 16832 22358 16836
rect 30495 16892 30559 16896
rect 30495 16836 30499 16892
rect 30499 16836 30555 16892
rect 30555 16836 30559 16892
rect 30495 16832 30559 16836
rect 30575 16892 30639 16896
rect 30575 16836 30579 16892
rect 30579 16836 30635 16892
rect 30635 16836 30639 16892
rect 30575 16832 30639 16836
rect 30655 16892 30719 16896
rect 30655 16836 30659 16892
rect 30659 16836 30715 16892
rect 30715 16836 30719 16892
rect 30655 16832 30719 16836
rect 30735 16892 30799 16896
rect 30735 16836 30739 16892
rect 30739 16836 30795 16892
rect 30795 16836 30799 16892
rect 30735 16832 30799 16836
rect 9392 16348 9456 16352
rect 9392 16292 9396 16348
rect 9396 16292 9452 16348
rect 9452 16292 9456 16348
rect 9392 16288 9456 16292
rect 9472 16348 9536 16352
rect 9472 16292 9476 16348
rect 9476 16292 9532 16348
rect 9532 16292 9536 16348
rect 9472 16288 9536 16292
rect 9552 16348 9616 16352
rect 9552 16292 9556 16348
rect 9556 16292 9612 16348
rect 9612 16292 9616 16348
rect 9552 16288 9616 16292
rect 9632 16348 9696 16352
rect 9632 16292 9636 16348
rect 9636 16292 9692 16348
rect 9692 16292 9696 16348
rect 9632 16288 9696 16292
rect 17833 16348 17897 16352
rect 17833 16292 17837 16348
rect 17837 16292 17893 16348
rect 17893 16292 17897 16348
rect 17833 16288 17897 16292
rect 17913 16348 17977 16352
rect 17913 16292 17917 16348
rect 17917 16292 17973 16348
rect 17973 16292 17977 16348
rect 17913 16288 17977 16292
rect 17993 16348 18057 16352
rect 17993 16292 17997 16348
rect 17997 16292 18053 16348
rect 18053 16292 18057 16348
rect 17993 16288 18057 16292
rect 18073 16348 18137 16352
rect 18073 16292 18077 16348
rect 18077 16292 18133 16348
rect 18133 16292 18137 16348
rect 18073 16288 18137 16292
rect 26274 16348 26338 16352
rect 26274 16292 26278 16348
rect 26278 16292 26334 16348
rect 26334 16292 26338 16348
rect 26274 16288 26338 16292
rect 26354 16348 26418 16352
rect 26354 16292 26358 16348
rect 26358 16292 26414 16348
rect 26414 16292 26418 16348
rect 26354 16288 26418 16292
rect 26434 16348 26498 16352
rect 26434 16292 26438 16348
rect 26438 16292 26494 16348
rect 26494 16292 26498 16348
rect 26434 16288 26498 16292
rect 26514 16348 26578 16352
rect 26514 16292 26518 16348
rect 26518 16292 26574 16348
rect 26574 16292 26578 16348
rect 26514 16288 26578 16292
rect 34715 16348 34779 16352
rect 34715 16292 34719 16348
rect 34719 16292 34775 16348
rect 34775 16292 34779 16348
rect 34715 16288 34779 16292
rect 34795 16348 34859 16352
rect 34795 16292 34799 16348
rect 34799 16292 34855 16348
rect 34855 16292 34859 16348
rect 34795 16288 34859 16292
rect 34875 16348 34939 16352
rect 34875 16292 34879 16348
rect 34879 16292 34935 16348
rect 34935 16292 34939 16348
rect 34875 16288 34939 16292
rect 34955 16348 35019 16352
rect 34955 16292 34959 16348
rect 34959 16292 35015 16348
rect 35015 16292 35019 16348
rect 34955 16288 35019 16292
rect 5172 15804 5236 15808
rect 5172 15748 5176 15804
rect 5176 15748 5232 15804
rect 5232 15748 5236 15804
rect 5172 15744 5236 15748
rect 5252 15804 5316 15808
rect 5252 15748 5256 15804
rect 5256 15748 5312 15804
rect 5312 15748 5316 15804
rect 5252 15744 5316 15748
rect 5332 15804 5396 15808
rect 5332 15748 5336 15804
rect 5336 15748 5392 15804
rect 5392 15748 5396 15804
rect 5332 15744 5396 15748
rect 5412 15804 5476 15808
rect 5412 15748 5416 15804
rect 5416 15748 5472 15804
rect 5472 15748 5476 15804
rect 5412 15744 5476 15748
rect 13613 15804 13677 15808
rect 13613 15748 13617 15804
rect 13617 15748 13673 15804
rect 13673 15748 13677 15804
rect 13613 15744 13677 15748
rect 13693 15804 13757 15808
rect 13693 15748 13697 15804
rect 13697 15748 13753 15804
rect 13753 15748 13757 15804
rect 13693 15744 13757 15748
rect 13773 15804 13837 15808
rect 13773 15748 13777 15804
rect 13777 15748 13833 15804
rect 13833 15748 13837 15804
rect 13773 15744 13837 15748
rect 13853 15804 13917 15808
rect 13853 15748 13857 15804
rect 13857 15748 13913 15804
rect 13913 15748 13917 15804
rect 13853 15744 13917 15748
rect 22054 15804 22118 15808
rect 22054 15748 22058 15804
rect 22058 15748 22114 15804
rect 22114 15748 22118 15804
rect 22054 15744 22118 15748
rect 22134 15804 22198 15808
rect 22134 15748 22138 15804
rect 22138 15748 22194 15804
rect 22194 15748 22198 15804
rect 22134 15744 22198 15748
rect 22214 15804 22278 15808
rect 22214 15748 22218 15804
rect 22218 15748 22274 15804
rect 22274 15748 22278 15804
rect 22214 15744 22278 15748
rect 22294 15804 22358 15808
rect 22294 15748 22298 15804
rect 22298 15748 22354 15804
rect 22354 15748 22358 15804
rect 22294 15744 22358 15748
rect 30495 15804 30559 15808
rect 30495 15748 30499 15804
rect 30499 15748 30555 15804
rect 30555 15748 30559 15804
rect 30495 15744 30559 15748
rect 30575 15804 30639 15808
rect 30575 15748 30579 15804
rect 30579 15748 30635 15804
rect 30635 15748 30639 15804
rect 30575 15744 30639 15748
rect 30655 15804 30719 15808
rect 30655 15748 30659 15804
rect 30659 15748 30715 15804
rect 30715 15748 30719 15804
rect 30655 15744 30719 15748
rect 30735 15804 30799 15808
rect 30735 15748 30739 15804
rect 30739 15748 30795 15804
rect 30795 15748 30799 15804
rect 30735 15744 30799 15748
rect 9392 15260 9456 15264
rect 9392 15204 9396 15260
rect 9396 15204 9452 15260
rect 9452 15204 9456 15260
rect 9392 15200 9456 15204
rect 9472 15260 9536 15264
rect 9472 15204 9476 15260
rect 9476 15204 9532 15260
rect 9532 15204 9536 15260
rect 9472 15200 9536 15204
rect 9552 15260 9616 15264
rect 9552 15204 9556 15260
rect 9556 15204 9612 15260
rect 9612 15204 9616 15260
rect 9552 15200 9616 15204
rect 9632 15260 9696 15264
rect 9632 15204 9636 15260
rect 9636 15204 9692 15260
rect 9692 15204 9696 15260
rect 9632 15200 9696 15204
rect 17833 15260 17897 15264
rect 17833 15204 17837 15260
rect 17837 15204 17893 15260
rect 17893 15204 17897 15260
rect 17833 15200 17897 15204
rect 17913 15260 17977 15264
rect 17913 15204 17917 15260
rect 17917 15204 17973 15260
rect 17973 15204 17977 15260
rect 17913 15200 17977 15204
rect 17993 15260 18057 15264
rect 17993 15204 17997 15260
rect 17997 15204 18053 15260
rect 18053 15204 18057 15260
rect 17993 15200 18057 15204
rect 18073 15260 18137 15264
rect 18073 15204 18077 15260
rect 18077 15204 18133 15260
rect 18133 15204 18137 15260
rect 18073 15200 18137 15204
rect 26274 15260 26338 15264
rect 26274 15204 26278 15260
rect 26278 15204 26334 15260
rect 26334 15204 26338 15260
rect 26274 15200 26338 15204
rect 26354 15260 26418 15264
rect 26354 15204 26358 15260
rect 26358 15204 26414 15260
rect 26414 15204 26418 15260
rect 26354 15200 26418 15204
rect 26434 15260 26498 15264
rect 26434 15204 26438 15260
rect 26438 15204 26494 15260
rect 26494 15204 26498 15260
rect 26434 15200 26498 15204
rect 26514 15260 26578 15264
rect 26514 15204 26518 15260
rect 26518 15204 26574 15260
rect 26574 15204 26578 15260
rect 26514 15200 26578 15204
rect 34715 15260 34779 15264
rect 34715 15204 34719 15260
rect 34719 15204 34775 15260
rect 34775 15204 34779 15260
rect 34715 15200 34779 15204
rect 34795 15260 34859 15264
rect 34795 15204 34799 15260
rect 34799 15204 34855 15260
rect 34855 15204 34859 15260
rect 34795 15200 34859 15204
rect 34875 15260 34939 15264
rect 34875 15204 34879 15260
rect 34879 15204 34935 15260
rect 34935 15204 34939 15260
rect 34875 15200 34939 15204
rect 34955 15260 35019 15264
rect 34955 15204 34959 15260
rect 34959 15204 35015 15260
rect 35015 15204 35019 15260
rect 34955 15200 35019 15204
rect 5172 14716 5236 14720
rect 5172 14660 5176 14716
rect 5176 14660 5232 14716
rect 5232 14660 5236 14716
rect 5172 14656 5236 14660
rect 5252 14716 5316 14720
rect 5252 14660 5256 14716
rect 5256 14660 5312 14716
rect 5312 14660 5316 14716
rect 5252 14656 5316 14660
rect 5332 14716 5396 14720
rect 5332 14660 5336 14716
rect 5336 14660 5392 14716
rect 5392 14660 5396 14716
rect 5332 14656 5396 14660
rect 5412 14716 5476 14720
rect 5412 14660 5416 14716
rect 5416 14660 5472 14716
rect 5472 14660 5476 14716
rect 5412 14656 5476 14660
rect 13613 14716 13677 14720
rect 13613 14660 13617 14716
rect 13617 14660 13673 14716
rect 13673 14660 13677 14716
rect 13613 14656 13677 14660
rect 13693 14716 13757 14720
rect 13693 14660 13697 14716
rect 13697 14660 13753 14716
rect 13753 14660 13757 14716
rect 13693 14656 13757 14660
rect 13773 14716 13837 14720
rect 13773 14660 13777 14716
rect 13777 14660 13833 14716
rect 13833 14660 13837 14716
rect 13773 14656 13837 14660
rect 13853 14716 13917 14720
rect 13853 14660 13857 14716
rect 13857 14660 13913 14716
rect 13913 14660 13917 14716
rect 13853 14656 13917 14660
rect 22054 14716 22118 14720
rect 22054 14660 22058 14716
rect 22058 14660 22114 14716
rect 22114 14660 22118 14716
rect 22054 14656 22118 14660
rect 22134 14716 22198 14720
rect 22134 14660 22138 14716
rect 22138 14660 22194 14716
rect 22194 14660 22198 14716
rect 22134 14656 22198 14660
rect 22214 14716 22278 14720
rect 22214 14660 22218 14716
rect 22218 14660 22274 14716
rect 22274 14660 22278 14716
rect 22214 14656 22278 14660
rect 22294 14716 22358 14720
rect 22294 14660 22298 14716
rect 22298 14660 22354 14716
rect 22354 14660 22358 14716
rect 22294 14656 22358 14660
rect 30495 14716 30559 14720
rect 30495 14660 30499 14716
rect 30499 14660 30555 14716
rect 30555 14660 30559 14716
rect 30495 14656 30559 14660
rect 30575 14716 30639 14720
rect 30575 14660 30579 14716
rect 30579 14660 30635 14716
rect 30635 14660 30639 14716
rect 30575 14656 30639 14660
rect 30655 14716 30719 14720
rect 30655 14660 30659 14716
rect 30659 14660 30715 14716
rect 30715 14660 30719 14716
rect 30655 14656 30719 14660
rect 30735 14716 30799 14720
rect 30735 14660 30739 14716
rect 30739 14660 30795 14716
rect 30795 14660 30799 14716
rect 30735 14656 30799 14660
rect 9392 14172 9456 14176
rect 9392 14116 9396 14172
rect 9396 14116 9452 14172
rect 9452 14116 9456 14172
rect 9392 14112 9456 14116
rect 9472 14172 9536 14176
rect 9472 14116 9476 14172
rect 9476 14116 9532 14172
rect 9532 14116 9536 14172
rect 9472 14112 9536 14116
rect 9552 14172 9616 14176
rect 9552 14116 9556 14172
rect 9556 14116 9612 14172
rect 9612 14116 9616 14172
rect 9552 14112 9616 14116
rect 9632 14172 9696 14176
rect 9632 14116 9636 14172
rect 9636 14116 9692 14172
rect 9692 14116 9696 14172
rect 9632 14112 9696 14116
rect 17833 14172 17897 14176
rect 17833 14116 17837 14172
rect 17837 14116 17893 14172
rect 17893 14116 17897 14172
rect 17833 14112 17897 14116
rect 17913 14172 17977 14176
rect 17913 14116 17917 14172
rect 17917 14116 17973 14172
rect 17973 14116 17977 14172
rect 17913 14112 17977 14116
rect 17993 14172 18057 14176
rect 17993 14116 17997 14172
rect 17997 14116 18053 14172
rect 18053 14116 18057 14172
rect 17993 14112 18057 14116
rect 18073 14172 18137 14176
rect 18073 14116 18077 14172
rect 18077 14116 18133 14172
rect 18133 14116 18137 14172
rect 18073 14112 18137 14116
rect 26274 14172 26338 14176
rect 26274 14116 26278 14172
rect 26278 14116 26334 14172
rect 26334 14116 26338 14172
rect 26274 14112 26338 14116
rect 26354 14172 26418 14176
rect 26354 14116 26358 14172
rect 26358 14116 26414 14172
rect 26414 14116 26418 14172
rect 26354 14112 26418 14116
rect 26434 14172 26498 14176
rect 26434 14116 26438 14172
rect 26438 14116 26494 14172
rect 26494 14116 26498 14172
rect 26434 14112 26498 14116
rect 26514 14172 26578 14176
rect 26514 14116 26518 14172
rect 26518 14116 26574 14172
rect 26574 14116 26578 14172
rect 26514 14112 26578 14116
rect 34715 14172 34779 14176
rect 34715 14116 34719 14172
rect 34719 14116 34775 14172
rect 34775 14116 34779 14172
rect 34715 14112 34779 14116
rect 34795 14172 34859 14176
rect 34795 14116 34799 14172
rect 34799 14116 34855 14172
rect 34855 14116 34859 14172
rect 34795 14112 34859 14116
rect 34875 14172 34939 14176
rect 34875 14116 34879 14172
rect 34879 14116 34935 14172
rect 34935 14116 34939 14172
rect 34875 14112 34939 14116
rect 34955 14172 35019 14176
rect 34955 14116 34959 14172
rect 34959 14116 35015 14172
rect 35015 14116 35019 14172
rect 34955 14112 35019 14116
rect 5172 13628 5236 13632
rect 5172 13572 5176 13628
rect 5176 13572 5232 13628
rect 5232 13572 5236 13628
rect 5172 13568 5236 13572
rect 5252 13628 5316 13632
rect 5252 13572 5256 13628
rect 5256 13572 5312 13628
rect 5312 13572 5316 13628
rect 5252 13568 5316 13572
rect 5332 13628 5396 13632
rect 5332 13572 5336 13628
rect 5336 13572 5392 13628
rect 5392 13572 5396 13628
rect 5332 13568 5396 13572
rect 5412 13628 5476 13632
rect 5412 13572 5416 13628
rect 5416 13572 5472 13628
rect 5472 13572 5476 13628
rect 5412 13568 5476 13572
rect 13613 13628 13677 13632
rect 13613 13572 13617 13628
rect 13617 13572 13673 13628
rect 13673 13572 13677 13628
rect 13613 13568 13677 13572
rect 13693 13628 13757 13632
rect 13693 13572 13697 13628
rect 13697 13572 13753 13628
rect 13753 13572 13757 13628
rect 13693 13568 13757 13572
rect 13773 13628 13837 13632
rect 13773 13572 13777 13628
rect 13777 13572 13833 13628
rect 13833 13572 13837 13628
rect 13773 13568 13837 13572
rect 13853 13628 13917 13632
rect 13853 13572 13857 13628
rect 13857 13572 13913 13628
rect 13913 13572 13917 13628
rect 13853 13568 13917 13572
rect 22054 13628 22118 13632
rect 22054 13572 22058 13628
rect 22058 13572 22114 13628
rect 22114 13572 22118 13628
rect 22054 13568 22118 13572
rect 22134 13628 22198 13632
rect 22134 13572 22138 13628
rect 22138 13572 22194 13628
rect 22194 13572 22198 13628
rect 22134 13568 22198 13572
rect 22214 13628 22278 13632
rect 22214 13572 22218 13628
rect 22218 13572 22274 13628
rect 22274 13572 22278 13628
rect 22214 13568 22278 13572
rect 22294 13628 22358 13632
rect 22294 13572 22298 13628
rect 22298 13572 22354 13628
rect 22354 13572 22358 13628
rect 22294 13568 22358 13572
rect 30495 13628 30559 13632
rect 30495 13572 30499 13628
rect 30499 13572 30555 13628
rect 30555 13572 30559 13628
rect 30495 13568 30559 13572
rect 30575 13628 30639 13632
rect 30575 13572 30579 13628
rect 30579 13572 30635 13628
rect 30635 13572 30639 13628
rect 30575 13568 30639 13572
rect 30655 13628 30719 13632
rect 30655 13572 30659 13628
rect 30659 13572 30715 13628
rect 30715 13572 30719 13628
rect 30655 13568 30719 13572
rect 30735 13628 30799 13632
rect 30735 13572 30739 13628
rect 30739 13572 30795 13628
rect 30795 13572 30799 13628
rect 30735 13568 30799 13572
rect 9392 13084 9456 13088
rect 9392 13028 9396 13084
rect 9396 13028 9452 13084
rect 9452 13028 9456 13084
rect 9392 13024 9456 13028
rect 9472 13084 9536 13088
rect 9472 13028 9476 13084
rect 9476 13028 9532 13084
rect 9532 13028 9536 13084
rect 9472 13024 9536 13028
rect 9552 13084 9616 13088
rect 9552 13028 9556 13084
rect 9556 13028 9612 13084
rect 9612 13028 9616 13084
rect 9552 13024 9616 13028
rect 9632 13084 9696 13088
rect 9632 13028 9636 13084
rect 9636 13028 9692 13084
rect 9692 13028 9696 13084
rect 9632 13024 9696 13028
rect 17833 13084 17897 13088
rect 17833 13028 17837 13084
rect 17837 13028 17893 13084
rect 17893 13028 17897 13084
rect 17833 13024 17897 13028
rect 17913 13084 17977 13088
rect 17913 13028 17917 13084
rect 17917 13028 17973 13084
rect 17973 13028 17977 13084
rect 17913 13024 17977 13028
rect 17993 13084 18057 13088
rect 17993 13028 17997 13084
rect 17997 13028 18053 13084
rect 18053 13028 18057 13084
rect 17993 13024 18057 13028
rect 18073 13084 18137 13088
rect 18073 13028 18077 13084
rect 18077 13028 18133 13084
rect 18133 13028 18137 13084
rect 18073 13024 18137 13028
rect 26274 13084 26338 13088
rect 26274 13028 26278 13084
rect 26278 13028 26334 13084
rect 26334 13028 26338 13084
rect 26274 13024 26338 13028
rect 26354 13084 26418 13088
rect 26354 13028 26358 13084
rect 26358 13028 26414 13084
rect 26414 13028 26418 13084
rect 26354 13024 26418 13028
rect 26434 13084 26498 13088
rect 26434 13028 26438 13084
rect 26438 13028 26494 13084
rect 26494 13028 26498 13084
rect 26434 13024 26498 13028
rect 26514 13084 26578 13088
rect 26514 13028 26518 13084
rect 26518 13028 26574 13084
rect 26574 13028 26578 13084
rect 26514 13024 26578 13028
rect 34715 13084 34779 13088
rect 34715 13028 34719 13084
rect 34719 13028 34775 13084
rect 34775 13028 34779 13084
rect 34715 13024 34779 13028
rect 34795 13084 34859 13088
rect 34795 13028 34799 13084
rect 34799 13028 34855 13084
rect 34855 13028 34859 13084
rect 34795 13024 34859 13028
rect 34875 13084 34939 13088
rect 34875 13028 34879 13084
rect 34879 13028 34935 13084
rect 34935 13028 34939 13084
rect 34875 13024 34939 13028
rect 34955 13084 35019 13088
rect 34955 13028 34959 13084
rect 34959 13028 35015 13084
rect 35015 13028 35019 13084
rect 34955 13024 35019 13028
rect 5172 12540 5236 12544
rect 5172 12484 5176 12540
rect 5176 12484 5232 12540
rect 5232 12484 5236 12540
rect 5172 12480 5236 12484
rect 5252 12540 5316 12544
rect 5252 12484 5256 12540
rect 5256 12484 5312 12540
rect 5312 12484 5316 12540
rect 5252 12480 5316 12484
rect 5332 12540 5396 12544
rect 5332 12484 5336 12540
rect 5336 12484 5392 12540
rect 5392 12484 5396 12540
rect 5332 12480 5396 12484
rect 5412 12540 5476 12544
rect 5412 12484 5416 12540
rect 5416 12484 5472 12540
rect 5472 12484 5476 12540
rect 5412 12480 5476 12484
rect 13613 12540 13677 12544
rect 13613 12484 13617 12540
rect 13617 12484 13673 12540
rect 13673 12484 13677 12540
rect 13613 12480 13677 12484
rect 13693 12540 13757 12544
rect 13693 12484 13697 12540
rect 13697 12484 13753 12540
rect 13753 12484 13757 12540
rect 13693 12480 13757 12484
rect 13773 12540 13837 12544
rect 13773 12484 13777 12540
rect 13777 12484 13833 12540
rect 13833 12484 13837 12540
rect 13773 12480 13837 12484
rect 13853 12540 13917 12544
rect 13853 12484 13857 12540
rect 13857 12484 13913 12540
rect 13913 12484 13917 12540
rect 13853 12480 13917 12484
rect 22054 12540 22118 12544
rect 22054 12484 22058 12540
rect 22058 12484 22114 12540
rect 22114 12484 22118 12540
rect 22054 12480 22118 12484
rect 22134 12540 22198 12544
rect 22134 12484 22138 12540
rect 22138 12484 22194 12540
rect 22194 12484 22198 12540
rect 22134 12480 22198 12484
rect 22214 12540 22278 12544
rect 22214 12484 22218 12540
rect 22218 12484 22274 12540
rect 22274 12484 22278 12540
rect 22214 12480 22278 12484
rect 22294 12540 22358 12544
rect 22294 12484 22298 12540
rect 22298 12484 22354 12540
rect 22354 12484 22358 12540
rect 22294 12480 22358 12484
rect 30495 12540 30559 12544
rect 30495 12484 30499 12540
rect 30499 12484 30555 12540
rect 30555 12484 30559 12540
rect 30495 12480 30559 12484
rect 30575 12540 30639 12544
rect 30575 12484 30579 12540
rect 30579 12484 30635 12540
rect 30635 12484 30639 12540
rect 30575 12480 30639 12484
rect 30655 12540 30719 12544
rect 30655 12484 30659 12540
rect 30659 12484 30715 12540
rect 30715 12484 30719 12540
rect 30655 12480 30719 12484
rect 30735 12540 30799 12544
rect 30735 12484 30739 12540
rect 30739 12484 30795 12540
rect 30795 12484 30799 12540
rect 30735 12480 30799 12484
rect 9392 11996 9456 12000
rect 9392 11940 9396 11996
rect 9396 11940 9452 11996
rect 9452 11940 9456 11996
rect 9392 11936 9456 11940
rect 9472 11996 9536 12000
rect 9472 11940 9476 11996
rect 9476 11940 9532 11996
rect 9532 11940 9536 11996
rect 9472 11936 9536 11940
rect 9552 11996 9616 12000
rect 9552 11940 9556 11996
rect 9556 11940 9612 11996
rect 9612 11940 9616 11996
rect 9552 11936 9616 11940
rect 9632 11996 9696 12000
rect 9632 11940 9636 11996
rect 9636 11940 9692 11996
rect 9692 11940 9696 11996
rect 9632 11936 9696 11940
rect 17833 11996 17897 12000
rect 17833 11940 17837 11996
rect 17837 11940 17893 11996
rect 17893 11940 17897 11996
rect 17833 11936 17897 11940
rect 17913 11996 17977 12000
rect 17913 11940 17917 11996
rect 17917 11940 17973 11996
rect 17973 11940 17977 11996
rect 17913 11936 17977 11940
rect 17993 11996 18057 12000
rect 17993 11940 17997 11996
rect 17997 11940 18053 11996
rect 18053 11940 18057 11996
rect 17993 11936 18057 11940
rect 18073 11996 18137 12000
rect 18073 11940 18077 11996
rect 18077 11940 18133 11996
rect 18133 11940 18137 11996
rect 18073 11936 18137 11940
rect 26274 11996 26338 12000
rect 26274 11940 26278 11996
rect 26278 11940 26334 11996
rect 26334 11940 26338 11996
rect 26274 11936 26338 11940
rect 26354 11996 26418 12000
rect 26354 11940 26358 11996
rect 26358 11940 26414 11996
rect 26414 11940 26418 11996
rect 26354 11936 26418 11940
rect 26434 11996 26498 12000
rect 26434 11940 26438 11996
rect 26438 11940 26494 11996
rect 26494 11940 26498 11996
rect 26434 11936 26498 11940
rect 26514 11996 26578 12000
rect 26514 11940 26518 11996
rect 26518 11940 26574 11996
rect 26574 11940 26578 11996
rect 26514 11936 26578 11940
rect 34715 11996 34779 12000
rect 34715 11940 34719 11996
rect 34719 11940 34775 11996
rect 34775 11940 34779 11996
rect 34715 11936 34779 11940
rect 34795 11996 34859 12000
rect 34795 11940 34799 11996
rect 34799 11940 34855 11996
rect 34855 11940 34859 11996
rect 34795 11936 34859 11940
rect 34875 11996 34939 12000
rect 34875 11940 34879 11996
rect 34879 11940 34935 11996
rect 34935 11940 34939 11996
rect 34875 11936 34939 11940
rect 34955 11996 35019 12000
rect 34955 11940 34959 11996
rect 34959 11940 35015 11996
rect 35015 11940 35019 11996
rect 34955 11936 35019 11940
rect 5172 11452 5236 11456
rect 5172 11396 5176 11452
rect 5176 11396 5232 11452
rect 5232 11396 5236 11452
rect 5172 11392 5236 11396
rect 5252 11452 5316 11456
rect 5252 11396 5256 11452
rect 5256 11396 5312 11452
rect 5312 11396 5316 11452
rect 5252 11392 5316 11396
rect 5332 11452 5396 11456
rect 5332 11396 5336 11452
rect 5336 11396 5392 11452
rect 5392 11396 5396 11452
rect 5332 11392 5396 11396
rect 5412 11452 5476 11456
rect 5412 11396 5416 11452
rect 5416 11396 5472 11452
rect 5472 11396 5476 11452
rect 5412 11392 5476 11396
rect 13613 11452 13677 11456
rect 13613 11396 13617 11452
rect 13617 11396 13673 11452
rect 13673 11396 13677 11452
rect 13613 11392 13677 11396
rect 13693 11452 13757 11456
rect 13693 11396 13697 11452
rect 13697 11396 13753 11452
rect 13753 11396 13757 11452
rect 13693 11392 13757 11396
rect 13773 11452 13837 11456
rect 13773 11396 13777 11452
rect 13777 11396 13833 11452
rect 13833 11396 13837 11452
rect 13773 11392 13837 11396
rect 13853 11452 13917 11456
rect 13853 11396 13857 11452
rect 13857 11396 13913 11452
rect 13913 11396 13917 11452
rect 13853 11392 13917 11396
rect 22054 11452 22118 11456
rect 22054 11396 22058 11452
rect 22058 11396 22114 11452
rect 22114 11396 22118 11452
rect 22054 11392 22118 11396
rect 22134 11452 22198 11456
rect 22134 11396 22138 11452
rect 22138 11396 22194 11452
rect 22194 11396 22198 11452
rect 22134 11392 22198 11396
rect 22214 11452 22278 11456
rect 22214 11396 22218 11452
rect 22218 11396 22274 11452
rect 22274 11396 22278 11452
rect 22214 11392 22278 11396
rect 22294 11452 22358 11456
rect 22294 11396 22298 11452
rect 22298 11396 22354 11452
rect 22354 11396 22358 11452
rect 22294 11392 22358 11396
rect 30495 11452 30559 11456
rect 30495 11396 30499 11452
rect 30499 11396 30555 11452
rect 30555 11396 30559 11452
rect 30495 11392 30559 11396
rect 30575 11452 30639 11456
rect 30575 11396 30579 11452
rect 30579 11396 30635 11452
rect 30635 11396 30639 11452
rect 30575 11392 30639 11396
rect 30655 11452 30719 11456
rect 30655 11396 30659 11452
rect 30659 11396 30715 11452
rect 30715 11396 30719 11452
rect 30655 11392 30719 11396
rect 30735 11452 30799 11456
rect 30735 11396 30739 11452
rect 30739 11396 30795 11452
rect 30795 11396 30799 11452
rect 30735 11392 30799 11396
rect 9392 10908 9456 10912
rect 9392 10852 9396 10908
rect 9396 10852 9452 10908
rect 9452 10852 9456 10908
rect 9392 10848 9456 10852
rect 9472 10908 9536 10912
rect 9472 10852 9476 10908
rect 9476 10852 9532 10908
rect 9532 10852 9536 10908
rect 9472 10848 9536 10852
rect 9552 10908 9616 10912
rect 9552 10852 9556 10908
rect 9556 10852 9612 10908
rect 9612 10852 9616 10908
rect 9552 10848 9616 10852
rect 9632 10908 9696 10912
rect 9632 10852 9636 10908
rect 9636 10852 9692 10908
rect 9692 10852 9696 10908
rect 9632 10848 9696 10852
rect 17833 10908 17897 10912
rect 17833 10852 17837 10908
rect 17837 10852 17893 10908
rect 17893 10852 17897 10908
rect 17833 10848 17897 10852
rect 17913 10908 17977 10912
rect 17913 10852 17917 10908
rect 17917 10852 17973 10908
rect 17973 10852 17977 10908
rect 17913 10848 17977 10852
rect 17993 10908 18057 10912
rect 17993 10852 17997 10908
rect 17997 10852 18053 10908
rect 18053 10852 18057 10908
rect 17993 10848 18057 10852
rect 18073 10908 18137 10912
rect 18073 10852 18077 10908
rect 18077 10852 18133 10908
rect 18133 10852 18137 10908
rect 18073 10848 18137 10852
rect 26274 10908 26338 10912
rect 26274 10852 26278 10908
rect 26278 10852 26334 10908
rect 26334 10852 26338 10908
rect 26274 10848 26338 10852
rect 26354 10908 26418 10912
rect 26354 10852 26358 10908
rect 26358 10852 26414 10908
rect 26414 10852 26418 10908
rect 26354 10848 26418 10852
rect 26434 10908 26498 10912
rect 26434 10852 26438 10908
rect 26438 10852 26494 10908
rect 26494 10852 26498 10908
rect 26434 10848 26498 10852
rect 26514 10908 26578 10912
rect 26514 10852 26518 10908
rect 26518 10852 26574 10908
rect 26574 10852 26578 10908
rect 26514 10848 26578 10852
rect 34715 10908 34779 10912
rect 34715 10852 34719 10908
rect 34719 10852 34775 10908
rect 34775 10852 34779 10908
rect 34715 10848 34779 10852
rect 34795 10908 34859 10912
rect 34795 10852 34799 10908
rect 34799 10852 34855 10908
rect 34855 10852 34859 10908
rect 34795 10848 34859 10852
rect 34875 10908 34939 10912
rect 34875 10852 34879 10908
rect 34879 10852 34935 10908
rect 34935 10852 34939 10908
rect 34875 10848 34939 10852
rect 34955 10908 35019 10912
rect 34955 10852 34959 10908
rect 34959 10852 35015 10908
rect 35015 10852 35019 10908
rect 34955 10848 35019 10852
rect 5172 10364 5236 10368
rect 5172 10308 5176 10364
rect 5176 10308 5232 10364
rect 5232 10308 5236 10364
rect 5172 10304 5236 10308
rect 5252 10364 5316 10368
rect 5252 10308 5256 10364
rect 5256 10308 5312 10364
rect 5312 10308 5316 10364
rect 5252 10304 5316 10308
rect 5332 10364 5396 10368
rect 5332 10308 5336 10364
rect 5336 10308 5392 10364
rect 5392 10308 5396 10364
rect 5332 10304 5396 10308
rect 5412 10364 5476 10368
rect 5412 10308 5416 10364
rect 5416 10308 5472 10364
rect 5472 10308 5476 10364
rect 5412 10304 5476 10308
rect 13613 10364 13677 10368
rect 13613 10308 13617 10364
rect 13617 10308 13673 10364
rect 13673 10308 13677 10364
rect 13613 10304 13677 10308
rect 13693 10364 13757 10368
rect 13693 10308 13697 10364
rect 13697 10308 13753 10364
rect 13753 10308 13757 10364
rect 13693 10304 13757 10308
rect 13773 10364 13837 10368
rect 13773 10308 13777 10364
rect 13777 10308 13833 10364
rect 13833 10308 13837 10364
rect 13773 10304 13837 10308
rect 13853 10364 13917 10368
rect 13853 10308 13857 10364
rect 13857 10308 13913 10364
rect 13913 10308 13917 10364
rect 13853 10304 13917 10308
rect 22054 10364 22118 10368
rect 22054 10308 22058 10364
rect 22058 10308 22114 10364
rect 22114 10308 22118 10364
rect 22054 10304 22118 10308
rect 22134 10364 22198 10368
rect 22134 10308 22138 10364
rect 22138 10308 22194 10364
rect 22194 10308 22198 10364
rect 22134 10304 22198 10308
rect 22214 10364 22278 10368
rect 22214 10308 22218 10364
rect 22218 10308 22274 10364
rect 22274 10308 22278 10364
rect 22214 10304 22278 10308
rect 22294 10364 22358 10368
rect 22294 10308 22298 10364
rect 22298 10308 22354 10364
rect 22354 10308 22358 10364
rect 22294 10304 22358 10308
rect 30495 10364 30559 10368
rect 30495 10308 30499 10364
rect 30499 10308 30555 10364
rect 30555 10308 30559 10364
rect 30495 10304 30559 10308
rect 30575 10364 30639 10368
rect 30575 10308 30579 10364
rect 30579 10308 30635 10364
rect 30635 10308 30639 10364
rect 30575 10304 30639 10308
rect 30655 10364 30719 10368
rect 30655 10308 30659 10364
rect 30659 10308 30715 10364
rect 30715 10308 30719 10364
rect 30655 10304 30719 10308
rect 30735 10364 30799 10368
rect 30735 10308 30739 10364
rect 30739 10308 30795 10364
rect 30795 10308 30799 10364
rect 30735 10304 30799 10308
rect 9392 9820 9456 9824
rect 9392 9764 9396 9820
rect 9396 9764 9452 9820
rect 9452 9764 9456 9820
rect 9392 9760 9456 9764
rect 9472 9820 9536 9824
rect 9472 9764 9476 9820
rect 9476 9764 9532 9820
rect 9532 9764 9536 9820
rect 9472 9760 9536 9764
rect 9552 9820 9616 9824
rect 9552 9764 9556 9820
rect 9556 9764 9612 9820
rect 9612 9764 9616 9820
rect 9552 9760 9616 9764
rect 9632 9820 9696 9824
rect 9632 9764 9636 9820
rect 9636 9764 9692 9820
rect 9692 9764 9696 9820
rect 9632 9760 9696 9764
rect 17833 9820 17897 9824
rect 17833 9764 17837 9820
rect 17837 9764 17893 9820
rect 17893 9764 17897 9820
rect 17833 9760 17897 9764
rect 17913 9820 17977 9824
rect 17913 9764 17917 9820
rect 17917 9764 17973 9820
rect 17973 9764 17977 9820
rect 17913 9760 17977 9764
rect 17993 9820 18057 9824
rect 17993 9764 17997 9820
rect 17997 9764 18053 9820
rect 18053 9764 18057 9820
rect 17993 9760 18057 9764
rect 18073 9820 18137 9824
rect 18073 9764 18077 9820
rect 18077 9764 18133 9820
rect 18133 9764 18137 9820
rect 18073 9760 18137 9764
rect 26274 9820 26338 9824
rect 26274 9764 26278 9820
rect 26278 9764 26334 9820
rect 26334 9764 26338 9820
rect 26274 9760 26338 9764
rect 26354 9820 26418 9824
rect 26354 9764 26358 9820
rect 26358 9764 26414 9820
rect 26414 9764 26418 9820
rect 26354 9760 26418 9764
rect 26434 9820 26498 9824
rect 26434 9764 26438 9820
rect 26438 9764 26494 9820
rect 26494 9764 26498 9820
rect 26434 9760 26498 9764
rect 26514 9820 26578 9824
rect 26514 9764 26518 9820
rect 26518 9764 26574 9820
rect 26574 9764 26578 9820
rect 26514 9760 26578 9764
rect 34715 9820 34779 9824
rect 34715 9764 34719 9820
rect 34719 9764 34775 9820
rect 34775 9764 34779 9820
rect 34715 9760 34779 9764
rect 34795 9820 34859 9824
rect 34795 9764 34799 9820
rect 34799 9764 34855 9820
rect 34855 9764 34859 9820
rect 34795 9760 34859 9764
rect 34875 9820 34939 9824
rect 34875 9764 34879 9820
rect 34879 9764 34935 9820
rect 34935 9764 34939 9820
rect 34875 9760 34939 9764
rect 34955 9820 35019 9824
rect 34955 9764 34959 9820
rect 34959 9764 35015 9820
rect 35015 9764 35019 9820
rect 34955 9760 35019 9764
rect 5172 9276 5236 9280
rect 5172 9220 5176 9276
rect 5176 9220 5232 9276
rect 5232 9220 5236 9276
rect 5172 9216 5236 9220
rect 5252 9276 5316 9280
rect 5252 9220 5256 9276
rect 5256 9220 5312 9276
rect 5312 9220 5316 9276
rect 5252 9216 5316 9220
rect 5332 9276 5396 9280
rect 5332 9220 5336 9276
rect 5336 9220 5392 9276
rect 5392 9220 5396 9276
rect 5332 9216 5396 9220
rect 5412 9276 5476 9280
rect 5412 9220 5416 9276
rect 5416 9220 5472 9276
rect 5472 9220 5476 9276
rect 5412 9216 5476 9220
rect 13613 9276 13677 9280
rect 13613 9220 13617 9276
rect 13617 9220 13673 9276
rect 13673 9220 13677 9276
rect 13613 9216 13677 9220
rect 13693 9276 13757 9280
rect 13693 9220 13697 9276
rect 13697 9220 13753 9276
rect 13753 9220 13757 9276
rect 13693 9216 13757 9220
rect 13773 9276 13837 9280
rect 13773 9220 13777 9276
rect 13777 9220 13833 9276
rect 13833 9220 13837 9276
rect 13773 9216 13837 9220
rect 13853 9276 13917 9280
rect 13853 9220 13857 9276
rect 13857 9220 13913 9276
rect 13913 9220 13917 9276
rect 13853 9216 13917 9220
rect 22054 9276 22118 9280
rect 22054 9220 22058 9276
rect 22058 9220 22114 9276
rect 22114 9220 22118 9276
rect 22054 9216 22118 9220
rect 22134 9276 22198 9280
rect 22134 9220 22138 9276
rect 22138 9220 22194 9276
rect 22194 9220 22198 9276
rect 22134 9216 22198 9220
rect 22214 9276 22278 9280
rect 22214 9220 22218 9276
rect 22218 9220 22274 9276
rect 22274 9220 22278 9276
rect 22214 9216 22278 9220
rect 22294 9276 22358 9280
rect 22294 9220 22298 9276
rect 22298 9220 22354 9276
rect 22354 9220 22358 9276
rect 22294 9216 22358 9220
rect 30495 9276 30559 9280
rect 30495 9220 30499 9276
rect 30499 9220 30555 9276
rect 30555 9220 30559 9276
rect 30495 9216 30559 9220
rect 30575 9276 30639 9280
rect 30575 9220 30579 9276
rect 30579 9220 30635 9276
rect 30635 9220 30639 9276
rect 30575 9216 30639 9220
rect 30655 9276 30719 9280
rect 30655 9220 30659 9276
rect 30659 9220 30715 9276
rect 30715 9220 30719 9276
rect 30655 9216 30719 9220
rect 30735 9276 30799 9280
rect 30735 9220 30739 9276
rect 30739 9220 30795 9276
rect 30795 9220 30799 9276
rect 30735 9216 30799 9220
rect 9392 8732 9456 8736
rect 9392 8676 9396 8732
rect 9396 8676 9452 8732
rect 9452 8676 9456 8732
rect 9392 8672 9456 8676
rect 9472 8732 9536 8736
rect 9472 8676 9476 8732
rect 9476 8676 9532 8732
rect 9532 8676 9536 8732
rect 9472 8672 9536 8676
rect 9552 8732 9616 8736
rect 9552 8676 9556 8732
rect 9556 8676 9612 8732
rect 9612 8676 9616 8732
rect 9552 8672 9616 8676
rect 9632 8732 9696 8736
rect 9632 8676 9636 8732
rect 9636 8676 9692 8732
rect 9692 8676 9696 8732
rect 9632 8672 9696 8676
rect 17833 8732 17897 8736
rect 17833 8676 17837 8732
rect 17837 8676 17893 8732
rect 17893 8676 17897 8732
rect 17833 8672 17897 8676
rect 17913 8732 17977 8736
rect 17913 8676 17917 8732
rect 17917 8676 17973 8732
rect 17973 8676 17977 8732
rect 17913 8672 17977 8676
rect 17993 8732 18057 8736
rect 17993 8676 17997 8732
rect 17997 8676 18053 8732
rect 18053 8676 18057 8732
rect 17993 8672 18057 8676
rect 18073 8732 18137 8736
rect 18073 8676 18077 8732
rect 18077 8676 18133 8732
rect 18133 8676 18137 8732
rect 18073 8672 18137 8676
rect 26274 8732 26338 8736
rect 26274 8676 26278 8732
rect 26278 8676 26334 8732
rect 26334 8676 26338 8732
rect 26274 8672 26338 8676
rect 26354 8732 26418 8736
rect 26354 8676 26358 8732
rect 26358 8676 26414 8732
rect 26414 8676 26418 8732
rect 26354 8672 26418 8676
rect 26434 8732 26498 8736
rect 26434 8676 26438 8732
rect 26438 8676 26494 8732
rect 26494 8676 26498 8732
rect 26434 8672 26498 8676
rect 26514 8732 26578 8736
rect 26514 8676 26518 8732
rect 26518 8676 26574 8732
rect 26574 8676 26578 8732
rect 26514 8672 26578 8676
rect 34715 8732 34779 8736
rect 34715 8676 34719 8732
rect 34719 8676 34775 8732
rect 34775 8676 34779 8732
rect 34715 8672 34779 8676
rect 34795 8732 34859 8736
rect 34795 8676 34799 8732
rect 34799 8676 34855 8732
rect 34855 8676 34859 8732
rect 34795 8672 34859 8676
rect 34875 8732 34939 8736
rect 34875 8676 34879 8732
rect 34879 8676 34935 8732
rect 34935 8676 34939 8732
rect 34875 8672 34939 8676
rect 34955 8732 35019 8736
rect 34955 8676 34959 8732
rect 34959 8676 35015 8732
rect 35015 8676 35019 8732
rect 34955 8672 35019 8676
rect 5172 8188 5236 8192
rect 5172 8132 5176 8188
rect 5176 8132 5232 8188
rect 5232 8132 5236 8188
rect 5172 8128 5236 8132
rect 5252 8188 5316 8192
rect 5252 8132 5256 8188
rect 5256 8132 5312 8188
rect 5312 8132 5316 8188
rect 5252 8128 5316 8132
rect 5332 8188 5396 8192
rect 5332 8132 5336 8188
rect 5336 8132 5392 8188
rect 5392 8132 5396 8188
rect 5332 8128 5396 8132
rect 5412 8188 5476 8192
rect 5412 8132 5416 8188
rect 5416 8132 5472 8188
rect 5472 8132 5476 8188
rect 5412 8128 5476 8132
rect 13613 8188 13677 8192
rect 13613 8132 13617 8188
rect 13617 8132 13673 8188
rect 13673 8132 13677 8188
rect 13613 8128 13677 8132
rect 13693 8188 13757 8192
rect 13693 8132 13697 8188
rect 13697 8132 13753 8188
rect 13753 8132 13757 8188
rect 13693 8128 13757 8132
rect 13773 8188 13837 8192
rect 13773 8132 13777 8188
rect 13777 8132 13833 8188
rect 13833 8132 13837 8188
rect 13773 8128 13837 8132
rect 13853 8188 13917 8192
rect 13853 8132 13857 8188
rect 13857 8132 13913 8188
rect 13913 8132 13917 8188
rect 13853 8128 13917 8132
rect 22054 8188 22118 8192
rect 22054 8132 22058 8188
rect 22058 8132 22114 8188
rect 22114 8132 22118 8188
rect 22054 8128 22118 8132
rect 22134 8188 22198 8192
rect 22134 8132 22138 8188
rect 22138 8132 22194 8188
rect 22194 8132 22198 8188
rect 22134 8128 22198 8132
rect 22214 8188 22278 8192
rect 22214 8132 22218 8188
rect 22218 8132 22274 8188
rect 22274 8132 22278 8188
rect 22214 8128 22278 8132
rect 22294 8188 22358 8192
rect 22294 8132 22298 8188
rect 22298 8132 22354 8188
rect 22354 8132 22358 8188
rect 22294 8128 22358 8132
rect 30495 8188 30559 8192
rect 30495 8132 30499 8188
rect 30499 8132 30555 8188
rect 30555 8132 30559 8188
rect 30495 8128 30559 8132
rect 30575 8188 30639 8192
rect 30575 8132 30579 8188
rect 30579 8132 30635 8188
rect 30635 8132 30639 8188
rect 30575 8128 30639 8132
rect 30655 8188 30719 8192
rect 30655 8132 30659 8188
rect 30659 8132 30715 8188
rect 30715 8132 30719 8188
rect 30655 8128 30719 8132
rect 30735 8188 30799 8192
rect 30735 8132 30739 8188
rect 30739 8132 30795 8188
rect 30795 8132 30799 8188
rect 30735 8128 30799 8132
rect 9392 7644 9456 7648
rect 9392 7588 9396 7644
rect 9396 7588 9452 7644
rect 9452 7588 9456 7644
rect 9392 7584 9456 7588
rect 9472 7644 9536 7648
rect 9472 7588 9476 7644
rect 9476 7588 9532 7644
rect 9532 7588 9536 7644
rect 9472 7584 9536 7588
rect 9552 7644 9616 7648
rect 9552 7588 9556 7644
rect 9556 7588 9612 7644
rect 9612 7588 9616 7644
rect 9552 7584 9616 7588
rect 9632 7644 9696 7648
rect 9632 7588 9636 7644
rect 9636 7588 9692 7644
rect 9692 7588 9696 7644
rect 9632 7584 9696 7588
rect 17833 7644 17897 7648
rect 17833 7588 17837 7644
rect 17837 7588 17893 7644
rect 17893 7588 17897 7644
rect 17833 7584 17897 7588
rect 17913 7644 17977 7648
rect 17913 7588 17917 7644
rect 17917 7588 17973 7644
rect 17973 7588 17977 7644
rect 17913 7584 17977 7588
rect 17993 7644 18057 7648
rect 17993 7588 17997 7644
rect 17997 7588 18053 7644
rect 18053 7588 18057 7644
rect 17993 7584 18057 7588
rect 18073 7644 18137 7648
rect 18073 7588 18077 7644
rect 18077 7588 18133 7644
rect 18133 7588 18137 7644
rect 18073 7584 18137 7588
rect 26274 7644 26338 7648
rect 26274 7588 26278 7644
rect 26278 7588 26334 7644
rect 26334 7588 26338 7644
rect 26274 7584 26338 7588
rect 26354 7644 26418 7648
rect 26354 7588 26358 7644
rect 26358 7588 26414 7644
rect 26414 7588 26418 7644
rect 26354 7584 26418 7588
rect 26434 7644 26498 7648
rect 26434 7588 26438 7644
rect 26438 7588 26494 7644
rect 26494 7588 26498 7644
rect 26434 7584 26498 7588
rect 26514 7644 26578 7648
rect 26514 7588 26518 7644
rect 26518 7588 26574 7644
rect 26574 7588 26578 7644
rect 26514 7584 26578 7588
rect 34715 7644 34779 7648
rect 34715 7588 34719 7644
rect 34719 7588 34775 7644
rect 34775 7588 34779 7644
rect 34715 7584 34779 7588
rect 34795 7644 34859 7648
rect 34795 7588 34799 7644
rect 34799 7588 34855 7644
rect 34855 7588 34859 7644
rect 34795 7584 34859 7588
rect 34875 7644 34939 7648
rect 34875 7588 34879 7644
rect 34879 7588 34935 7644
rect 34935 7588 34939 7644
rect 34875 7584 34939 7588
rect 34955 7644 35019 7648
rect 34955 7588 34959 7644
rect 34959 7588 35015 7644
rect 35015 7588 35019 7644
rect 34955 7584 35019 7588
rect 5172 7100 5236 7104
rect 5172 7044 5176 7100
rect 5176 7044 5232 7100
rect 5232 7044 5236 7100
rect 5172 7040 5236 7044
rect 5252 7100 5316 7104
rect 5252 7044 5256 7100
rect 5256 7044 5312 7100
rect 5312 7044 5316 7100
rect 5252 7040 5316 7044
rect 5332 7100 5396 7104
rect 5332 7044 5336 7100
rect 5336 7044 5392 7100
rect 5392 7044 5396 7100
rect 5332 7040 5396 7044
rect 5412 7100 5476 7104
rect 5412 7044 5416 7100
rect 5416 7044 5472 7100
rect 5472 7044 5476 7100
rect 5412 7040 5476 7044
rect 13613 7100 13677 7104
rect 13613 7044 13617 7100
rect 13617 7044 13673 7100
rect 13673 7044 13677 7100
rect 13613 7040 13677 7044
rect 13693 7100 13757 7104
rect 13693 7044 13697 7100
rect 13697 7044 13753 7100
rect 13753 7044 13757 7100
rect 13693 7040 13757 7044
rect 13773 7100 13837 7104
rect 13773 7044 13777 7100
rect 13777 7044 13833 7100
rect 13833 7044 13837 7100
rect 13773 7040 13837 7044
rect 13853 7100 13917 7104
rect 13853 7044 13857 7100
rect 13857 7044 13913 7100
rect 13913 7044 13917 7100
rect 13853 7040 13917 7044
rect 22054 7100 22118 7104
rect 22054 7044 22058 7100
rect 22058 7044 22114 7100
rect 22114 7044 22118 7100
rect 22054 7040 22118 7044
rect 22134 7100 22198 7104
rect 22134 7044 22138 7100
rect 22138 7044 22194 7100
rect 22194 7044 22198 7100
rect 22134 7040 22198 7044
rect 22214 7100 22278 7104
rect 22214 7044 22218 7100
rect 22218 7044 22274 7100
rect 22274 7044 22278 7100
rect 22214 7040 22278 7044
rect 22294 7100 22358 7104
rect 22294 7044 22298 7100
rect 22298 7044 22354 7100
rect 22354 7044 22358 7100
rect 22294 7040 22358 7044
rect 30495 7100 30559 7104
rect 30495 7044 30499 7100
rect 30499 7044 30555 7100
rect 30555 7044 30559 7100
rect 30495 7040 30559 7044
rect 30575 7100 30639 7104
rect 30575 7044 30579 7100
rect 30579 7044 30635 7100
rect 30635 7044 30639 7100
rect 30575 7040 30639 7044
rect 30655 7100 30719 7104
rect 30655 7044 30659 7100
rect 30659 7044 30715 7100
rect 30715 7044 30719 7100
rect 30655 7040 30719 7044
rect 30735 7100 30799 7104
rect 30735 7044 30739 7100
rect 30739 7044 30795 7100
rect 30795 7044 30799 7100
rect 30735 7040 30799 7044
rect 9392 6556 9456 6560
rect 9392 6500 9396 6556
rect 9396 6500 9452 6556
rect 9452 6500 9456 6556
rect 9392 6496 9456 6500
rect 9472 6556 9536 6560
rect 9472 6500 9476 6556
rect 9476 6500 9532 6556
rect 9532 6500 9536 6556
rect 9472 6496 9536 6500
rect 9552 6556 9616 6560
rect 9552 6500 9556 6556
rect 9556 6500 9612 6556
rect 9612 6500 9616 6556
rect 9552 6496 9616 6500
rect 9632 6556 9696 6560
rect 9632 6500 9636 6556
rect 9636 6500 9692 6556
rect 9692 6500 9696 6556
rect 9632 6496 9696 6500
rect 17833 6556 17897 6560
rect 17833 6500 17837 6556
rect 17837 6500 17893 6556
rect 17893 6500 17897 6556
rect 17833 6496 17897 6500
rect 17913 6556 17977 6560
rect 17913 6500 17917 6556
rect 17917 6500 17973 6556
rect 17973 6500 17977 6556
rect 17913 6496 17977 6500
rect 17993 6556 18057 6560
rect 17993 6500 17997 6556
rect 17997 6500 18053 6556
rect 18053 6500 18057 6556
rect 17993 6496 18057 6500
rect 18073 6556 18137 6560
rect 18073 6500 18077 6556
rect 18077 6500 18133 6556
rect 18133 6500 18137 6556
rect 18073 6496 18137 6500
rect 26274 6556 26338 6560
rect 26274 6500 26278 6556
rect 26278 6500 26334 6556
rect 26334 6500 26338 6556
rect 26274 6496 26338 6500
rect 26354 6556 26418 6560
rect 26354 6500 26358 6556
rect 26358 6500 26414 6556
rect 26414 6500 26418 6556
rect 26354 6496 26418 6500
rect 26434 6556 26498 6560
rect 26434 6500 26438 6556
rect 26438 6500 26494 6556
rect 26494 6500 26498 6556
rect 26434 6496 26498 6500
rect 26514 6556 26578 6560
rect 26514 6500 26518 6556
rect 26518 6500 26574 6556
rect 26574 6500 26578 6556
rect 26514 6496 26578 6500
rect 34715 6556 34779 6560
rect 34715 6500 34719 6556
rect 34719 6500 34775 6556
rect 34775 6500 34779 6556
rect 34715 6496 34779 6500
rect 34795 6556 34859 6560
rect 34795 6500 34799 6556
rect 34799 6500 34855 6556
rect 34855 6500 34859 6556
rect 34795 6496 34859 6500
rect 34875 6556 34939 6560
rect 34875 6500 34879 6556
rect 34879 6500 34935 6556
rect 34935 6500 34939 6556
rect 34875 6496 34939 6500
rect 34955 6556 35019 6560
rect 34955 6500 34959 6556
rect 34959 6500 35015 6556
rect 35015 6500 35019 6556
rect 34955 6496 35019 6500
rect 5172 6012 5236 6016
rect 5172 5956 5176 6012
rect 5176 5956 5232 6012
rect 5232 5956 5236 6012
rect 5172 5952 5236 5956
rect 5252 6012 5316 6016
rect 5252 5956 5256 6012
rect 5256 5956 5312 6012
rect 5312 5956 5316 6012
rect 5252 5952 5316 5956
rect 5332 6012 5396 6016
rect 5332 5956 5336 6012
rect 5336 5956 5392 6012
rect 5392 5956 5396 6012
rect 5332 5952 5396 5956
rect 5412 6012 5476 6016
rect 5412 5956 5416 6012
rect 5416 5956 5472 6012
rect 5472 5956 5476 6012
rect 5412 5952 5476 5956
rect 13613 6012 13677 6016
rect 13613 5956 13617 6012
rect 13617 5956 13673 6012
rect 13673 5956 13677 6012
rect 13613 5952 13677 5956
rect 13693 6012 13757 6016
rect 13693 5956 13697 6012
rect 13697 5956 13753 6012
rect 13753 5956 13757 6012
rect 13693 5952 13757 5956
rect 13773 6012 13837 6016
rect 13773 5956 13777 6012
rect 13777 5956 13833 6012
rect 13833 5956 13837 6012
rect 13773 5952 13837 5956
rect 13853 6012 13917 6016
rect 13853 5956 13857 6012
rect 13857 5956 13913 6012
rect 13913 5956 13917 6012
rect 13853 5952 13917 5956
rect 22054 6012 22118 6016
rect 22054 5956 22058 6012
rect 22058 5956 22114 6012
rect 22114 5956 22118 6012
rect 22054 5952 22118 5956
rect 22134 6012 22198 6016
rect 22134 5956 22138 6012
rect 22138 5956 22194 6012
rect 22194 5956 22198 6012
rect 22134 5952 22198 5956
rect 22214 6012 22278 6016
rect 22214 5956 22218 6012
rect 22218 5956 22274 6012
rect 22274 5956 22278 6012
rect 22214 5952 22278 5956
rect 22294 6012 22358 6016
rect 22294 5956 22298 6012
rect 22298 5956 22354 6012
rect 22354 5956 22358 6012
rect 22294 5952 22358 5956
rect 30495 6012 30559 6016
rect 30495 5956 30499 6012
rect 30499 5956 30555 6012
rect 30555 5956 30559 6012
rect 30495 5952 30559 5956
rect 30575 6012 30639 6016
rect 30575 5956 30579 6012
rect 30579 5956 30635 6012
rect 30635 5956 30639 6012
rect 30575 5952 30639 5956
rect 30655 6012 30719 6016
rect 30655 5956 30659 6012
rect 30659 5956 30715 6012
rect 30715 5956 30719 6012
rect 30655 5952 30719 5956
rect 30735 6012 30799 6016
rect 30735 5956 30739 6012
rect 30739 5956 30795 6012
rect 30795 5956 30799 6012
rect 30735 5952 30799 5956
rect 9392 5468 9456 5472
rect 9392 5412 9396 5468
rect 9396 5412 9452 5468
rect 9452 5412 9456 5468
rect 9392 5408 9456 5412
rect 9472 5468 9536 5472
rect 9472 5412 9476 5468
rect 9476 5412 9532 5468
rect 9532 5412 9536 5468
rect 9472 5408 9536 5412
rect 9552 5468 9616 5472
rect 9552 5412 9556 5468
rect 9556 5412 9612 5468
rect 9612 5412 9616 5468
rect 9552 5408 9616 5412
rect 9632 5468 9696 5472
rect 9632 5412 9636 5468
rect 9636 5412 9692 5468
rect 9692 5412 9696 5468
rect 9632 5408 9696 5412
rect 17833 5468 17897 5472
rect 17833 5412 17837 5468
rect 17837 5412 17893 5468
rect 17893 5412 17897 5468
rect 17833 5408 17897 5412
rect 17913 5468 17977 5472
rect 17913 5412 17917 5468
rect 17917 5412 17973 5468
rect 17973 5412 17977 5468
rect 17913 5408 17977 5412
rect 17993 5468 18057 5472
rect 17993 5412 17997 5468
rect 17997 5412 18053 5468
rect 18053 5412 18057 5468
rect 17993 5408 18057 5412
rect 18073 5468 18137 5472
rect 18073 5412 18077 5468
rect 18077 5412 18133 5468
rect 18133 5412 18137 5468
rect 18073 5408 18137 5412
rect 26274 5468 26338 5472
rect 26274 5412 26278 5468
rect 26278 5412 26334 5468
rect 26334 5412 26338 5468
rect 26274 5408 26338 5412
rect 26354 5468 26418 5472
rect 26354 5412 26358 5468
rect 26358 5412 26414 5468
rect 26414 5412 26418 5468
rect 26354 5408 26418 5412
rect 26434 5468 26498 5472
rect 26434 5412 26438 5468
rect 26438 5412 26494 5468
rect 26494 5412 26498 5468
rect 26434 5408 26498 5412
rect 26514 5468 26578 5472
rect 26514 5412 26518 5468
rect 26518 5412 26574 5468
rect 26574 5412 26578 5468
rect 26514 5408 26578 5412
rect 34715 5468 34779 5472
rect 34715 5412 34719 5468
rect 34719 5412 34775 5468
rect 34775 5412 34779 5468
rect 34715 5408 34779 5412
rect 34795 5468 34859 5472
rect 34795 5412 34799 5468
rect 34799 5412 34855 5468
rect 34855 5412 34859 5468
rect 34795 5408 34859 5412
rect 34875 5468 34939 5472
rect 34875 5412 34879 5468
rect 34879 5412 34935 5468
rect 34935 5412 34939 5468
rect 34875 5408 34939 5412
rect 34955 5468 35019 5472
rect 34955 5412 34959 5468
rect 34959 5412 35015 5468
rect 35015 5412 35019 5468
rect 34955 5408 35019 5412
rect 5172 4924 5236 4928
rect 5172 4868 5176 4924
rect 5176 4868 5232 4924
rect 5232 4868 5236 4924
rect 5172 4864 5236 4868
rect 5252 4924 5316 4928
rect 5252 4868 5256 4924
rect 5256 4868 5312 4924
rect 5312 4868 5316 4924
rect 5252 4864 5316 4868
rect 5332 4924 5396 4928
rect 5332 4868 5336 4924
rect 5336 4868 5392 4924
rect 5392 4868 5396 4924
rect 5332 4864 5396 4868
rect 5412 4924 5476 4928
rect 5412 4868 5416 4924
rect 5416 4868 5472 4924
rect 5472 4868 5476 4924
rect 5412 4864 5476 4868
rect 13613 4924 13677 4928
rect 13613 4868 13617 4924
rect 13617 4868 13673 4924
rect 13673 4868 13677 4924
rect 13613 4864 13677 4868
rect 13693 4924 13757 4928
rect 13693 4868 13697 4924
rect 13697 4868 13753 4924
rect 13753 4868 13757 4924
rect 13693 4864 13757 4868
rect 13773 4924 13837 4928
rect 13773 4868 13777 4924
rect 13777 4868 13833 4924
rect 13833 4868 13837 4924
rect 13773 4864 13837 4868
rect 13853 4924 13917 4928
rect 13853 4868 13857 4924
rect 13857 4868 13913 4924
rect 13913 4868 13917 4924
rect 13853 4864 13917 4868
rect 22054 4924 22118 4928
rect 22054 4868 22058 4924
rect 22058 4868 22114 4924
rect 22114 4868 22118 4924
rect 22054 4864 22118 4868
rect 22134 4924 22198 4928
rect 22134 4868 22138 4924
rect 22138 4868 22194 4924
rect 22194 4868 22198 4924
rect 22134 4864 22198 4868
rect 22214 4924 22278 4928
rect 22214 4868 22218 4924
rect 22218 4868 22274 4924
rect 22274 4868 22278 4924
rect 22214 4864 22278 4868
rect 22294 4924 22358 4928
rect 22294 4868 22298 4924
rect 22298 4868 22354 4924
rect 22354 4868 22358 4924
rect 22294 4864 22358 4868
rect 30495 4924 30559 4928
rect 30495 4868 30499 4924
rect 30499 4868 30555 4924
rect 30555 4868 30559 4924
rect 30495 4864 30559 4868
rect 30575 4924 30639 4928
rect 30575 4868 30579 4924
rect 30579 4868 30635 4924
rect 30635 4868 30639 4924
rect 30575 4864 30639 4868
rect 30655 4924 30719 4928
rect 30655 4868 30659 4924
rect 30659 4868 30715 4924
rect 30715 4868 30719 4924
rect 30655 4864 30719 4868
rect 30735 4924 30799 4928
rect 30735 4868 30739 4924
rect 30739 4868 30795 4924
rect 30795 4868 30799 4924
rect 30735 4864 30799 4868
rect 9392 4380 9456 4384
rect 9392 4324 9396 4380
rect 9396 4324 9452 4380
rect 9452 4324 9456 4380
rect 9392 4320 9456 4324
rect 9472 4380 9536 4384
rect 9472 4324 9476 4380
rect 9476 4324 9532 4380
rect 9532 4324 9536 4380
rect 9472 4320 9536 4324
rect 9552 4380 9616 4384
rect 9552 4324 9556 4380
rect 9556 4324 9612 4380
rect 9612 4324 9616 4380
rect 9552 4320 9616 4324
rect 9632 4380 9696 4384
rect 9632 4324 9636 4380
rect 9636 4324 9692 4380
rect 9692 4324 9696 4380
rect 9632 4320 9696 4324
rect 17833 4380 17897 4384
rect 17833 4324 17837 4380
rect 17837 4324 17893 4380
rect 17893 4324 17897 4380
rect 17833 4320 17897 4324
rect 17913 4380 17977 4384
rect 17913 4324 17917 4380
rect 17917 4324 17973 4380
rect 17973 4324 17977 4380
rect 17913 4320 17977 4324
rect 17993 4380 18057 4384
rect 17993 4324 17997 4380
rect 17997 4324 18053 4380
rect 18053 4324 18057 4380
rect 17993 4320 18057 4324
rect 18073 4380 18137 4384
rect 18073 4324 18077 4380
rect 18077 4324 18133 4380
rect 18133 4324 18137 4380
rect 18073 4320 18137 4324
rect 26274 4380 26338 4384
rect 26274 4324 26278 4380
rect 26278 4324 26334 4380
rect 26334 4324 26338 4380
rect 26274 4320 26338 4324
rect 26354 4380 26418 4384
rect 26354 4324 26358 4380
rect 26358 4324 26414 4380
rect 26414 4324 26418 4380
rect 26354 4320 26418 4324
rect 26434 4380 26498 4384
rect 26434 4324 26438 4380
rect 26438 4324 26494 4380
rect 26494 4324 26498 4380
rect 26434 4320 26498 4324
rect 26514 4380 26578 4384
rect 26514 4324 26518 4380
rect 26518 4324 26574 4380
rect 26574 4324 26578 4380
rect 26514 4320 26578 4324
rect 34715 4380 34779 4384
rect 34715 4324 34719 4380
rect 34719 4324 34775 4380
rect 34775 4324 34779 4380
rect 34715 4320 34779 4324
rect 34795 4380 34859 4384
rect 34795 4324 34799 4380
rect 34799 4324 34855 4380
rect 34855 4324 34859 4380
rect 34795 4320 34859 4324
rect 34875 4380 34939 4384
rect 34875 4324 34879 4380
rect 34879 4324 34935 4380
rect 34935 4324 34939 4380
rect 34875 4320 34939 4324
rect 34955 4380 35019 4384
rect 34955 4324 34959 4380
rect 34959 4324 35015 4380
rect 35015 4324 35019 4380
rect 34955 4320 35019 4324
rect 5172 3836 5236 3840
rect 5172 3780 5176 3836
rect 5176 3780 5232 3836
rect 5232 3780 5236 3836
rect 5172 3776 5236 3780
rect 5252 3836 5316 3840
rect 5252 3780 5256 3836
rect 5256 3780 5312 3836
rect 5312 3780 5316 3836
rect 5252 3776 5316 3780
rect 5332 3836 5396 3840
rect 5332 3780 5336 3836
rect 5336 3780 5392 3836
rect 5392 3780 5396 3836
rect 5332 3776 5396 3780
rect 5412 3836 5476 3840
rect 5412 3780 5416 3836
rect 5416 3780 5472 3836
rect 5472 3780 5476 3836
rect 5412 3776 5476 3780
rect 13613 3836 13677 3840
rect 13613 3780 13617 3836
rect 13617 3780 13673 3836
rect 13673 3780 13677 3836
rect 13613 3776 13677 3780
rect 13693 3836 13757 3840
rect 13693 3780 13697 3836
rect 13697 3780 13753 3836
rect 13753 3780 13757 3836
rect 13693 3776 13757 3780
rect 13773 3836 13837 3840
rect 13773 3780 13777 3836
rect 13777 3780 13833 3836
rect 13833 3780 13837 3836
rect 13773 3776 13837 3780
rect 13853 3836 13917 3840
rect 13853 3780 13857 3836
rect 13857 3780 13913 3836
rect 13913 3780 13917 3836
rect 13853 3776 13917 3780
rect 22054 3836 22118 3840
rect 22054 3780 22058 3836
rect 22058 3780 22114 3836
rect 22114 3780 22118 3836
rect 22054 3776 22118 3780
rect 22134 3836 22198 3840
rect 22134 3780 22138 3836
rect 22138 3780 22194 3836
rect 22194 3780 22198 3836
rect 22134 3776 22198 3780
rect 22214 3836 22278 3840
rect 22214 3780 22218 3836
rect 22218 3780 22274 3836
rect 22274 3780 22278 3836
rect 22214 3776 22278 3780
rect 22294 3836 22358 3840
rect 22294 3780 22298 3836
rect 22298 3780 22354 3836
rect 22354 3780 22358 3836
rect 22294 3776 22358 3780
rect 30495 3836 30559 3840
rect 30495 3780 30499 3836
rect 30499 3780 30555 3836
rect 30555 3780 30559 3836
rect 30495 3776 30559 3780
rect 30575 3836 30639 3840
rect 30575 3780 30579 3836
rect 30579 3780 30635 3836
rect 30635 3780 30639 3836
rect 30575 3776 30639 3780
rect 30655 3836 30719 3840
rect 30655 3780 30659 3836
rect 30659 3780 30715 3836
rect 30715 3780 30719 3836
rect 30655 3776 30719 3780
rect 30735 3836 30799 3840
rect 30735 3780 30739 3836
rect 30739 3780 30795 3836
rect 30795 3780 30799 3836
rect 30735 3776 30799 3780
rect 9392 3292 9456 3296
rect 9392 3236 9396 3292
rect 9396 3236 9452 3292
rect 9452 3236 9456 3292
rect 9392 3232 9456 3236
rect 9472 3292 9536 3296
rect 9472 3236 9476 3292
rect 9476 3236 9532 3292
rect 9532 3236 9536 3292
rect 9472 3232 9536 3236
rect 9552 3292 9616 3296
rect 9552 3236 9556 3292
rect 9556 3236 9612 3292
rect 9612 3236 9616 3292
rect 9552 3232 9616 3236
rect 9632 3292 9696 3296
rect 9632 3236 9636 3292
rect 9636 3236 9692 3292
rect 9692 3236 9696 3292
rect 9632 3232 9696 3236
rect 17833 3292 17897 3296
rect 17833 3236 17837 3292
rect 17837 3236 17893 3292
rect 17893 3236 17897 3292
rect 17833 3232 17897 3236
rect 17913 3292 17977 3296
rect 17913 3236 17917 3292
rect 17917 3236 17973 3292
rect 17973 3236 17977 3292
rect 17913 3232 17977 3236
rect 17993 3292 18057 3296
rect 17993 3236 17997 3292
rect 17997 3236 18053 3292
rect 18053 3236 18057 3292
rect 17993 3232 18057 3236
rect 18073 3292 18137 3296
rect 18073 3236 18077 3292
rect 18077 3236 18133 3292
rect 18133 3236 18137 3292
rect 18073 3232 18137 3236
rect 26274 3292 26338 3296
rect 26274 3236 26278 3292
rect 26278 3236 26334 3292
rect 26334 3236 26338 3292
rect 26274 3232 26338 3236
rect 26354 3292 26418 3296
rect 26354 3236 26358 3292
rect 26358 3236 26414 3292
rect 26414 3236 26418 3292
rect 26354 3232 26418 3236
rect 26434 3292 26498 3296
rect 26434 3236 26438 3292
rect 26438 3236 26494 3292
rect 26494 3236 26498 3292
rect 26434 3232 26498 3236
rect 26514 3292 26578 3296
rect 26514 3236 26518 3292
rect 26518 3236 26574 3292
rect 26574 3236 26578 3292
rect 26514 3232 26578 3236
rect 34715 3292 34779 3296
rect 34715 3236 34719 3292
rect 34719 3236 34775 3292
rect 34775 3236 34779 3292
rect 34715 3232 34779 3236
rect 34795 3292 34859 3296
rect 34795 3236 34799 3292
rect 34799 3236 34855 3292
rect 34855 3236 34859 3292
rect 34795 3232 34859 3236
rect 34875 3292 34939 3296
rect 34875 3236 34879 3292
rect 34879 3236 34935 3292
rect 34935 3236 34939 3292
rect 34875 3232 34939 3236
rect 34955 3292 35019 3296
rect 34955 3236 34959 3292
rect 34959 3236 35015 3292
rect 35015 3236 35019 3292
rect 34955 3232 35019 3236
rect 5172 2748 5236 2752
rect 5172 2692 5176 2748
rect 5176 2692 5232 2748
rect 5232 2692 5236 2748
rect 5172 2688 5236 2692
rect 5252 2748 5316 2752
rect 5252 2692 5256 2748
rect 5256 2692 5312 2748
rect 5312 2692 5316 2748
rect 5252 2688 5316 2692
rect 5332 2748 5396 2752
rect 5332 2692 5336 2748
rect 5336 2692 5392 2748
rect 5392 2692 5396 2748
rect 5332 2688 5396 2692
rect 5412 2748 5476 2752
rect 5412 2692 5416 2748
rect 5416 2692 5472 2748
rect 5472 2692 5476 2748
rect 5412 2688 5476 2692
rect 13613 2748 13677 2752
rect 13613 2692 13617 2748
rect 13617 2692 13673 2748
rect 13673 2692 13677 2748
rect 13613 2688 13677 2692
rect 13693 2748 13757 2752
rect 13693 2692 13697 2748
rect 13697 2692 13753 2748
rect 13753 2692 13757 2748
rect 13693 2688 13757 2692
rect 13773 2748 13837 2752
rect 13773 2692 13777 2748
rect 13777 2692 13833 2748
rect 13833 2692 13837 2748
rect 13773 2688 13837 2692
rect 13853 2748 13917 2752
rect 13853 2692 13857 2748
rect 13857 2692 13913 2748
rect 13913 2692 13917 2748
rect 13853 2688 13917 2692
rect 22054 2748 22118 2752
rect 22054 2692 22058 2748
rect 22058 2692 22114 2748
rect 22114 2692 22118 2748
rect 22054 2688 22118 2692
rect 22134 2748 22198 2752
rect 22134 2692 22138 2748
rect 22138 2692 22194 2748
rect 22194 2692 22198 2748
rect 22134 2688 22198 2692
rect 22214 2748 22278 2752
rect 22214 2692 22218 2748
rect 22218 2692 22274 2748
rect 22274 2692 22278 2748
rect 22214 2688 22278 2692
rect 22294 2748 22358 2752
rect 22294 2692 22298 2748
rect 22298 2692 22354 2748
rect 22354 2692 22358 2748
rect 22294 2688 22358 2692
rect 30495 2748 30559 2752
rect 30495 2692 30499 2748
rect 30499 2692 30555 2748
rect 30555 2692 30559 2748
rect 30495 2688 30559 2692
rect 30575 2748 30639 2752
rect 30575 2692 30579 2748
rect 30579 2692 30635 2748
rect 30635 2692 30639 2748
rect 30575 2688 30639 2692
rect 30655 2748 30719 2752
rect 30655 2692 30659 2748
rect 30659 2692 30715 2748
rect 30715 2692 30719 2748
rect 30655 2688 30719 2692
rect 30735 2748 30799 2752
rect 30735 2692 30739 2748
rect 30739 2692 30795 2748
rect 30795 2692 30799 2748
rect 30735 2688 30799 2692
rect 9392 2204 9456 2208
rect 9392 2148 9396 2204
rect 9396 2148 9452 2204
rect 9452 2148 9456 2204
rect 9392 2144 9456 2148
rect 9472 2204 9536 2208
rect 9472 2148 9476 2204
rect 9476 2148 9532 2204
rect 9532 2148 9536 2204
rect 9472 2144 9536 2148
rect 9552 2204 9616 2208
rect 9552 2148 9556 2204
rect 9556 2148 9612 2204
rect 9612 2148 9616 2204
rect 9552 2144 9616 2148
rect 9632 2204 9696 2208
rect 9632 2148 9636 2204
rect 9636 2148 9692 2204
rect 9692 2148 9696 2204
rect 9632 2144 9696 2148
rect 17833 2204 17897 2208
rect 17833 2148 17837 2204
rect 17837 2148 17893 2204
rect 17893 2148 17897 2204
rect 17833 2144 17897 2148
rect 17913 2204 17977 2208
rect 17913 2148 17917 2204
rect 17917 2148 17973 2204
rect 17973 2148 17977 2204
rect 17913 2144 17977 2148
rect 17993 2204 18057 2208
rect 17993 2148 17997 2204
rect 17997 2148 18053 2204
rect 18053 2148 18057 2204
rect 17993 2144 18057 2148
rect 18073 2204 18137 2208
rect 18073 2148 18077 2204
rect 18077 2148 18133 2204
rect 18133 2148 18137 2204
rect 18073 2144 18137 2148
rect 26274 2204 26338 2208
rect 26274 2148 26278 2204
rect 26278 2148 26334 2204
rect 26334 2148 26338 2204
rect 26274 2144 26338 2148
rect 26354 2204 26418 2208
rect 26354 2148 26358 2204
rect 26358 2148 26414 2204
rect 26414 2148 26418 2204
rect 26354 2144 26418 2148
rect 26434 2204 26498 2208
rect 26434 2148 26438 2204
rect 26438 2148 26494 2204
rect 26494 2148 26498 2204
rect 26434 2144 26498 2148
rect 26514 2204 26578 2208
rect 26514 2148 26518 2204
rect 26518 2148 26574 2204
rect 26574 2148 26578 2204
rect 26514 2144 26578 2148
rect 34715 2204 34779 2208
rect 34715 2148 34719 2204
rect 34719 2148 34775 2204
rect 34775 2148 34779 2204
rect 34715 2144 34779 2148
rect 34795 2204 34859 2208
rect 34795 2148 34799 2204
rect 34799 2148 34855 2204
rect 34855 2148 34859 2204
rect 34795 2144 34859 2148
rect 34875 2204 34939 2208
rect 34875 2148 34879 2204
rect 34879 2148 34935 2204
rect 34935 2148 34939 2204
rect 34875 2144 34939 2148
rect 34955 2204 35019 2208
rect 34955 2148 34959 2204
rect 34959 2148 35015 2204
rect 35015 2148 35019 2204
rect 34955 2144 35019 2148
<< metal4 >>
rect 5164 39744 5484 39760
rect 5164 39680 5172 39744
rect 5236 39680 5252 39744
rect 5316 39680 5332 39744
rect 5396 39680 5412 39744
rect 5476 39680 5484 39744
rect 5164 38656 5484 39680
rect 5164 38592 5172 38656
rect 5236 38592 5252 38656
rect 5316 38592 5332 38656
rect 5396 38592 5412 38656
rect 5476 38592 5484 38656
rect 5164 37568 5484 38592
rect 5164 37504 5172 37568
rect 5236 37504 5252 37568
rect 5316 37504 5332 37568
rect 5396 37504 5412 37568
rect 5476 37504 5484 37568
rect 5164 36480 5484 37504
rect 5164 36416 5172 36480
rect 5236 36416 5252 36480
rect 5316 36416 5332 36480
rect 5396 36416 5412 36480
rect 5476 36416 5484 36480
rect 5164 35392 5484 36416
rect 5164 35328 5172 35392
rect 5236 35328 5252 35392
rect 5316 35328 5332 35392
rect 5396 35328 5412 35392
rect 5476 35328 5484 35392
rect 5164 34304 5484 35328
rect 5164 34240 5172 34304
rect 5236 34240 5252 34304
rect 5316 34240 5332 34304
rect 5396 34240 5412 34304
rect 5476 34240 5484 34304
rect 5164 33216 5484 34240
rect 5164 33152 5172 33216
rect 5236 33152 5252 33216
rect 5316 33152 5332 33216
rect 5396 33152 5412 33216
rect 5476 33152 5484 33216
rect 5164 32128 5484 33152
rect 5164 32064 5172 32128
rect 5236 32064 5252 32128
rect 5316 32064 5332 32128
rect 5396 32064 5412 32128
rect 5476 32064 5484 32128
rect 5164 31040 5484 32064
rect 5164 30976 5172 31040
rect 5236 30976 5252 31040
rect 5316 30976 5332 31040
rect 5396 30976 5412 31040
rect 5476 30976 5484 31040
rect 5164 29952 5484 30976
rect 5164 29888 5172 29952
rect 5236 29888 5252 29952
rect 5316 29888 5332 29952
rect 5396 29888 5412 29952
rect 5476 29888 5484 29952
rect 5164 28864 5484 29888
rect 5164 28800 5172 28864
rect 5236 28800 5252 28864
rect 5316 28800 5332 28864
rect 5396 28800 5412 28864
rect 5476 28800 5484 28864
rect 5164 27776 5484 28800
rect 5164 27712 5172 27776
rect 5236 27712 5252 27776
rect 5316 27712 5332 27776
rect 5396 27712 5412 27776
rect 5476 27712 5484 27776
rect 5164 26688 5484 27712
rect 5164 26624 5172 26688
rect 5236 26624 5252 26688
rect 5316 26624 5332 26688
rect 5396 26624 5412 26688
rect 5476 26624 5484 26688
rect 5164 25600 5484 26624
rect 5164 25536 5172 25600
rect 5236 25536 5252 25600
rect 5316 25536 5332 25600
rect 5396 25536 5412 25600
rect 5476 25536 5484 25600
rect 5164 24512 5484 25536
rect 5164 24448 5172 24512
rect 5236 24448 5252 24512
rect 5316 24448 5332 24512
rect 5396 24448 5412 24512
rect 5476 24448 5484 24512
rect 5164 23424 5484 24448
rect 5164 23360 5172 23424
rect 5236 23360 5252 23424
rect 5316 23360 5332 23424
rect 5396 23360 5412 23424
rect 5476 23360 5484 23424
rect 5164 22336 5484 23360
rect 5164 22272 5172 22336
rect 5236 22272 5252 22336
rect 5316 22272 5332 22336
rect 5396 22272 5412 22336
rect 5476 22272 5484 22336
rect 5164 21248 5484 22272
rect 5164 21184 5172 21248
rect 5236 21184 5252 21248
rect 5316 21184 5332 21248
rect 5396 21184 5412 21248
rect 5476 21184 5484 21248
rect 5164 20160 5484 21184
rect 5164 20096 5172 20160
rect 5236 20096 5252 20160
rect 5316 20096 5332 20160
rect 5396 20096 5412 20160
rect 5476 20096 5484 20160
rect 5164 19072 5484 20096
rect 5164 19008 5172 19072
rect 5236 19008 5252 19072
rect 5316 19008 5332 19072
rect 5396 19008 5412 19072
rect 5476 19008 5484 19072
rect 5164 17984 5484 19008
rect 5164 17920 5172 17984
rect 5236 17920 5252 17984
rect 5316 17920 5332 17984
rect 5396 17920 5412 17984
rect 5476 17920 5484 17984
rect 5164 16896 5484 17920
rect 5164 16832 5172 16896
rect 5236 16832 5252 16896
rect 5316 16832 5332 16896
rect 5396 16832 5412 16896
rect 5476 16832 5484 16896
rect 5164 15808 5484 16832
rect 5164 15744 5172 15808
rect 5236 15744 5252 15808
rect 5316 15744 5332 15808
rect 5396 15744 5412 15808
rect 5476 15744 5484 15808
rect 5164 14720 5484 15744
rect 5164 14656 5172 14720
rect 5236 14656 5252 14720
rect 5316 14656 5332 14720
rect 5396 14656 5412 14720
rect 5476 14656 5484 14720
rect 5164 13632 5484 14656
rect 5164 13568 5172 13632
rect 5236 13568 5252 13632
rect 5316 13568 5332 13632
rect 5396 13568 5412 13632
rect 5476 13568 5484 13632
rect 5164 12544 5484 13568
rect 5164 12480 5172 12544
rect 5236 12480 5252 12544
rect 5316 12480 5332 12544
rect 5396 12480 5412 12544
rect 5476 12480 5484 12544
rect 5164 11456 5484 12480
rect 5164 11392 5172 11456
rect 5236 11392 5252 11456
rect 5316 11392 5332 11456
rect 5396 11392 5412 11456
rect 5476 11392 5484 11456
rect 5164 10368 5484 11392
rect 5164 10304 5172 10368
rect 5236 10304 5252 10368
rect 5316 10304 5332 10368
rect 5396 10304 5412 10368
rect 5476 10304 5484 10368
rect 5164 9280 5484 10304
rect 5164 9216 5172 9280
rect 5236 9216 5252 9280
rect 5316 9216 5332 9280
rect 5396 9216 5412 9280
rect 5476 9216 5484 9280
rect 5164 8192 5484 9216
rect 5164 8128 5172 8192
rect 5236 8128 5252 8192
rect 5316 8128 5332 8192
rect 5396 8128 5412 8192
rect 5476 8128 5484 8192
rect 5164 7104 5484 8128
rect 5164 7040 5172 7104
rect 5236 7040 5252 7104
rect 5316 7040 5332 7104
rect 5396 7040 5412 7104
rect 5476 7040 5484 7104
rect 5164 6016 5484 7040
rect 5164 5952 5172 6016
rect 5236 5952 5252 6016
rect 5316 5952 5332 6016
rect 5396 5952 5412 6016
rect 5476 5952 5484 6016
rect 5164 4928 5484 5952
rect 5164 4864 5172 4928
rect 5236 4864 5252 4928
rect 5316 4864 5332 4928
rect 5396 4864 5412 4928
rect 5476 4864 5484 4928
rect 5164 3840 5484 4864
rect 5164 3776 5172 3840
rect 5236 3776 5252 3840
rect 5316 3776 5332 3840
rect 5396 3776 5412 3840
rect 5476 3776 5484 3840
rect 5164 2752 5484 3776
rect 5164 2688 5172 2752
rect 5236 2688 5252 2752
rect 5316 2688 5332 2752
rect 5396 2688 5412 2752
rect 5476 2688 5484 2752
rect 5164 2128 5484 2688
rect 9384 39200 9704 39760
rect 9384 39136 9392 39200
rect 9456 39136 9472 39200
rect 9536 39136 9552 39200
rect 9616 39136 9632 39200
rect 9696 39136 9704 39200
rect 9384 38112 9704 39136
rect 9384 38048 9392 38112
rect 9456 38048 9472 38112
rect 9536 38048 9552 38112
rect 9616 38048 9632 38112
rect 9696 38048 9704 38112
rect 9384 37024 9704 38048
rect 9384 36960 9392 37024
rect 9456 36960 9472 37024
rect 9536 36960 9552 37024
rect 9616 36960 9632 37024
rect 9696 36960 9704 37024
rect 9384 35936 9704 36960
rect 9384 35872 9392 35936
rect 9456 35872 9472 35936
rect 9536 35872 9552 35936
rect 9616 35872 9632 35936
rect 9696 35872 9704 35936
rect 9384 34848 9704 35872
rect 9384 34784 9392 34848
rect 9456 34784 9472 34848
rect 9536 34784 9552 34848
rect 9616 34784 9632 34848
rect 9696 34784 9704 34848
rect 9384 33760 9704 34784
rect 9384 33696 9392 33760
rect 9456 33696 9472 33760
rect 9536 33696 9552 33760
rect 9616 33696 9632 33760
rect 9696 33696 9704 33760
rect 9384 32672 9704 33696
rect 9384 32608 9392 32672
rect 9456 32608 9472 32672
rect 9536 32608 9552 32672
rect 9616 32608 9632 32672
rect 9696 32608 9704 32672
rect 9384 31584 9704 32608
rect 9384 31520 9392 31584
rect 9456 31520 9472 31584
rect 9536 31520 9552 31584
rect 9616 31520 9632 31584
rect 9696 31520 9704 31584
rect 9384 30496 9704 31520
rect 9384 30432 9392 30496
rect 9456 30432 9472 30496
rect 9536 30432 9552 30496
rect 9616 30432 9632 30496
rect 9696 30432 9704 30496
rect 9384 29408 9704 30432
rect 9384 29344 9392 29408
rect 9456 29344 9472 29408
rect 9536 29344 9552 29408
rect 9616 29344 9632 29408
rect 9696 29344 9704 29408
rect 9384 28320 9704 29344
rect 9384 28256 9392 28320
rect 9456 28256 9472 28320
rect 9536 28256 9552 28320
rect 9616 28256 9632 28320
rect 9696 28256 9704 28320
rect 9384 27232 9704 28256
rect 9384 27168 9392 27232
rect 9456 27168 9472 27232
rect 9536 27168 9552 27232
rect 9616 27168 9632 27232
rect 9696 27168 9704 27232
rect 9384 26144 9704 27168
rect 9384 26080 9392 26144
rect 9456 26080 9472 26144
rect 9536 26080 9552 26144
rect 9616 26080 9632 26144
rect 9696 26080 9704 26144
rect 9384 25056 9704 26080
rect 9384 24992 9392 25056
rect 9456 24992 9472 25056
rect 9536 24992 9552 25056
rect 9616 24992 9632 25056
rect 9696 24992 9704 25056
rect 9384 23968 9704 24992
rect 9384 23904 9392 23968
rect 9456 23904 9472 23968
rect 9536 23904 9552 23968
rect 9616 23904 9632 23968
rect 9696 23904 9704 23968
rect 9384 22880 9704 23904
rect 9384 22816 9392 22880
rect 9456 22816 9472 22880
rect 9536 22816 9552 22880
rect 9616 22816 9632 22880
rect 9696 22816 9704 22880
rect 9384 21792 9704 22816
rect 9384 21728 9392 21792
rect 9456 21728 9472 21792
rect 9536 21728 9552 21792
rect 9616 21728 9632 21792
rect 9696 21728 9704 21792
rect 9384 20704 9704 21728
rect 9384 20640 9392 20704
rect 9456 20640 9472 20704
rect 9536 20640 9552 20704
rect 9616 20640 9632 20704
rect 9696 20640 9704 20704
rect 9384 19616 9704 20640
rect 9384 19552 9392 19616
rect 9456 19552 9472 19616
rect 9536 19552 9552 19616
rect 9616 19552 9632 19616
rect 9696 19552 9704 19616
rect 9384 18528 9704 19552
rect 9384 18464 9392 18528
rect 9456 18464 9472 18528
rect 9536 18464 9552 18528
rect 9616 18464 9632 18528
rect 9696 18464 9704 18528
rect 9384 17440 9704 18464
rect 9384 17376 9392 17440
rect 9456 17376 9472 17440
rect 9536 17376 9552 17440
rect 9616 17376 9632 17440
rect 9696 17376 9704 17440
rect 9384 16352 9704 17376
rect 9384 16288 9392 16352
rect 9456 16288 9472 16352
rect 9536 16288 9552 16352
rect 9616 16288 9632 16352
rect 9696 16288 9704 16352
rect 9384 15264 9704 16288
rect 9384 15200 9392 15264
rect 9456 15200 9472 15264
rect 9536 15200 9552 15264
rect 9616 15200 9632 15264
rect 9696 15200 9704 15264
rect 9384 14176 9704 15200
rect 9384 14112 9392 14176
rect 9456 14112 9472 14176
rect 9536 14112 9552 14176
rect 9616 14112 9632 14176
rect 9696 14112 9704 14176
rect 9384 13088 9704 14112
rect 9384 13024 9392 13088
rect 9456 13024 9472 13088
rect 9536 13024 9552 13088
rect 9616 13024 9632 13088
rect 9696 13024 9704 13088
rect 9384 12000 9704 13024
rect 9384 11936 9392 12000
rect 9456 11936 9472 12000
rect 9536 11936 9552 12000
rect 9616 11936 9632 12000
rect 9696 11936 9704 12000
rect 9384 10912 9704 11936
rect 9384 10848 9392 10912
rect 9456 10848 9472 10912
rect 9536 10848 9552 10912
rect 9616 10848 9632 10912
rect 9696 10848 9704 10912
rect 9384 9824 9704 10848
rect 9384 9760 9392 9824
rect 9456 9760 9472 9824
rect 9536 9760 9552 9824
rect 9616 9760 9632 9824
rect 9696 9760 9704 9824
rect 9384 8736 9704 9760
rect 9384 8672 9392 8736
rect 9456 8672 9472 8736
rect 9536 8672 9552 8736
rect 9616 8672 9632 8736
rect 9696 8672 9704 8736
rect 9384 7648 9704 8672
rect 9384 7584 9392 7648
rect 9456 7584 9472 7648
rect 9536 7584 9552 7648
rect 9616 7584 9632 7648
rect 9696 7584 9704 7648
rect 9384 6560 9704 7584
rect 9384 6496 9392 6560
rect 9456 6496 9472 6560
rect 9536 6496 9552 6560
rect 9616 6496 9632 6560
rect 9696 6496 9704 6560
rect 9384 5472 9704 6496
rect 9384 5408 9392 5472
rect 9456 5408 9472 5472
rect 9536 5408 9552 5472
rect 9616 5408 9632 5472
rect 9696 5408 9704 5472
rect 9384 4384 9704 5408
rect 9384 4320 9392 4384
rect 9456 4320 9472 4384
rect 9536 4320 9552 4384
rect 9616 4320 9632 4384
rect 9696 4320 9704 4384
rect 9384 3296 9704 4320
rect 9384 3232 9392 3296
rect 9456 3232 9472 3296
rect 9536 3232 9552 3296
rect 9616 3232 9632 3296
rect 9696 3232 9704 3296
rect 9384 2208 9704 3232
rect 9384 2144 9392 2208
rect 9456 2144 9472 2208
rect 9536 2144 9552 2208
rect 9616 2144 9632 2208
rect 9696 2144 9704 2208
rect 9384 2128 9704 2144
rect 13605 39744 13925 39760
rect 13605 39680 13613 39744
rect 13677 39680 13693 39744
rect 13757 39680 13773 39744
rect 13837 39680 13853 39744
rect 13917 39680 13925 39744
rect 13605 38656 13925 39680
rect 13605 38592 13613 38656
rect 13677 38592 13693 38656
rect 13757 38592 13773 38656
rect 13837 38592 13853 38656
rect 13917 38592 13925 38656
rect 13605 37568 13925 38592
rect 13605 37504 13613 37568
rect 13677 37504 13693 37568
rect 13757 37504 13773 37568
rect 13837 37504 13853 37568
rect 13917 37504 13925 37568
rect 13605 36480 13925 37504
rect 13605 36416 13613 36480
rect 13677 36416 13693 36480
rect 13757 36416 13773 36480
rect 13837 36416 13853 36480
rect 13917 36416 13925 36480
rect 13605 35392 13925 36416
rect 13605 35328 13613 35392
rect 13677 35328 13693 35392
rect 13757 35328 13773 35392
rect 13837 35328 13853 35392
rect 13917 35328 13925 35392
rect 13605 34304 13925 35328
rect 13605 34240 13613 34304
rect 13677 34240 13693 34304
rect 13757 34240 13773 34304
rect 13837 34240 13853 34304
rect 13917 34240 13925 34304
rect 13605 33216 13925 34240
rect 13605 33152 13613 33216
rect 13677 33152 13693 33216
rect 13757 33152 13773 33216
rect 13837 33152 13853 33216
rect 13917 33152 13925 33216
rect 13605 32128 13925 33152
rect 13605 32064 13613 32128
rect 13677 32064 13693 32128
rect 13757 32064 13773 32128
rect 13837 32064 13853 32128
rect 13917 32064 13925 32128
rect 13605 31040 13925 32064
rect 13605 30976 13613 31040
rect 13677 30976 13693 31040
rect 13757 30976 13773 31040
rect 13837 30976 13853 31040
rect 13917 30976 13925 31040
rect 13605 29952 13925 30976
rect 13605 29888 13613 29952
rect 13677 29888 13693 29952
rect 13757 29888 13773 29952
rect 13837 29888 13853 29952
rect 13917 29888 13925 29952
rect 13605 28864 13925 29888
rect 13605 28800 13613 28864
rect 13677 28800 13693 28864
rect 13757 28800 13773 28864
rect 13837 28800 13853 28864
rect 13917 28800 13925 28864
rect 13605 27776 13925 28800
rect 13605 27712 13613 27776
rect 13677 27712 13693 27776
rect 13757 27712 13773 27776
rect 13837 27712 13853 27776
rect 13917 27712 13925 27776
rect 13605 26688 13925 27712
rect 13605 26624 13613 26688
rect 13677 26624 13693 26688
rect 13757 26624 13773 26688
rect 13837 26624 13853 26688
rect 13917 26624 13925 26688
rect 13605 25600 13925 26624
rect 13605 25536 13613 25600
rect 13677 25536 13693 25600
rect 13757 25536 13773 25600
rect 13837 25536 13853 25600
rect 13917 25536 13925 25600
rect 13605 24512 13925 25536
rect 13605 24448 13613 24512
rect 13677 24448 13693 24512
rect 13757 24448 13773 24512
rect 13837 24448 13853 24512
rect 13917 24448 13925 24512
rect 13605 23424 13925 24448
rect 13605 23360 13613 23424
rect 13677 23360 13693 23424
rect 13757 23360 13773 23424
rect 13837 23360 13853 23424
rect 13917 23360 13925 23424
rect 13605 22336 13925 23360
rect 13605 22272 13613 22336
rect 13677 22272 13693 22336
rect 13757 22272 13773 22336
rect 13837 22272 13853 22336
rect 13917 22272 13925 22336
rect 13605 21248 13925 22272
rect 13605 21184 13613 21248
rect 13677 21184 13693 21248
rect 13757 21184 13773 21248
rect 13837 21184 13853 21248
rect 13917 21184 13925 21248
rect 13605 20160 13925 21184
rect 13605 20096 13613 20160
rect 13677 20096 13693 20160
rect 13757 20096 13773 20160
rect 13837 20096 13853 20160
rect 13917 20096 13925 20160
rect 13605 19072 13925 20096
rect 13605 19008 13613 19072
rect 13677 19008 13693 19072
rect 13757 19008 13773 19072
rect 13837 19008 13853 19072
rect 13917 19008 13925 19072
rect 13605 17984 13925 19008
rect 13605 17920 13613 17984
rect 13677 17920 13693 17984
rect 13757 17920 13773 17984
rect 13837 17920 13853 17984
rect 13917 17920 13925 17984
rect 13605 16896 13925 17920
rect 13605 16832 13613 16896
rect 13677 16832 13693 16896
rect 13757 16832 13773 16896
rect 13837 16832 13853 16896
rect 13917 16832 13925 16896
rect 13605 15808 13925 16832
rect 13605 15744 13613 15808
rect 13677 15744 13693 15808
rect 13757 15744 13773 15808
rect 13837 15744 13853 15808
rect 13917 15744 13925 15808
rect 13605 14720 13925 15744
rect 13605 14656 13613 14720
rect 13677 14656 13693 14720
rect 13757 14656 13773 14720
rect 13837 14656 13853 14720
rect 13917 14656 13925 14720
rect 13605 13632 13925 14656
rect 13605 13568 13613 13632
rect 13677 13568 13693 13632
rect 13757 13568 13773 13632
rect 13837 13568 13853 13632
rect 13917 13568 13925 13632
rect 13605 12544 13925 13568
rect 13605 12480 13613 12544
rect 13677 12480 13693 12544
rect 13757 12480 13773 12544
rect 13837 12480 13853 12544
rect 13917 12480 13925 12544
rect 13605 11456 13925 12480
rect 13605 11392 13613 11456
rect 13677 11392 13693 11456
rect 13757 11392 13773 11456
rect 13837 11392 13853 11456
rect 13917 11392 13925 11456
rect 13605 10368 13925 11392
rect 13605 10304 13613 10368
rect 13677 10304 13693 10368
rect 13757 10304 13773 10368
rect 13837 10304 13853 10368
rect 13917 10304 13925 10368
rect 13605 9280 13925 10304
rect 13605 9216 13613 9280
rect 13677 9216 13693 9280
rect 13757 9216 13773 9280
rect 13837 9216 13853 9280
rect 13917 9216 13925 9280
rect 13605 8192 13925 9216
rect 13605 8128 13613 8192
rect 13677 8128 13693 8192
rect 13757 8128 13773 8192
rect 13837 8128 13853 8192
rect 13917 8128 13925 8192
rect 13605 7104 13925 8128
rect 13605 7040 13613 7104
rect 13677 7040 13693 7104
rect 13757 7040 13773 7104
rect 13837 7040 13853 7104
rect 13917 7040 13925 7104
rect 13605 6016 13925 7040
rect 13605 5952 13613 6016
rect 13677 5952 13693 6016
rect 13757 5952 13773 6016
rect 13837 5952 13853 6016
rect 13917 5952 13925 6016
rect 13605 4928 13925 5952
rect 13605 4864 13613 4928
rect 13677 4864 13693 4928
rect 13757 4864 13773 4928
rect 13837 4864 13853 4928
rect 13917 4864 13925 4928
rect 13605 3840 13925 4864
rect 13605 3776 13613 3840
rect 13677 3776 13693 3840
rect 13757 3776 13773 3840
rect 13837 3776 13853 3840
rect 13917 3776 13925 3840
rect 13605 2752 13925 3776
rect 13605 2688 13613 2752
rect 13677 2688 13693 2752
rect 13757 2688 13773 2752
rect 13837 2688 13853 2752
rect 13917 2688 13925 2752
rect 13605 2128 13925 2688
rect 17825 39200 18145 39760
rect 17825 39136 17833 39200
rect 17897 39136 17913 39200
rect 17977 39136 17993 39200
rect 18057 39136 18073 39200
rect 18137 39136 18145 39200
rect 17825 38112 18145 39136
rect 17825 38048 17833 38112
rect 17897 38048 17913 38112
rect 17977 38048 17993 38112
rect 18057 38048 18073 38112
rect 18137 38048 18145 38112
rect 17825 37024 18145 38048
rect 17825 36960 17833 37024
rect 17897 36960 17913 37024
rect 17977 36960 17993 37024
rect 18057 36960 18073 37024
rect 18137 36960 18145 37024
rect 17825 35936 18145 36960
rect 17825 35872 17833 35936
rect 17897 35872 17913 35936
rect 17977 35872 17993 35936
rect 18057 35872 18073 35936
rect 18137 35872 18145 35936
rect 17825 34848 18145 35872
rect 17825 34784 17833 34848
rect 17897 34784 17913 34848
rect 17977 34784 17993 34848
rect 18057 34784 18073 34848
rect 18137 34784 18145 34848
rect 17825 33760 18145 34784
rect 17825 33696 17833 33760
rect 17897 33696 17913 33760
rect 17977 33696 17993 33760
rect 18057 33696 18073 33760
rect 18137 33696 18145 33760
rect 17825 32672 18145 33696
rect 17825 32608 17833 32672
rect 17897 32608 17913 32672
rect 17977 32608 17993 32672
rect 18057 32608 18073 32672
rect 18137 32608 18145 32672
rect 17825 31584 18145 32608
rect 17825 31520 17833 31584
rect 17897 31520 17913 31584
rect 17977 31520 17993 31584
rect 18057 31520 18073 31584
rect 18137 31520 18145 31584
rect 17825 30496 18145 31520
rect 17825 30432 17833 30496
rect 17897 30432 17913 30496
rect 17977 30432 17993 30496
rect 18057 30432 18073 30496
rect 18137 30432 18145 30496
rect 17825 29408 18145 30432
rect 17825 29344 17833 29408
rect 17897 29344 17913 29408
rect 17977 29344 17993 29408
rect 18057 29344 18073 29408
rect 18137 29344 18145 29408
rect 17825 28320 18145 29344
rect 17825 28256 17833 28320
rect 17897 28256 17913 28320
rect 17977 28256 17993 28320
rect 18057 28256 18073 28320
rect 18137 28256 18145 28320
rect 17825 27232 18145 28256
rect 17825 27168 17833 27232
rect 17897 27168 17913 27232
rect 17977 27168 17993 27232
rect 18057 27168 18073 27232
rect 18137 27168 18145 27232
rect 17825 26144 18145 27168
rect 17825 26080 17833 26144
rect 17897 26080 17913 26144
rect 17977 26080 17993 26144
rect 18057 26080 18073 26144
rect 18137 26080 18145 26144
rect 17825 25056 18145 26080
rect 17825 24992 17833 25056
rect 17897 24992 17913 25056
rect 17977 24992 17993 25056
rect 18057 24992 18073 25056
rect 18137 24992 18145 25056
rect 17825 23968 18145 24992
rect 17825 23904 17833 23968
rect 17897 23904 17913 23968
rect 17977 23904 17993 23968
rect 18057 23904 18073 23968
rect 18137 23904 18145 23968
rect 17825 22880 18145 23904
rect 17825 22816 17833 22880
rect 17897 22816 17913 22880
rect 17977 22816 17993 22880
rect 18057 22816 18073 22880
rect 18137 22816 18145 22880
rect 17825 21792 18145 22816
rect 17825 21728 17833 21792
rect 17897 21728 17913 21792
rect 17977 21728 17993 21792
rect 18057 21728 18073 21792
rect 18137 21728 18145 21792
rect 17825 20704 18145 21728
rect 17825 20640 17833 20704
rect 17897 20640 17913 20704
rect 17977 20640 17993 20704
rect 18057 20640 18073 20704
rect 18137 20640 18145 20704
rect 17825 19616 18145 20640
rect 17825 19552 17833 19616
rect 17897 19552 17913 19616
rect 17977 19552 17993 19616
rect 18057 19552 18073 19616
rect 18137 19552 18145 19616
rect 17825 18528 18145 19552
rect 17825 18464 17833 18528
rect 17897 18464 17913 18528
rect 17977 18464 17993 18528
rect 18057 18464 18073 18528
rect 18137 18464 18145 18528
rect 17825 17440 18145 18464
rect 17825 17376 17833 17440
rect 17897 17376 17913 17440
rect 17977 17376 17993 17440
rect 18057 17376 18073 17440
rect 18137 17376 18145 17440
rect 17825 16352 18145 17376
rect 17825 16288 17833 16352
rect 17897 16288 17913 16352
rect 17977 16288 17993 16352
rect 18057 16288 18073 16352
rect 18137 16288 18145 16352
rect 17825 15264 18145 16288
rect 17825 15200 17833 15264
rect 17897 15200 17913 15264
rect 17977 15200 17993 15264
rect 18057 15200 18073 15264
rect 18137 15200 18145 15264
rect 17825 14176 18145 15200
rect 17825 14112 17833 14176
rect 17897 14112 17913 14176
rect 17977 14112 17993 14176
rect 18057 14112 18073 14176
rect 18137 14112 18145 14176
rect 17825 13088 18145 14112
rect 17825 13024 17833 13088
rect 17897 13024 17913 13088
rect 17977 13024 17993 13088
rect 18057 13024 18073 13088
rect 18137 13024 18145 13088
rect 17825 12000 18145 13024
rect 17825 11936 17833 12000
rect 17897 11936 17913 12000
rect 17977 11936 17993 12000
rect 18057 11936 18073 12000
rect 18137 11936 18145 12000
rect 17825 10912 18145 11936
rect 17825 10848 17833 10912
rect 17897 10848 17913 10912
rect 17977 10848 17993 10912
rect 18057 10848 18073 10912
rect 18137 10848 18145 10912
rect 17825 9824 18145 10848
rect 17825 9760 17833 9824
rect 17897 9760 17913 9824
rect 17977 9760 17993 9824
rect 18057 9760 18073 9824
rect 18137 9760 18145 9824
rect 17825 8736 18145 9760
rect 17825 8672 17833 8736
rect 17897 8672 17913 8736
rect 17977 8672 17993 8736
rect 18057 8672 18073 8736
rect 18137 8672 18145 8736
rect 17825 7648 18145 8672
rect 17825 7584 17833 7648
rect 17897 7584 17913 7648
rect 17977 7584 17993 7648
rect 18057 7584 18073 7648
rect 18137 7584 18145 7648
rect 17825 6560 18145 7584
rect 17825 6496 17833 6560
rect 17897 6496 17913 6560
rect 17977 6496 17993 6560
rect 18057 6496 18073 6560
rect 18137 6496 18145 6560
rect 17825 5472 18145 6496
rect 17825 5408 17833 5472
rect 17897 5408 17913 5472
rect 17977 5408 17993 5472
rect 18057 5408 18073 5472
rect 18137 5408 18145 5472
rect 17825 4384 18145 5408
rect 17825 4320 17833 4384
rect 17897 4320 17913 4384
rect 17977 4320 17993 4384
rect 18057 4320 18073 4384
rect 18137 4320 18145 4384
rect 17825 3296 18145 4320
rect 17825 3232 17833 3296
rect 17897 3232 17913 3296
rect 17977 3232 17993 3296
rect 18057 3232 18073 3296
rect 18137 3232 18145 3296
rect 17825 2208 18145 3232
rect 17825 2144 17833 2208
rect 17897 2144 17913 2208
rect 17977 2144 17993 2208
rect 18057 2144 18073 2208
rect 18137 2144 18145 2208
rect 17825 2128 18145 2144
rect 22046 39744 22366 39760
rect 22046 39680 22054 39744
rect 22118 39680 22134 39744
rect 22198 39680 22214 39744
rect 22278 39680 22294 39744
rect 22358 39680 22366 39744
rect 22046 38656 22366 39680
rect 22046 38592 22054 38656
rect 22118 38592 22134 38656
rect 22198 38592 22214 38656
rect 22278 38592 22294 38656
rect 22358 38592 22366 38656
rect 22046 37568 22366 38592
rect 22046 37504 22054 37568
rect 22118 37504 22134 37568
rect 22198 37504 22214 37568
rect 22278 37504 22294 37568
rect 22358 37504 22366 37568
rect 22046 36480 22366 37504
rect 22046 36416 22054 36480
rect 22118 36416 22134 36480
rect 22198 36416 22214 36480
rect 22278 36416 22294 36480
rect 22358 36416 22366 36480
rect 22046 35392 22366 36416
rect 22046 35328 22054 35392
rect 22118 35328 22134 35392
rect 22198 35328 22214 35392
rect 22278 35328 22294 35392
rect 22358 35328 22366 35392
rect 22046 34304 22366 35328
rect 22046 34240 22054 34304
rect 22118 34240 22134 34304
rect 22198 34240 22214 34304
rect 22278 34240 22294 34304
rect 22358 34240 22366 34304
rect 22046 33216 22366 34240
rect 22046 33152 22054 33216
rect 22118 33152 22134 33216
rect 22198 33152 22214 33216
rect 22278 33152 22294 33216
rect 22358 33152 22366 33216
rect 22046 32128 22366 33152
rect 22046 32064 22054 32128
rect 22118 32064 22134 32128
rect 22198 32064 22214 32128
rect 22278 32064 22294 32128
rect 22358 32064 22366 32128
rect 22046 31040 22366 32064
rect 22046 30976 22054 31040
rect 22118 30976 22134 31040
rect 22198 30976 22214 31040
rect 22278 30976 22294 31040
rect 22358 30976 22366 31040
rect 22046 29952 22366 30976
rect 22046 29888 22054 29952
rect 22118 29888 22134 29952
rect 22198 29888 22214 29952
rect 22278 29888 22294 29952
rect 22358 29888 22366 29952
rect 22046 28864 22366 29888
rect 22046 28800 22054 28864
rect 22118 28800 22134 28864
rect 22198 28800 22214 28864
rect 22278 28800 22294 28864
rect 22358 28800 22366 28864
rect 22046 27776 22366 28800
rect 22046 27712 22054 27776
rect 22118 27712 22134 27776
rect 22198 27712 22214 27776
rect 22278 27712 22294 27776
rect 22358 27712 22366 27776
rect 22046 26688 22366 27712
rect 22046 26624 22054 26688
rect 22118 26624 22134 26688
rect 22198 26624 22214 26688
rect 22278 26624 22294 26688
rect 22358 26624 22366 26688
rect 22046 25600 22366 26624
rect 22046 25536 22054 25600
rect 22118 25536 22134 25600
rect 22198 25536 22214 25600
rect 22278 25536 22294 25600
rect 22358 25536 22366 25600
rect 22046 24512 22366 25536
rect 22046 24448 22054 24512
rect 22118 24448 22134 24512
rect 22198 24448 22214 24512
rect 22278 24448 22294 24512
rect 22358 24448 22366 24512
rect 22046 23424 22366 24448
rect 22046 23360 22054 23424
rect 22118 23360 22134 23424
rect 22198 23360 22214 23424
rect 22278 23360 22294 23424
rect 22358 23360 22366 23424
rect 22046 22336 22366 23360
rect 22046 22272 22054 22336
rect 22118 22272 22134 22336
rect 22198 22272 22214 22336
rect 22278 22272 22294 22336
rect 22358 22272 22366 22336
rect 22046 21248 22366 22272
rect 22046 21184 22054 21248
rect 22118 21184 22134 21248
rect 22198 21184 22214 21248
rect 22278 21184 22294 21248
rect 22358 21184 22366 21248
rect 22046 20160 22366 21184
rect 22046 20096 22054 20160
rect 22118 20096 22134 20160
rect 22198 20096 22214 20160
rect 22278 20096 22294 20160
rect 22358 20096 22366 20160
rect 22046 19072 22366 20096
rect 22046 19008 22054 19072
rect 22118 19008 22134 19072
rect 22198 19008 22214 19072
rect 22278 19008 22294 19072
rect 22358 19008 22366 19072
rect 22046 17984 22366 19008
rect 22046 17920 22054 17984
rect 22118 17920 22134 17984
rect 22198 17920 22214 17984
rect 22278 17920 22294 17984
rect 22358 17920 22366 17984
rect 22046 16896 22366 17920
rect 22046 16832 22054 16896
rect 22118 16832 22134 16896
rect 22198 16832 22214 16896
rect 22278 16832 22294 16896
rect 22358 16832 22366 16896
rect 22046 15808 22366 16832
rect 22046 15744 22054 15808
rect 22118 15744 22134 15808
rect 22198 15744 22214 15808
rect 22278 15744 22294 15808
rect 22358 15744 22366 15808
rect 22046 14720 22366 15744
rect 22046 14656 22054 14720
rect 22118 14656 22134 14720
rect 22198 14656 22214 14720
rect 22278 14656 22294 14720
rect 22358 14656 22366 14720
rect 22046 13632 22366 14656
rect 22046 13568 22054 13632
rect 22118 13568 22134 13632
rect 22198 13568 22214 13632
rect 22278 13568 22294 13632
rect 22358 13568 22366 13632
rect 22046 12544 22366 13568
rect 22046 12480 22054 12544
rect 22118 12480 22134 12544
rect 22198 12480 22214 12544
rect 22278 12480 22294 12544
rect 22358 12480 22366 12544
rect 22046 11456 22366 12480
rect 22046 11392 22054 11456
rect 22118 11392 22134 11456
rect 22198 11392 22214 11456
rect 22278 11392 22294 11456
rect 22358 11392 22366 11456
rect 22046 10368 22366 11392
rect 22046 10304 22054 10368
rect 22118 10304 22134 10368
rect 22198 10304 22214 10368
rect 22278 10304 22294 10368
rect 22358 10304 22366 10368
rect 22046 9280 22366 10304
rect 22046 9216 22054 9280
rect 22118 9216 22134 9280
rect 22198 9216 22214 9280
rect 22278 9216 22294 9280
rect 22358 9216 22366 9280
rect 22046 8192 22366 9216
rect 22046 8128 22054 8192
rect 22118 8128 22134 8192
rect 22198 8128 22214 8192
rect 22278 8128 22294 8192
rect 22358 8128 22366 8192
rect 22046 7104 22366 8128
rect 22046 7040 22054 7104
rect 22118 7040 22134 7104
rect 22198 7040 22214 7104
rect 22278 7040 22294 7104
rect 22358 7040 22366 7104
rect 22046 6016 22366 7040
rect 22046 5952 22054 6016
rect 22118 5952 22134 6016
rect 22198 5952 22214 6016
rect 22278 5952 22294 6016
rect 22358 5952 22366 6016
rect 22046 4928 22366 5952
rect 22046 4864 22054 4928
rect 22118 4864 22134 4928
rect 22198 4864 22214 4928
rect 22278 4864 22294 4928
rect 22358 4864 22366 4928
rect 22046 3840 22366 4864
rect 22046 3776 22054 3840
rect 22118 3776 22134 3840
rect 22198 3776 22214 3840
rect 22278 3776 22294 3840
rect 22358 3776 22366 3840
rect 22046 2752 22366 3776
rect 22046 2688 22054 2752
rect 22118 2688 22134 2752
rect 22198 2688 22214 2752
rect 22278 2688 22294 2752
rect 22358 2688 22366 2752
rect 22046 2128 22366 2688
rect 26266 39200 26586 39760
rect 26266 39136 26274 39200
rect 26338 39136 26354 39200
rect 26418 39136 26434 39200
rect 26498 39136 26514 39200
rect 26578 39136 26586 39200
rect 26266 38112 26586 39136
rect 26266 38048 26274 38112
rect 26338 38048 26354 38112
rect 26418 38048 26434 38112
rect 26498 38048 26514 38112
rect 26578 38048 26586 38112
rect 26266 37024 26586 38048
rect 26266 36960 26274 37024
rect 26338 36960 26354 37024
rect 26418 36960 26434 37024
rect 26498 36960 26514 37024
rect 26578 36960 26586 37024
rect 26266 35936 26586 36960
rect 26266 35872 26274 35936
rect 26338 35872 26354 35936
rect 26418 35872 26434 35936
rect 26498 35872 26514 35936
rect 26578 35872 26586 35936
rect 26266 34848 26586 35872
rect 26266 34784 26274 34848
rect 26338 34784 26354 34848
rect 26418 34784 26434 34848
rect 26498 34784 26514 34848
rect 26578 34784 26586 34848
rect 26266 33760 26586 34784
rect 26266 33696 26274 33760
rect 26338 33696 26354 33760
rect 26418 33696 26434 33760
rect 26498 33696 26514 33760
rect 26578 33696 26586 33760
rect 26266 32672 26586 33696
rect 26266 32608 26274 32672
rect 26338 32608 26354 32672
rect 26418 32608 26434 32672
rect 26498 32608 26514 32672
rect 26578 32608 26586 32672
rect 26266 31584 26586 32608
rect 26266 31520 26274 31584
rect 26338 31520 26354 31584
rect 26418 31520 26434 31584
rect 26498 31520 26514 31584
rect 26578 31520 26586 31584
rect 26266 30496 26586 31520
rect 26266 30432 26274 30496
rect 26338 30432 26354 30496
rect 26418 30432 26434 30496
rect 26498 30432 26514 30496
rect 26578 30432 26586 30496
rect 26266 29408 26586 30432
rect 26266 29344 26274 29408
rect 26338 29344 26354 29408
rect 26418 29344 26434 29408
rect 26498 29344 26514 29408
rect 26578 29344 26586 29408
rect 26266 28320 26586 29344
rect 26266 28256 26274 28320
rect 26338 28256 26354 28320
rect 26418 28256 26434 28320
rect 26498 28256 26514 28320
rect 26578 28256 26586 28320
rect 26266 27232 26586 28256
rect 26266 27168 26274 27232
rect 26338 27168 26354 27232
rect 26418 27168 26434 27232
rect 26498 27168 26514 27232
rect 26578 27168 26586 27232
rect 26266 26144 26586 27168
rect 26266 26080 26274 26144
rect 26338 26080 26354 26144
rect 26418 26080 26434 26144
rect 26498 26080 26514 26144
rect 26578 26080 26586 26144
rect 26266 25056 26586 26080
rect 26266 24992 26274 25056
rect 26338 24992 26354 25056
rect 26418 24992 26434 25056
rect 26498 24992 26514 25056
rect 26578 24992 26586 25056
rect 26266 23968 26586 24992
rect 26266 23904 26274 23968
rect 26338 23904 26354 23968
rect 26418 23904 26434 23968
rect 26498 23904 26514 23968
rect 26578 23904 26586 23968
rect 26266 22880 26586 23904
rect 26266 22816 26274 22880
rect 26338 22816 26354 22880
rect 26418 22816 26434 22880
rect 26498 22816 26514 22880
rect 26578 22816 26586 22880
rect 26266 21792 26586 22816
rect 26266 21728 26274 21792
rect 26338 21728 26354 21792
rect 26418 21728 26434 21792
rect 26498 21728 26514 21792
rect 26578 21728 26586 21792
rect 26266 20704 26586 21728
rect 26266 20640 26274 20704
rect 26338 20640 26354 20704
rect 26418 20640 26434 20704
rect 26498 20640 26514 20704
rect 26578 20640 26586 20704
rect 26266 19616 26586 20640
rect 26266 19552 26274 19616
rect 26338 19552 26354 19616
rect 26418 19552 26434 19616
rect 26498 19552 26514 19616
rect 26578 19552 26586 19616
rect 26266 18528 26586 19552
rect 26266 18464 26274 18528
rect 26338 18464 26354 18528
rect 26418 18464 26434 18528
rect 26498 18464 26514 18528
rect 26578 18464 26586 18528
rect 26266 17440 26586 18464
rect 26266 17376 26274 17440
rect 26338 17376 26354 17440
rect 26418 17376 26434 17440
rect 26498 17376 26514 17440
rect 26578 17376 26586 17440
rect 26266 16352 26586 17376
rect 26266 16288 26274 16352
rect 26338 16288 26354 16352
rect 26418 16288 26434 16352
rect 26498 16288 26514 16352
rect 26578 16288 26586 16352
rect 26266 15264 26586 16288
rect 26266 15200 26274 15264
rect 26338 15200 26354 15264
rect 26418 15200 26434 15264
rect 26498 15200 26514 15264
rect 26578 15200 26586 15264
rect 26266 14176 26586 15200
rect 26266 14112 26274 14176
rect 26338 14112 26354 14176
rect 26418 14112 26434 14176
rect 26498 14112 26514 14176
rect 26578 14112 26586 14176
rect 26266 13088 26586 14112
rect 26266 13024 26274 13088
rect 26338 13024 26354 13088
rect 26418 13024 26434 13088
rect 26498 13024 26514 13088
rect 26578 13024 26586 13088
rect 26266 12000 26586 13024
rect 26266 11936 26274 12000
rect 26338 11936 26354 12000
rect 26418 11936 26434 12000
rect 26498 11936 26514 12000
rect 26578 11936 26586 12000
rect 26266 10912 26586 11936
rect 26266 10848 26274 10912
rect 26338 10848 26354 10912
rect 26418 10848 26434 10912
rect 26498 10848 26514 10912
rect 26578 10848 26586 10912
rect 26266 9824 26586 10848
rect 26266 9760 26274 9824
rect 26338 9760 26354 9824
rect 26418 9760 26434 9824
rect 26498 9760 26514 9824
rect 26578 9760 26586 9824
rect 26266 8736 26586 9760
rect 26266 8672 26274 8736
rect 26338 8672 26354 8736
rect 26418 8672 26434 8736
rect 26498 8672 26514 8736
rect 26578 8672 26586 8736
rect 26266 7648 26586 8672
rect 26266 7584 26274 7648
rect 26338 7584 26354 7648
rect 26418 7584 26434 7648
rect 26498 7584 26514 7648
rect 26578 7584 26586 7648
rect 26266 6560 26586 7584
rect 26266 6496 26274 6560
rect 26338 6496 26354 6560
rect 26418 6496 26434 6560
rect 26498 6496 26514 6560
rect 26578 6496 26586 6560
rect 26266 5472 26586 6496
rect 26266 5408 26274 5472
rect 26338 5408 26354 5472
rect 26418 5408 26434 5472
rect 26498 5408 26514 5472
rect 26578 5408 26586 5472
rect 26266 4384 26586 5408
rect 26266 4320 26274 4384
rect 26338 4320 26354 4384
rect 26418 4320 26434 4384
rect 26498 4320 26514 4384
rect 26578 4320 26586 4384
rect 26266 3296 26586 4320
rect 26266 3232 26274 3296
rect 26338 3232 26354 3296
rect 26418 3232 26434 3296
rect 26498 3232 26514 3296
rect 26578 3232 26586 3296
rect 26266 2208 26586 3232
rect 26266 2144 26274 2208
rect 26338 2144 26354 2208
rect 26418 2144 26434 2208
rect 26498 2144 26514 2208
rect 26578 2144 26586 2208
rect 26266 2128 26586 2144
rect 30487 39744 30807 39760
rect 30487 39680 30495 39744
rect 30559 39680 30575 39744
rect 30639 39680 30655 39744
rect 30719 39680 30735 39744
rect 30799 39680 30807 39744
rect 30487 38656 30807 39680
rect 30487 38592 30495 38656
rect 30559 38592 30575 38656
rect 30639 38592 30655 38656
rect 30719 38592 30735 38656
rect 30799 38592 30807 38656
rect 30487 37568 30807 38592
rect 30487 37504 30495 37568
rect 30559 37504 30575 37568
rect 30639 37504 30655 37568
rect 30719 37504 30735 37568
rect 30799 37504 30807 37568
rect 30487 36480 30807 37504
rect 30487 36416 30495 36480
rect 30559 36416 30575 36480
rect 30639 36416 30655 36480
rect 30719 36416 30735 36480
rect 30799 36416 30807 36480
rect 30487 35392 30807 36416
rect 30487 35328 30495 35392
rect 30559 35328 30575 35392
rect 30639 35328 30655 35392
rect 30719 35328 30735 35392
rect 30799 35328 30807 35392
rect 30487 34304 30807 35328
rect 30487 34240 30495 34304
rect 30559 34240 30575 34304
rect 30639 34240 30655 34304
rect 30719 34240 30735 34304
rect 30799 34240 30807 34304
rect 30487 33216 30807 34240
rect 30487 33152 30495 33216
rect 30559 33152 30575 33216
rect 30639 33152 30655 33216
rect 30719 33152 30735 33216
rect 30799 33152 30807 33216
rect 30487 32128 30807 33152
rect 30487 32064 30495 32128
rect 30559 32064 30575 32128
rect 30639 32064 30655 32128
rect 30719 32064 30735 32128
rect 30799 32064 30807 32128
rect 30487 31040 30807 32064
rect 30487 30976 30495 31040
rect 30559 30976 30575 31040
rect 30639 30976 30655 31040
rect 30719 30976 30735 31040
rect 30799 30976 30807 31040
rect 30487 29952 30807 30976
rect 30487 29888 30495 29952
rect 30559 29888 30575 29952
rect 30639 29888 30655 29952
rect 30719 29888 30735 29952
rect 30799 29888 30807 29952
rect 30487 28864 30807 29888
rect 30487 28800 30495 28864
rect 30559 28800 30575 28864
rect 30639 28800 30655 28864
rect 30719 28800 30735 28864
rect 30799 28800 30807 28864
rect 30487 27776 30807 28800
rect 30487 27712 30495 27776
rect 30559 27712 30575 27776
rect 30639 27712 30655 27776
rect 30719 27712 30735 27776
rect 30799 27712 30807 27776
rect 30487 26688 30807 27712
rect 30487 26624 30495 26688
rect 30559 26624 30575 26688
rect 30639 26624 30655 26688
rect 30719 26624 30735 26688
rect 30799 26624 30807 26688
rect 30487 25600 30807 26624
rect 30487 25536 30495 25600
rect 30559 25536 30575 25600
rect 30639 25536 30655 25600
rect 30719 25536 30735 25600
rect 30799 25536 30807 25600
rect 30487 24512 30807 25536
rect 30487 24448 30495 24512
rect 30559 24448 30575 24512
rect 30639 24448 30655 24512
rect 30719 24448 30735 24512
rect 30799 24448 30807 24512
rect 30487 23424 30807 24448
rect 30487 23360 30495 23424
rect 30559 23360 30575 23424
rect 30639 23360 30655 23424
rect 30719 23360 30735 23424
rect 30799 23360 30807 23424
rect 30487 22336 30807 23360
rect 30487 22272 30495 22336
rect 30559 22272 30575 22336
rect 30639 22272 30655 22336
rect 30719 22272 30735 22336
rect 30799 22272 30807 22336
rect 30487 21248 30807 22272
rect 30487 21184 30495 21248
rect 30559 21184 30575 21248
rect 30639 21184 30655 21248
rect 30719 21184 30735 21248
rect 30799 21184 30807 21248
rect 30487 20160 30807 21184
rect 30487 20096 30495 20160
rect 30559 20096 30575 20160
rect 30639 20096 30655 20160
rect 30719 20096 30735 20160
rect 30799 20096 30807 20160
rect 30487 19072 30807 20096
rect 30487 19008 30495 19072
rect 30559 19008 30575 19072
rect 30639 19008 30655 19072
rect 30719 19008 30735 19072
rect 30799 19008 30807 19072
rect 30487 17984 30807 19008
rect 30487 17920 30495 17984
rect 30559 17920 30575 17984
rect 30639 17920 30655 17984
rect 30719 17920 30735 17984
rect 30799 17920 30807 17984
rect 30487 16896 30807 17920
rect 30487 16832 30495 16896
rect 30559 16832 30575 16896
rect 30639 16832 30655 16896
rect 30719 16832 30735 16896
rect 30799 16832 30807 16896
rect 30487 15808 30807 16832
rect 30487 15744 30495 15808
rect 30559 15744 30575 15808
rect 30639 15744 30655 15808
rect 30719 15744 30735 15808
rect 30799 15744 30807 15808
rect 30487 14720 30807 15744
rect 30487 14656 30495 14720
rect 30559 14656 30575 14720
rect 30639 14656 30655 14720
rect 30719 14656 30735 14720
rect 30799 14656 30807 14720
rect 30487 13632 30807 14656
rect 30487 13568 30495 13632
rect 30559 13568 30575 13632
rect 30639 13568 30655 13632
rect 30719 13568 30735 13632
rect 30799 13568 30807 13632
rect 30487 12544 30807 13568
rect 30487 12480 30495 12544
rect 30559 12480 30575 12544
rect 30639 12480 30655 12544
rect 30719 12480 30735 12544
rect 30799 12480 30807 12544
rect 30487 11456 30807 12480
rect 30487 11392 30495 11456
rect 30559 11392 30575 11456
rect 30639 11392 30655 11456
rect 30719 11392 30735 11456
rect 30799 11392 30807 11456
rect 30487 10368 30807 11392
rect 30487 10304 30495 10368
rect 30559 10304 30575 10368
rect 30639 10304 30655 10368
rect 30719 10304 30735 10368
rect 30799 10304 30807 10368
rect 30487 9280 30807 10304
rect 30487 9216 30495 9280
rect 30559 9216 30575 9280
rect 30639 9216 30655 9280
rect 30719 9216 30735 9280
rect 30799 9216 30807 9280
rect 30487 8192 30807 9216
rect 30487 8128 30495 8192
rect 30559 8128 30575 8192
rect 30639 8128 30655 8192
rect 30719 8128 30735 8192
rect 30799 8128 30807 8192
rect 30487 7104 30807 8128
rect 30487 7040 30495 7104
rect 30559 7040 30575 7104
rect 30639 7040 30655 7104
rect 30719 7040 30735 7104
rect 30799 7040 30807 7104
rect 30487 6016 30807 7040
rect 30487 5952 30495 6016
rect 30559 5952 30575 6016
rect 30639 5952 30655 6016
rect 30719 5952 30735 6016
rect 30799 5952 30807 6016
rect 30487 4928 30807 5952
rect 30487 4864 30495 4928
rect 30559 4864 30575 4928
rect 30639 4864 30655 4928
rect 30719 4864 30735 4928
rect 30799 4864 30807 4928
rect 30487 3840 30807 4864
rect 30487 3776 30495 3840
rect 30559 3776 30575 3840
rect 30639 3776 30655 3840
rect 30719 3776 30735 3840
rect 30799 3776 30807 3840
rect 30487 2752 30807 3776
rect 30487 2688 30495 2752
rect 30559 2688 30575 2752
rect 30639 2688 30655 2752
rect 30719 2688 30735 2752
rect 30799 2688 30807 2752
rect 30487 2128 30807 2688
rect 34707 39200 35027 39760
rect 34707 39136 34715 39200
rect 34779 39136 34795 39200
rect 34859 39136 34875 39200
rect 34939 39136 34955 39200
rect 35019 39136 35027 39200
rect 34707 38112 35027 39136
rect 34707 38048 34715 38112
rect 34779 38048 34795 38112
rect 34859 38048 34875 38112
rect 34939 38048 34955 38112
rect 35019 38048 35027 38112
rect 34707 37024 35027 38048
rect 34707 36960 34715 37024
rect 34779 36960 34795 37024
rect 34859 36960 34875 37024
rect 34939 36960 34955 37024
rect 35019 36960 35027 37024
rect 34707 35936 35027 36960
rect 34707 35872 34715 35936
rect 34779 35872 34795 35936
rect 34859 35872 34875 35936
rect 34939 35872 34955 35936
rect 35019 35872 35027 35936
rect 34707 34848 35027 35872
rect 34707 34784 34715 34848
rect 34779 34784 34795 34848
rect 34859 34784 34875 34848
rect 34939 34784 34955 34848
rect 35019 34784 35027 34848
rect 34707 33760 35027 34784
rect 34707 33696 34715 33760
rect 34779 33696 34795 33760
rect 34859 33696 34875 33760
rect 34939 33696 34955 33760
rect 35019 33696 35027 33760
rect 34707 32672 35027 33696
rect 34707 32608 34715 32672
rect 34779 32608 34795 32672
rect 34859 32608 34875 32672
rect 34939 32608 34955 32672
rect 35019 32608 35027 32672
rect 34707 31584 35027 32608
rect 34707 31520 34715 31584
rect 34779 31520 34795 31584
rect 34859 31520 34875 31584
rect 34939 31520 34955 31584
rect 35019 31520 35027 31584
rect 34707 30496 35027 31520
rect 34707 30432 34715 30496
rect 34779 30432 34795 30496
rect 34859 30432 34875 30496
rect 34939 30432 34955 30496
rect 35019 30432 35027 30496
rect 34707 29408 35027 30432
rect 34707 29344 34715 29408
rect 34779 29344 34795 29408
rect 34859 29344 34875 29408
rect 34939 29344 34955 29408
rect 35019 29344 35027 29408
rect 34707 28320 35027 29344
rect 34707 28256 34715 28320
rect 34779 28256 34795 28320
rect 34859 28256 34875 28320
rect 34939 28256 34955 28320
rect 35019 28256 35027 28320
rect 34707 27232 35027 28256
rect 34707 27168 34715 27232
rect 34779 27168 34795 27232
rect 34859 27168 34875 27232
rect 34939 27168 34955 27232
rect 35019 27168 35027 27232
rect 34707 26144 35027 27168
rect 34707 26080 34715 26144
rect 34779 26080 34795 26144
rect 34859 26080 34875 26144
rect 34939 26080 34955 26144
rect 35019 26080 35027 26144
rect 34707 25056 35027 26080
rect 34707 24992 34715 25056
rect 34779 24992 34795 25056
rect 34859 24992 34875 25056
rect 34939 24992 34955 25056
rect 35019 24992 35027 25056
rect 34707 23968 35027 24992
rect 34707 23904 34715 23968
rect 34779 23904 34795 23968
rect 34859 23904 34875 23968
rect 34939 23904 34955 23968
rect 35019 23904 35027 23968
rect 34707 22880 35027 23904
rect 34707 22816 34715 22880
rect 34779 22816 34795 22880
rect 34859 22816 34875 22880
rect 34939 22816 34955 22880
rect 35019 22816 35027 22880
rect 34707 21792 35027 22816
rect 34707 21728 34715 21792
rect 34779 21728 34795 21792
rect 34859 21728 34875 21792
rect 34939 21728 34955 21792
rect 35019 21728 35027 21792
rect 34707 20704 35027 21728
rect 34707 20640 34715 20704
rect 34779 20640 34795 20704
rect 34859 20640 34875 20704
rect 34939 20640 34955 20704
rect 35019 20640 35027 20704
rect 34707 19616 35027 20640
rect 34707 19552 34715 19616
rect 34779 19552 34795 19616
rect 34859 19552 34875 19616
rect 34939 19552 34955 19616
rect 35019 19552 35027 19616
rect 34707 18528 35027 19552
rect 34707 18464 34715 18528
rect 34779 18464 34795 18528
rect 34859 18464 34875 18528
rect 34939 18464 34955 18528
rect 35019 18464 35027 18528
rect 34707 17440 35027 18464
rect 34707 17376 34715 17440
rect 34779 17376 34795 17440
rect 34859 17376 34875 17440
rect 34939 17376 34955 17440
rect 35019 17376 35027 17440
rect 34707 16352 35027 17376
rect 34707 16288 34715 16352
rect 34779 16288 34795 16352
rect 34859 16288 34875 16352
rect 34939 16288 34955 16352
rect 35019 16288 35027 16352
rect 34707 15264 35027 16288
rect 34707 15200 34715 15264
rect 34779 15200 34795 15264
rect 34859 15200 34875 15264
rect 34939 15200 34955 15264
rect 35019 15200 35027 15264
rect 34707 14176 35027 15200
rect 34707 14112 34715 14176
rect 34779 14112 34795 14176
rect 34859 14112 34875 14176
rect 34939 14112 34955 14176
rect 35019 14112 35027 14176
rect 34707 13088 35027 14112
rect 34707 13024 34715 13088
rect 34779 13024 34795 13088
rect 34859 13024 34875 13088
rect 34939 13024 34955 13088
rect 35019 13024 35027 13088
rect 34707 12000 35027 13024
rect 34707 11936 34715 12000
rect 34779 11936 34795 12000
rect 34859 11936 34875 12000
rect 34939 11936 34955 12000
rect 35019 11936 35027 12000
rect 34707 10912 35027 11936
rect 34707 10848 34715 10912
rect 34779 10848 34795 10912
rect 34859 10848 34875 10912
rect 34939 10848 34955 10912
rect 35019 10848 35027 10912
rect 34707 9824 35027 10848
rect 34707 9760 34715 9824
rect 34779 9760 34795 9824
rect 34859 9760 34875 9824
rect 34939 9760 34955 9824
rect 35019 9760 35027 9824
rect 34707 8736 35027 9760
rect 34707 8672 34715 8736
rect 34779 8672 34795 8736
rect 34859 8672 34875 8736
rect 34939 8672 34955 8736
rect 35019 8672 35027 8736
rect 34707 7648 35027 8672
rect 34707 7584 34715 7648
rect 34779 7584 34795 7648
rect 34859 7584 34875 7648
rect 34939 7584 34955 7648
rect 35019 7584 35027 7648
rect 34707 6560 35027 7584
rect 34707 6496 34715 6560
rect 34779 6496 34795 6560
rect 34859 6496 34875 6560
rect 34939 6496 34955 6560
rect 35019 6496 35027 6560
rect 34707 5472 35027 6496
rect 34707 5408 34715 5472
rect 34779 5408 34795 5472
rect 34859 5408 34875 5472
rect 34939 5408 34955 5472
rect 35019 5408 35027 5472
rect 34707 4384 35027 5408
rect 34707 4320 34715 4384
rect 34779 4320 34795 4384
rect 34859 4320 34875 4384
rect 34939 4320 34955 4384
rect 35019 4320 35027 4384
rect 34707 3296 35027 4320
rect 34707 3232 34715 3296
rect 34779 3232 34795 3296
rect 34859 3232 34875 3296
rect 34939 3232 34955 3296
rect 35019 3232 35027 3296
rect 34707 2208 35027 3232
rect 34707 2144 34715 2208
rect 34779 2144 34795 2208
rect 34859 2144 34875 2208
rect 34939 2144 34955 2208
rect 35019 2144 35027 2208
rect 34707 2128 35027 2144
use sky130_fd_sc_hd__inv_2  _427_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 20700 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _428_
timestamp 1688980957
transform 1 0 20608 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _429_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 19320 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _430_
timestamp 1688980957
transform -1 0 19136 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _431_
timestamp 1688980957
transform -1 0 17664 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _432_
timestamp 1688980957
transform -1 0 16100 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _433_
timestamp 1688980957
transform 1 0 14352 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _434_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 18032 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _435_
timestamp 1688980957
transform -1 0 14352 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _436_
timestamp 1688980957
transform 1 0 15272 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _437_
timestamp 1688980957
transform -1 0 14076 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _438_
timestamp 1688980957
transform 1 0 14352 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _439_
timestamp 1688980957
transform 1 0 15548 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _440_
timestamp 1688980957
transform 1 0 16652 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _441_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 17020 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _442_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 17940 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _443_
timestamp 1688980957
transform 1 0 18952 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  _444_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 9568 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _445_
timestamp 1688980957
transform -1 0 11960 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _446_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 11592 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _447_
timestamp 1688980957
transform 1 0 14720 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _448_
timestamp 1688980957
transform 1 0 19964 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _449_
timestamp 1688980957
transform -1 0 22448 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _450_
timestamp 1688980957
transform -1 0 20884 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _451_
timestamp 1688980957
transform -1 0 20608 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _452_
timestamp 1688980957
transform -1 0 20608 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _453_
timestamp 1688980957
transform -1 0 19412 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _454_
timestamp 1688980957
transform 1 0 19412 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _455_
timestamp 1688980957
transform -1 0 21160 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _456_
timestamp 1688980957
transform -1 0 20884 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _457_
timestamp 1688980957
transform -1 0 19872 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _458_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 20424 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _459_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 19872 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _460_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 20056 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _461_
timestamp 1688980957
transform -1 0 19964 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _462_
timestamp 1688980957
transform -1 0 20332 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _463_
timestamp 1688980957
transform 1 0 19412 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _464_
timestamp 1688980957
transform -1 0 20424 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _465_
timestamp 1688980957
transform 1 0 19872 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  _466_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 16836 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__a211oi_4  _467_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 21344 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  _468_
timestamp 1688980957
transform -1 0 11316 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _469_
timestamp 1688980957
transform -1 0 10764 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _470_
timestamp 1688980957
transform 1 0 11500 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _471_
timestamp 1688980957
transform -1 0 12696 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _472_
timestamp 1688980957
transform -1 0 13432 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _473_
timestamp 1688980957
transform -1 0 13432 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _474_
timestamp 1688980957
transform -1 0 14168 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _475_
timestamp 1688980957
transform -1 0 14444 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _476_
timestamp 1688980957
transform -1 0 14720 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _477_
timestamp 1688980957
transform 1 0 14720 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _478_
timestamp 1688980957
transform -1 0 15456 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _479_
timestamp 1688980957
transform -1 0 15088 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _480_
timestamp 1688980957
transform -1 0 14812 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _481_
timestamp 1688980957
transform -1 0 13064 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _482_
timestamp 1688980957
transform -1 0 12696 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _483_
timestamp 1688980957
transform -1 0 12236 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _484_
timestamp 1688980957
transform -1 0 11224 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__a211oi_2  _485_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 11316 0 1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__inv_2  _486_
timestamp 1688980957
transform 1 0 7820 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _487_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 17848 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__o41a_1  _488_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 16928 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__and4_1  _489_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 17756 0 1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__a41o_1  _490_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 17204 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  _491_
timestamp 1688980957
transform 1 0 13432 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _492_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 16744 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  _493_
timestamp 1688980957
transform 1 0 13432 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _494_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 14720 0 1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _495_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 14076 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _496_
timestamp 1688980957
transform -1 0 15732 0 1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _497_
timestamp 1688980957
transform -1 0 13984 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _498_
timestamp 1688980957
transform -1 0 15456 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _499_
timestamp 1688980957
transform -1 0 14720 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _500_
timestamp 1688980957
transform -1 0 17112 0 -1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _501_
timestamp 1688980957
transform -1 0 15824 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _502_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 18952 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _503_
timestamp 1688980957
transform -1 0 18308 0 1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _504_
timestamp 1688980957
transform -1 0 17112 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _505_
timestamp 1688980957
transform 1 0 16284 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _506_
timestamp 1688980957
transform -1 0 17664 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _507_
timestamp 1688980957
transform 1 0 17572 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _508_
timestamp 1688980957
transform -1 0 19136 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _509_
timestamp 1688980957
transform -1 0 19872 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _510_
timestamp 1688980957
transform -1 0 15824 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _511_
timestamp 1688980957
transform -1 0 21712 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__o41a_1  _512_
timestamp 1688980957
transform 1 0 21804 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__and4_1  _513_
timestamp 1688980957
transform 1 0 21804 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__a41o_1  _514_
timestamp 1688980957
transform 1 0 21712 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _515_
timestamp 1688980957
transform -1 0 20792 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _516_
timestamp 1688980957
transform 1 0 23460 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _517_
timestamp 1688980957
transform -1 0 24380 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _518_
timestamp 1688980957
transform 1 0 20240 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _519_
timestamp 1688980957
transform 1 0 20700 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _520_
timestamp 1688980957
transform -1 0 23184 0 1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _521_
timestamp 1688980957
transform 1 0 20516 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _522_
timestamp 1688980957
transform -1 0 23644 0 1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _523_
timestamp 1688980957
transform -1 0 21528 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _524_
timestamp 1688980957
transform 1 0 22356 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _525_
timestamp 1688980957
transform -1 0 23092 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _526_
timestamp 1688980957
transform -1 0 21620 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _527_
timestamp 1688980957
transform 1 0 20056 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _528_
timestamp 1688980957
transform 1 0 20700 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _529_
timestamp 1688980957
transform 1 0 21344 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _530_
timestamp 1688980957
transform -1 0 9752 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _531_
timestamp 1688980957
transform 1 0 23368 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _532_
timestamp 1688980957
transform 1 0 23828 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _533_
timestamp 1688980957
transform -1 0 24288 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__o41a_1  _534_
timestamp 1688980957
transform 1 0 22908 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__and4_1  _535_
timestamp 1688980957
transform -1 0 24564 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__a41o_1  _536_
timestamp 1688980957
transform 1 0 23276 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _537_
timestamp 1688980957
transform 1 0 22540 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _538_
timestamp 1688980957
transform 1 0 23736 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _539_
timestamp 1688980957
transform 1 0 23828 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _540_
timestamp 1688980957
transform -1 0 25024 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _541_
timestamp 1688980957
transform -1 0 23920 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _542_
timestamp 1688980957
transform 1 0 23000 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _543_
timestamp 1688980957
transform 1 0 24380 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _544_
timestamp 1688980957
transform 1 0 24104 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _545_
timestamp 1688980957
transform 1 0 24564 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _546_
timestamp 1688980957
transform -1 0 24840 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _547_
timestamp 1688980957
transform 1 0 23920 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _548_
timestamp 1688980957
transform 1 0 21988 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _549_
timestamp 1688980957
transform 1 0 22264 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _550_
timestamp 1688980957
transform 1 0 21804 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _551_
timestamp 1688980957
transform -1 0 22816 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _552_
timestamp 1688980957
transform -1 0 23092 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _553_
timestamp 1688980957
transform -1 0 21436 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _554_
timestamp 1688980957
transform 1 0 10856 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__o41a_1  _555_
timestamp 1688980957
transform -1 0 13708 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__and4_1  _556_
timestamp 1688980957
transform 1 0 11684 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__a41o_1  _557_
timestamp 1688980957
transform -1 0 13248 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _558_
timestamp 1688980957
transform -1 0 13340 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _559_
timestamp 1688980957
transform 1 0 8280 0 1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _560_
timestamp 1688980957
transform -1 0 9108 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _561_
timestamp 1688980957
transform -1 0 11316 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _562_
timestamp 1688980957
transform -1 0 9016 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _563_
timestamp 1688980957
transform -1 0 10672 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _564_
timestamp 1688980957
transform 1 0 9936 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _565_
timestamp 1688980957
transform 1 0 11592 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _566_
timestamp 1688980957
transform -1 0 10856 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _567_
timestamp 1688980957
transform 1 0 10120 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _568_
timestamp 1688980957
transform -1 0 12788 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _569_
timestamp 1688980957
transform 1 0 11500 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _570_
timestamp 1688980957
transform -1 0 12604 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _571_
timestamp 1688980957
transform -1 0 11408 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _572_
timestamp 1688980957
transform 1 0 12052 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _573_
timestamp 1688980957
transform 1 0 14076 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _574_
timestamp 1688980957
transform -1 0 14536 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _575_
timestamp 1688980957
transform 1 0 12880 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _576_
timestamp 1688980957
transform 1 0 9660 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__o41a_1  _577_
timestamp 1688980957
transform 1 0 10488 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__and4_1  _578_
timestamp 1688980957
transform -1 0 8280 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__a41o_1  _579_
timestamp 1688980957
transform 1 0 9752 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _580_
timestamp 1688980957
transform 1 0 9016 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _581_
timestamp 1688980957
transform 1 0 5888 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _582_
timestamp 1688980957
transform -1 0 6808 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _583_
timestamp 1688980957
transform -1 0 8740 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _584_
timestamp 1688980957
transform 1 0 8004 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _585_
timestamp 1688980957
transform -1 0 9936 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _586_
timestamp 1688980957
transform -1 0 7636 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _587_
timestamp 1688980957
transform 1 0 7636 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _588_
timestamp 1688980957
transform 1 0 8280 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _589_
timestamp 1688980957
transform -1 0 9384 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _590_
timestamp 1688980957
transform -1 0 8832 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _591_
timestamp 1688980957
transform 1 0 9752 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _592_
timestamp 1688980957
transform 1 0 11132 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _593_
timestamp 1688980957
transform 1 0 12696 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _594_
timestamp 1688980957
transform 1 0 10948 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _595_
timestamp 1688980957
transform -1 0 11592 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _596_
timestamp 1688980957
transform -1 0 12696 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _597_
timestamp 1688980957
transform -1 0 11592 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _598_
timestamp 1688980957
transform -1 0 8832 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__o41a_1  _599_
timestamp 1688980957
transform -1 0 10948 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__and4_1  _600_
timestamp 1688980957
transform 1 0 9200 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a41o_1  _601_
timestamp 1688980957
transform -1 0 10856 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _602_
timestamp 1688980957
transform -1 0 12236 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _603_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 16376 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _604_
timestamp 1688980957
transform 1 0 12972 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _605_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 16560 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _606_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 13984 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _607_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 15548 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _608_
timestamp 1688980957
transform -1 0 14536 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_1  _609_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14260 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _610_
timestamp 1688980957
transform -1 0 13524 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _611_
timestamp 1688980957
transform -1 0 13800 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _612_
timestamp 1688980957
transform -1 0 13340 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _613_
timestamp 1688980957
transform 1 0 15272 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _614_
timestamp 1688980957
transform -1 0 13984 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _615_
timestamp 1688980957
transform 1 0 13524 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _616_
timestamp 1688980957
transform 1 0 12236 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _617_
timestamp 1688980957
transform -1 0 12696 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _618_
timestamp 1688980957
transform -1 0 9844 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _619_
timestamp 1688980957
transform 1 0 10764 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _620_
timestamp 1688980957
transform -1 0 12052 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _621_
timestamp 1688980957
transform 1 0 9016 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _622_
timestamp 1688980957
transform 1 0 8280 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _623_
timestamp 1688980957
transform 1 0 9844 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _624_
timestamp 1688980957
transform -1 0 9476 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _625_
timestamp 1688980957
transform 1 0 14352 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _626_
timestamp 1688980957
transform 1 0 14996 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _627_
timestamp 1688980957
transform 1 0 5796 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _628_
timestamp 1688980957
transform -1 0 6624 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _629_
timestamp 1688980957
transform -1 0 8464 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _630_
timestamp 1688980957
transform 1 0 7912 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _631_
timestamp 1688980957
transform -1 0 7820 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _632_
timestamp 1688980957
transform -1 0 7268 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _633_
timestamp 1688980957
transform -1 0 8280 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _634_
timestamp 1688980957
transform -1 0 7544 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _635_
timestamp 1688980957
transform 1 0 9016 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _636_
timestamp 1688980957
transform 1 0 9844 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _637_
timestamp 1688980957
transform 1 0 10028 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _638_
timestamp 1688980957
transform 1 0 10488 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _639_
timestamp 1688980957
transform 1 0 9108 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _640_
timestamp 1688980957
transform 1 0 10028 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _641_
timestamp 1688980957
transform -1 0 11960 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _642_
timestamp 1688980957
transform -1 0 10028 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _643_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 16744 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _644_
timestamp 1688980957
transform 1 0 16744 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _645_
timestamp 1688980957
transform 1 0 16008 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _646_
timestamp 1688980957
transform -1 0 16560 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_2  _647_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 16468 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  _648_
timestamp 1688980957
transform -1 0 14536 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _649_
timestamp 1688980957
transform -1 0 14444 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _650_
timestamp 1688980957
transform 1 0 14168 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _651_
timestamp 1688980957
transform -1 0 19136 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _652_
timestamp 1688980957
transform -1 0 14536 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _653_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 15088 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _654_
timestamp 1688980957
transform 1 0 14444 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _655_
timestamp 1688980957
transform -1 0 13984 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _656_
timestamp 1688980957
transform 1 0 13156 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _657_
timestamp 1688980957
transform 1 0 13340 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__a21boi_2  _658_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14076 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _659_
timestamp 1688980957
transform 1 0 15732 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _660_
timestamp 1688980957
transform 1 0 16192 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _661_
timestamp 1688980957
transform -1 0 17204 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _662_
timestamp 1688980957
transform 1 0 15916 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _663_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 15548 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _664_
timestamp 1688980957
transform -1 0 14812 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _665_
timestamp 1688980957
transform -1 0 15548 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _666_
timestamp 1688980957
transform -1 0 16376 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _667_
timestamp 1688980957
transform 1 0 15548 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _668_
timestamp 1688980957
transform -1 0 15732 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _669_
timestamp 1688980957
transform -1 0 17204 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _670_
timestamp 1688980957
transform 1 0 14812 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _671_
timestamp 1688980957
transform 1 0 17204 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_1  _672_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 15732 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _673_
timestamp 1688980957
transform -1 0 17572 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _674_
timestamp 1688980957
transform -1 0 19688 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _675_
timestamp 1688980957
transform -1 0 16928 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _676_
timestamp 1688980957
transform -1 0 18124 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _677_
timestamp 1688980957
transform 1 0 17664 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _678_
timestamp 1688980957
transform -1 0 18952 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _679_
timestamp 1688980957
transform 1 0 18492 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _680_
timestamp 1688980957
transform -1 0 17756 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _681_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 18308 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _682_
timestamp 1688980957
transform 1 0 17572 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _683_
timestamp 1688980957
transform -1 0 20976 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _684_
timestamp 1688980957
transform 1 0 21160 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _685_
timestamp 1688980957
transform 1 0 19688 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _686_
timestamp 1688980957
transform 1 0 20700 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _687_
timestamp 1688980957
transform 1 0 18952 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_1  _688_
timestamp 1688980957
transform -1 0 18216 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _689_
timestamp 1688980957
transform 1 0 20424 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _690_
timestamp 1688980957
transform 1 0 19688 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__o22ai_1  _691_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 19688 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _692_
timestamp 1688980957
transform -1 0 20976 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _693_
timestamp 1688980957
transform -1 0 19228 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _694_
timestamp 1688980957
transform -1 0 20516 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _695_
timestamp 1688980957
transform 1 0 20148 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__o31ai_1  _696_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 19872 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _697_
timestamp 1688980957
transform 1 0 19504 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _698_
timestamp 1688980957
transform -1 0 23828 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _699_
timestamp 1688980957
transform -1 0 22080 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _700_
timestamp 1688980957
transform 1 0 15824 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _701_
timestamp 1688980957
transform 1 0 16008 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _702_
timestamp 1688980957
transform 1 0 22080 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _703_
timestamp 1688980957
transform 1 0 21344 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _704_
timestamp 1688980957
transform -1 0 23736 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _705_
timestamp 1688980957
transform 1 0 24196 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_2  _706_
timestamp 1688980957
transform 1 0 22172 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _707_
timestamp 1688980957
transform 1 0 21804 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _708_
timestamp 1688980957
transform 1 0 20332 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _709_
timestamp 1688980957
transform 1 0 21068 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _710_
timestamp 1688980957
transform -1 0 23552 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _711_
timestamp 1688980957
transform -1 0 22264 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _712_
timestamp 1688980957
transform 1 0 20700 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _713_
timestamp 1688980957
transform -1 0 21712 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _714_
timestamp 1688980957
transform -1 0 21528 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _715_
timestamp 1688980957
transform 1 0 20424 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _716_
timestamp 1688980957
transform 1 0 20976 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__a21boi_2  _717_
timestamp 1688980957
transform 1 0 20792 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _718_
timestamp 1688980957
transform 1 0 22172 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _719_
timestamp 1688980957
transform -1 0 22172 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _720_
timestamp 1688980957
transform 1 0 23000 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _721_
timestamp 1688980957
transform -1 0 23552 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _722_
timestamp 1688980957
transform 1 0 21804 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _723_
timestamp 1688980957
transform -1 0 23184 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _724_
timestamp 1688980957
transform -1 0 23184 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _725_
timestamp 1688980957
transform 1 0 21804 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _726_
timestamp 1688980957
transform 1 0 22632 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _727_
timestamp 1688980957
transform -1 0 24288 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _728_
timestamp 1688980957
transform 1 0 22632 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _729_
timestamp 1688980957
transform -1 0 23368 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _730_
timestamp 1688980957
transform -1 0 21712 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_1  _731_
timestamp 1688980957
transform -1 0 22632 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _732_
timestamp 1688980957
transform -1 0 21712 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _733_
timestamp 1688980957
transform 1 0 21160 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _734_
timestamp 1688980957
transform 1 0 23644 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _735_
timestamp 1688980957
transform 1 0 22172 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _736_
timestamp 1688980957
transform 1 0 24288 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _737_
timestamp 1688980957
transform 1 0 22632 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _738_
timestamp 1688980957
transform -1 0 23092 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _739_
timestamp 1688980957
transform 1 0 20700 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _740_
timestamp 1688980957
transform -1 0 22356 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__o31ai_1  _741_
timestamp 1688980957
transform -1 0 22816 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _742_
timestamp 1688980957
transform 1 0 21988 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _743_
timestamp 1688980957
transform -1 0 20608 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _744_
timestamp 1688980957
transform 1 0 21252 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _745_
timestamp 1688980957
transform 1 0 22264 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _746_
timestamp 1688980957
transform -1 0 23644 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_1  _747_
timestamp 1688980957
transform 1 0 21620 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _748_
timestamp 1688980957
transform 1 0 22448 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _749_
timestamp 1688980957
transform -1 0 21620 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _750_
timestamp 1688980957
transform -1 0 21344 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _751_
timestamp 1688980957
transform -1 0 20332 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _752_
timestamp 1688980957
transform 1 0 21804 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _753_
timestamp 1688980957
transform 1 0 21712 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__o31ai_1  _754_
timestamp 1688980957
transform 1 0 23184 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _755_
timestamp 1688980957
transform 1 0 21528 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _756_
timestamp 1688980957
transform 1 0 12236 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _757_
timestamp 1688980957
transform 1 0 14076 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _758_
timestamp 1688980957
transform 1 0 20884 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _759_
timestamp 1688980957
transform -1 0 21344 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _760_
timestamp 1688980957
transform 1 0 12236 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _761_
timestamp 1688980957
transform 1 0 12144 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _762_
timestamp 1688980957
transform -1 0 13340 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _763_
timestamp 1688980957
transform -1 0 13616 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_2  _764_
timestamp 1688980957
transform -1 0 13984 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _765_
timestamp 1688980957
transform 1 0 14260 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _766_
timestamp 1688980957
transform -1 0 14996 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _767_
timestamp 1688980957
transform -1 0 14904 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _768_
timestamp 1688980957
transform -1 0 13340 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _769_
timestamp 1688980957
transform 1 0 15088 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _770_
timestamp 1688980957
transform 1 0 14996 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _771_
timestamp 1688980957
transform 1 0 14536 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _772_
timestamp 1688980957
transform 1 0 15272 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _773_
timestamp 1688980957
transform 1 0 15548 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _774_
timestamp 1688980957
transform -1 0 16468 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__a21boi_2  _775_
timestamp 1688980957
transform 1 0 14904 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _776_
timestamp 1688980957
transform 1 0 14260 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _777_
timestamp 1688980957
transform 1 0 13432 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _778_
timestamp 1688980957
transform 1 0 14076 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _779_
timestamp 1688980957
transform -1 0 14996 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _780_
timestamp 1688980957
transform 1 0 14076 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _781_
timestamp 1688980957
transform 1 0 15456 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _782_
timestamp 1688980957
transform -1 0 15456 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _783_
timestamp 1688980957
transform 1 0 12788 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _784_
timestamp 1688980957
transform 1 0 13616 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _785_
timestamp 1688980957
transform -1 0 14628 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _786_
timestamp 1688980957
transform 1 0 14076 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _787_
timestamp 1688980957
transform 1 0 12788 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _788_
timestamp 1688980957
transform 1 0 13616 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_1  _789_
timestamp 1688980957
transform 1 0 13432 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _790_
timestamp 1688980957
transform 1 0 13340 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _791_
timestamp 1688980957
transform -1 0 13340 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _792_
timestamp 1688980957
transform 1 0 12144 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _793_
timestamp 1688980957
transform 1 0 12236 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _794_
timestamp 1688980957
transform -1 0 12420 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _795_
timestamp 1688980957
transform 1 0 13432 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _796_
timestamp 1688980957
transform 1 0 12696 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _797_
timestamp 1688980957
transform 1 0 10580 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _798_
timestamp 1688980957
transform 1 0 12052 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__o31ai_1  _799_
timestamp 1688980957
transform -1 0 12052 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _800_
timestamp 1688980957
transform -1 0 12052 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _801_
timestamp 1688980957
transform -1 0 10028 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _802_
timestamp 1688980957
transform -1 0 12604 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _803_
timestamp 1688980957
transform -1 0 12236 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _804_
timestamp 1688980957
transform 1 0 12696 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_1  _805_
timestamp 1688980957
transform 1 0 12236 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _806_
timestamp 1688980957
transform -1 0 10580 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _807_
timestamp 1688980957
transform -1 0 11408 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _808_
timestamp 1688980957
transform 1 0 10028 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _809_
timestamp 1688980957
transform 1 0 9660 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _810_
timestamp 1688980957
transform 1 0 10028 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _811_
timestamp 1688980957
transform 1 0 11224 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__o31ai_1  _812_
timestamp 1688980957
transform -1 0 12144 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _813_
timestamp 1688980957
transform 1 0 11500 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _814_
timestamp 1688980957
transform 1 0 10948 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _815_
timestamp 1688980957
transform -1 0 11776 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _816_
timestamp 1688980957
transform -1 0 13984 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _817_
timestamp 1688980957
transform -1 0 16100 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _818_
timestamp 1688980957
transform 1 0 13524 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _819_
timestamp 1688980957
transform 1 0 14628 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _820_
timestamp 1688980957
transform -1 0 16008 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_1  _821_
timestamp 1688980957
transform 1 0 16192 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _822_
timestamp 1688980957
transform 1 0 16100 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _823_
timestamp 1688980957
transform 1 0 17664 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _824_
timestamp 1688980957
transform -1 0 17020 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _825_
timestamp 1688980957
transform 1 0 17204 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _826_
timestamp 1688980957
transform -1 0 16008 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _827_
timestamp 1688980957
transform 1 0 16652 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _828_
timestamp 1688980957
transform -1 0 19596 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _829_
timestamp 1688980957
transform -1 0 18768 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _830_
timestamp 1688980957
transform -1 0 18584 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _831_
timestamp 1688980957
transform -1 0 19688 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _832_
timestamp 1688980957
transform -1 0 18952 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _833_
timestamp 1688980957
transform 1 0 18584 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _834_
timestamp 1688980957
transform -1 0 20332 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _835_
timestamp 1688980957
transform 1 0 20148 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _836_
timestamp 1688980957
transform -1 0 15456 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _837_
timestamp 1688980957
transform -1 0 15824 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _838_
timestamp 1688980957
transform 1 0 15456 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _839_
timestamp 1688980957
transform -1 0 19044 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _840_
timestamp 1688980957
transform -1 0 17112 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_1  _841_
timestamp 1688980957
transform 1 0 17112 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _842_
timestamp 1688980957
transform -1 0 18676 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _843_
timestamp 1688980957
transform -1 0 19044 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _844_
timestamp 1688980957
transform -1 0 18216 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _845_
timestamp 1688980957
transform 1 0 19228 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _846_
timestamp 1688980957
transform 1 0 17664 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _847_
timestamp 1688980957
transform 1 0 16744 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _848_
timestamp 1688980957
transform -1 0 19596 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _849_
timestamp 1688980957
transform 1 0 17848 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _850_
timestamp 1688980957
transform 1 0 15548 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _851_
timestamp 1688980957
transform -1 0 19688 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _852_
timestamp 1688980957
transform -1 0 19136 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _853_
timestamp 1688980957
transform 1 0 17388 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _854_
timestamp 1688980957
transform 1 0 18676 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _855_
timestamp 1688980957
transform 1 0 18400 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _856__12 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 7636 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__dfstp_1  _856_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 6900 0 1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__dfxtp_1  _857_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 16652 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _858_
timestamp 1688980957
transform 1 0 14076 0 -1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _859_
timestamp 1688980957
transform 1 0 14168 0 1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _860_
timestamp 1688980957
transform 1 0 14720 0 -1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _861_
timestamp 1688980957
transform 1 0 15824 0 1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _862_
timestamp 1688980957
transform 1 0 17112 0 -1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _863_
timestamp 1688980957
transform 1 0 17664 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _864_
timestamp 1688980957
transform -1 0 20700 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _865_
timestamp 1688980957
transform -1 0 19412 0 -1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _866_
timestamp 1688980957
transform -1 0 21712 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _867_
timestamp 1688980957
transform -1 0 24840 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _868_
timestamp 1688980957
transform 1 0 19596 0 1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _869_
timestamp 1688980957
transform 1 0 20148 0 -1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _870_
timestamp 1688980957
transform -1 0 23276 0 -1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _871_
timestamp 1688980957
transform -1 0 23368 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _872_
timestamp 1688980957
transform 1 0 19136 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _873_
timestamp 1688980957
transform 1 0 20792 0 1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _874_
timestamp 1688980957
transform -1 0 23828 0 1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _875_
timestamp 1688980957
transform -1 0 22908 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _876_
timestamp 1688980957
transform 1 0 23276 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _877_
timestamp 1688980957
transform 1 0 24380 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _878_
timestamp 1688980957
transform 1 0 24012 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _879_
timestamp 1688980957
transform -1 0 24840 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _880_
timestamp 1688980957
transform -1 0 24104 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _881_
timestamp 1688980957
transform -1 0 22448 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _882_
timestamp 1688980957
transform 1 0 22448 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _883_
timestamp 1688980957
transform 1 0 21804 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _884_
timestamp 1688980957
transform 1 0 14076 0 1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _885_
timestamp 1688980957
transform 1 0 8740 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _886_
timestamp 1688980957
transform 1 0 9568 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _887_
timestamp 1688980957
transform 1 0 9384 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _888_
timestamp 1688980957
transform 1 0 9568 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _889_
timestamp 1688980957
transform 1 0 11040 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _890_
timestamp 1688980957
transform 1 0 11960 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _891_
timestamp 1688980957
transform -1 0 13984 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _892_
timestamp 1688980957
transform 1 0 12512 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _893_
timestamp 1688980957
transform 1 0 10856 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _894_
timestamp 1688980957
transform 1 0 6808 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _895_
timestamp 1688980957
transform 1 0 7360 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _896_
timestamp 1688980957
transform 1 0 8924 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _897_
timestamp 1688980957
transform 1 0 7360 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _898_
timestamp 1688980957
transform 1 0 8924 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _899_
timestamp 1688980957
transform -1 0 11132 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _900_
timestamp 1688980957
transform -1 0 12972 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _901_
timestamp 1688980957
transform -1 0 12972 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _902_
timestamp 1688980957
transform -1 0 12236 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _903_
timestamp 1688980957
transform -1 0 16560 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _904_
timestamp 1688980957
transform -1 0 17112 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _905_
timestamp 1688980957
transform 1 0 14168 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _906_
timestamp 1688980957
transform 1 0 12788 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _907_
timestamp 1688980957
transform -1 0 13064 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _908_
timestamp 1688980957
transform 1 0 10120 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _909_
timestamp 1688980957
transform 1 0 9292 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _910_
timestamp 1688980957
transform 1 0 8924 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _911_
timestamp 1688980957
transform 1 0 14536 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _912_
timestamp 1688980957
transform 1 0 6532 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _913_
timestamp 1688980957
transform 1 0 7360 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _914_
timestamp 1688980957
transform 1 0 7360 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _915_
timestamp 1688980957
transform 1 0 7544 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _916_
timestamp 1688980957
transform 1 0 9200 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _917_
timestamp 1688980957
transform 1 0 8924 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _918_
timestamp 1688980957
transform 1 0 9568 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _919_
timestamp 1688980957
transform 1 0 9844 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _920_
timestamp 1688980957
transform 1 0 12696 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _921_
timestamp 1688980957
transform 1 0 12512 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _922_
timestamp 1688980957
transform 1 0 14720 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _923_
timestamp 1688980957
transform 1 0 15824 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _924_
timestamp 1688980957
transform -1 0 19044 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _925_
timestamp 1688980957
transform -1 0 19136 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _926_
timestamp 1688980957
transform 1 0 19228 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _927_
timestamp 1688980957
transform -1 0 21344 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _928_
timestamp 1688980957
transform 1 0 21896 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _929_
timestamp 1688980957
transform 1 0 14812 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _930_
timestamp 1688980957
transform 1 0 19964 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _931_
timestamp 1688980957
transform -1 0 21344 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _932_
timestamp 1688980957
transform 1 0 23184 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _933_
timestamp 1688980957
transform 1 0 22816 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _934_
timestamp 1688980957
transform 1 0 23092 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _935_
timestamp 1688980957
transform 1 0 22816 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _936_
timestamp 1688980957
transform 1 0 19412 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _937_
timestamp 1688980957
transform 1 0 22356 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _938_
timestamp 1688980957
transform 1 0 11868 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _939_
timestamp 1688980957
transform 1 0 21804 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _940_
timestamp 1688980957
transform 1 0 14720 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _941_
timestamp 1688980957
transform -1 0 17388 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _942_
timestamp 1688980957
transform -1 0 16192 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _943_
timestamp 1688980957
transform 1 0 12512 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _944_
timestamp 1688980957
transform -1 0 14168 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _945_
timestamp 1688980957
transform 1 0 9752 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _946_
timestamp 1688980957
transform 1 0 8924 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _947_
timestamp 1688980957
transform -1 0 12512 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _948_
timestamp 1688980957
transform 1 0 11776 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _949_
timestamp 1688980957
transform 1 0 13892 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _950_
timestamp 1688980957
transform 1 0 14076 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _951_
timestamp 1688980957
transform -1 0 15732 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _952_
timestamp 1688980957
transform -1 0 17480 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _953_
timestamp 1688980957
transform 1 0 16652 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _954_
timestamp 1688980957
transform 1 0 17664 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _955_
timestamp 1688980957
transform 1 0 18308 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _956_
timestamp 1688980957
transform 1 0 19596 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _957_
timestamp 1688980957
transform 1 0 16192 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _958_
timestamp 1688980957
transform 1 0 16652 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _959_
timestamp 1688980957
transform 1 0 17664 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _960_
timestamp 1688980957
transform 1 0 18216 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _961_
timestamp 1688980957
transform 1 0 16744 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _962_
timestamp 1688980957
transform 1 0 16928 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _963_
timestamp 1688980957
transform 1 0 17664 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _964_
timestamp 1688980957
transform 1 0 17664 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  _976_
timestamp 1688980957
transform 1 0 7452 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 18032 0 1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_0__f_clk
timestamp 1688980957
transform 1 0 10396 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_1__f_clk
timestamp 1688980957
transform -1 0 9660 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_2__f_clk
timestamp 1688980957
transform -1 0 20056 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_3__f_clk
timestamp 1688980957
transform 1 0 18216 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_4__f_clk
timestamp 1688980957
transform 1 0 10396 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_5__f_clk
timestamp 1688980957
transform 1 0 10396 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_6__f_clk
timestamp 1688980957
transform 1 0 20792 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_7__f_clk
timestamp 1688980957
transform -1 0 20056 0 -1 36992
box -38 -48 1878 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_6 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1656 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_18 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2760 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_26 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3496 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_29
timestamp 1688980957
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_41
timestamp 1688980957
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_53 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_57
timestamp 1688980957
transform 1 0 6348 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_62
timestamp 1688980957
transform 1 0 6808 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_74
timestamp 1688980957
transform 1 0 7912 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_82
timestamp 1688980957
transform 1 0 8648 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_85
timestamp 1688980957
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_97
timestamp 1688980957
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_109
timestamp 1688980957
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_113
timestamp 1688980957
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_125
timestamp 1688980957
transform 1 0 12604 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_133
timestamp 1688980957
transform 1 0 13340 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_139 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 13892 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_141
timestamp 1688980957
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_153
timestamp 1688980957
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_165
timestamp 1688980957
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_169
timestamp 1688980957
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_181
timestamp 1688980957
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_193
timestamp 1688980957
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_197
timestamp 1688980957
transform 1 0 19228 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_205
timestamp 1688980957
transform 1 0 19964 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_225
timestamp 1688980957
transform 1 0 21804 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_237
timestamp 1688980957
transform 1 0 22908 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_249
timestamp 1688980957
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_253
timestamp 1688980957
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_265
timestamp 1688980957
transform 1 0 25484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_277
timestamp 1688980957
transform 1 0 26588 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_281
timestamp 1688980957
transform 1 0 26956 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_286
timestamp 1688980957
transform 1 0 27416 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_298
timestamp 1688980957
transform 1 0 28520 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_306
timestamp 1688980957
transform 1 0 29256 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_309
timestamp 1688980957
transform 1 0 29532 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_321
timestamp 1688980957
transform 1 0 30636 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_333
timestamp 1688980957
transform 1 0 31740 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_337
timestamp 1688980957
transform 1 0 32108 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_349
timestamp 1688980957
transform 1 0 33212 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_357
timestamp 1688980957
transform 1 0 33948 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_363
timestamp 1688980957
transform 1 0 34500 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 1688980957
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 1688980957
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp 1688980957
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_39
timestamp 1688980957
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_51 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 1688980957
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_57
timestamp 1688980957
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_69
timestamp 1688980957
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_81
timestamp 1688980957
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_93
timestamp 1688980957
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_105 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_111
timestamp 1688980957
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_113
timestamp 1688980957
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_125
timestamp 1688980957
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_137
timestamp 1688980957
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_149
timestamp 1688980957
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_161
timestamp 1688980957
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_167
timestamp 1688980957
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_169
timestamp 1688980957
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_181
timestamp 1688980957
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_193
timestamp 1688980957
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_205
timestamp 1688980957
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_217
timestamp 1688980957
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_223
timestamp 1688980957
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_225
timestamp 1688980957
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_237
timestamp 1688980957
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_249
timestamp 1688980957
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_261
timestamp 1688980957
transform 1 0 25116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_273
timestamp 1688980957
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_279
timestamp 1688980957
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_281
timestamp 1688980957
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_293
timestamp 1688980957
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_305
timestamp 1688980957
transform 1 0 29164 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_317
timestamp 1688980957
transform 1 0 30268 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_329
timestamp 1688980957
transform 1 0 31372 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_335
timestamp 1688980957
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_337
timestamp 1688980957
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_349
timestamp 1688980957
transform 1 0 33212 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_361
timestamp 1688980957
transform 1 0 34316 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1688980957
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1688980957
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1688980957
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 1688980957
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 1688980957
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_53
timestamp 1688980957
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_65
timestamp 1688980957
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_77
timestamp 1688980957
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 1688980957
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_85
timestamp 1688980957
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_97
timestamp 1688980957
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_109
timestamp 1688980957
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_121
timestamp 1688980957
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_133
timestamp 1688980957
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_139
timestamp 1688980957
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_141
timestamp 1688980957
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_153
timestamp 1688980957
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_165
timestamp 1688980957
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_177
timestamp 1688980957
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_189
timestamp 1688980957
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_195
timestamp 1688980957
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_197
timestamp 1688980957
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_209
timestamp 1688980957
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_221
timestamp 1688980957
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_233
timestamp 1688980957
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_245
timestamp 1688980957
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_251
timestamp 1688980957
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_253
timestamp 1688980957
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_265
timestamp 1688980957
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_277
timestamp 1688980957
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_289
timestamp 1688980957
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_301
timestamp 1688980957
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_307
timestamp 1688980957
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_309
timestamp 1688980957
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_321
timestamp 1688980957
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_333
timestamp 1688980957
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_345
timestamp 1688980957
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_357
timestamp 1688980957
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_363
timestamp 1688980957
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1688980957
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1688980957
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 1688980957
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 1688980957
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 1688980957
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1688980957
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 1688980957
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_69
timestamp 1688980957
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_81
timestamp 1688980957
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_93
timestamp 1688980957
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_105
timestamp 1688980957
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_111
timestamp 1688980957
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_113
timestamp 1688980957
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_125
timestamp 1688980957
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_137
timestamp 1688980957
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_149
timestamp 1688980957
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_161
timestamp 1688980957
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_167
timestamp 1688980957
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_169
timestamp 1688980957
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_181
timestamp 1688980957
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_193
timestamp 1688980957
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_205
timestamp 1688980957
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_217
timestamp 1688980957
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_223
timestamp 1688980957
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_225
timestamp 1688980957
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_237
timestamp 1688980957
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_249
timestamp 1688980957
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_261
timestamp 1688980957
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_273
timestamp 1688980957
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_279
timestamp 1688980957
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_281
timestamp 1688980957
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_293
timestamp 1688980957
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_305
timestamp 1688980957
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_317
timestamp 1688980957
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_329
timestamp 1688980957
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_335
timestamp 1688980957
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_337
timestamp 1688980957
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_349
timestamp 1688980957
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_361
timestamp 1688980957
transform 1 0 34316 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1688980957
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 1688980957
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1688980957
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1688980957
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 1688980957
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_53
timestamp 1688980957
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_65
timestamp 1688980957
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_77
timestamp 1688980957
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 1688980957
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_85
timestamp 1688980957
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_97
timestamp 1688980957
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_109
timestamp 1688980957
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_121
timestamp 1688980957
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_133
timestamp 1688980957
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_139
timestamp 1688980957
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_141
timestamp 1688980957
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_153
timestamp 1688980957
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_165
timestamp 1688980957
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_177
timestamp 1688980957
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_189
timestamp 1688980957
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_195
timestamp 1688980957
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_197
timestamp 1688980957
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_209
timestamp 1688980957
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_221
timestamp 1688980957
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_233
timestamp 1688980957
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_245
timestamp 1688980957
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_251
timestamp 1688980957
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_253
timestamp 1688980957
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_265
timestamp 1688980957
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_277
timestamp 1688980957
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_289
timestamp 1688980957
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_301
timestamp 1688980957
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_307
timestamp 1688980957
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_309
timestamp 1688980957
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_321
timestamp 1688980957
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_333
timestamp 1688980957
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_345
timestamp 1688980957
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_357
timestamp 1688980957
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_363
timestamp 1688980957
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 1688980957
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 1688980957
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_27
timestamp 1688980957
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_39
timestamp 1688980957
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_51
timestamp 1688980957
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 1688980957
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 1688980957
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_69
timestamp 1688980957
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_81
timestamp 1688980957
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_93
timestamp 1688980957
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_105
timestamp 1688980957
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_111
timestamp 1688980957
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_113
timestamp 1688980957
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_125
timestamp 1688980957
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_137
timestamp 1688980957
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_149
timestamp 1688980957
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_161
timestamp 1688980957
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_167
timestamp 1688980957
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_169
timestamp 1688980957
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_181
timestamp 1688980957
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_193
timestamp 1688980957
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_205
timestamp 1688980957
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_217
timestamp 1688980957
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_223
timestamp 1688980957
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_225
timestamp 1688980957
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_237
timestamp 1688980957
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_249
timestamp 1688980957
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_261
timestamp 1688980957
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_273
timestamp 1688980957
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_279
timestamp 1688980957
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_281
timestamp 1688980957
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_293
timestamp 1688980957
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_305
timestamp 1688980957
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_317
timestamp 1688980957
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_329
timestamp 1688980957
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_335
timestamp 1688980957
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_337
timestamp 1688980957
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_349
timestamp 1688980957
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_361
timestamp 1688980957
transform 1 0 34316 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 1688980957
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp 1688980957
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1688980957
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 1688980957
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_41
timestamp 1688980957
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_53
timestamp 1688980957
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_65
timestamp 1688980957
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_77
timestamp 1688980957
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp 1688980957
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_85
timestamp 1688980957
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_97
timestamp 1688980957
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_109
timestamp 1688980957
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_121
timestamp 1688980957
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_133
timestamp 1688980957
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_139
timestamp 1688980957
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_141
timestamp 1688980957
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_153
timestamp 1688980957
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_165
timestamp 1688980957
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_177
timestamp 1688980957
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_189
timestamp 1688980957
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_195
timestamp 1688980957
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_197
timestamp 1688980957
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_209
timestamp 1688980957
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_221
timestamp 1688980957
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_233
timestamp 1688980957
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_245
timestamp 1688980957
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_251
timestamp 1688980957
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_253
timestamp 1688980957
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_265
timestamp 1688980957
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_277
timestamp 1688980957
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_289
timestamp 1688980957
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_301
timestamp 1688980957
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_307
timestamp 1688980957
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_309
timestamp 1688980957
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_321
timestamp 1688980957
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_333
timestamp 1688980957
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_345
timestamp 1688980957
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_357
timestamp 1688980957
transform 1 0 33948 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 1688980957
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 1688980957
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_27
timestamp 1688980957
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_39
timestamp 1688980957
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_51
timestamp 1688980957
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 1688980957
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_57
timestamp 1688980957
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_69
timestamp 1688980957
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_81
timestamp 1688980957
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_93
timestamp 1688980957
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_105
timestamp 1688980957
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_111
timestamp 1688980957
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_113
timestamp 1688980957
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_125
timestamp 1688980957
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_137
timestamp 1688980957
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_149
timestamp 1688980957
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_161
timestamp 1688980957
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_167
timestamp 1688980957
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_169
timestamp 1688980957
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_181
timestamp 1688980957
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_193
timestamp 1688980957
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_205
timestamp 1688980957
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_217
timestamp 1688980957
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_223
timestamp 1688980957
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_225
timestamp 1688980957
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_237
timestamp 1688980957
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_249
timestamp 1688980957
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_261
timestamp 1688980957
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_273
timestamp 1688980957
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_279
timestamp 1688980957
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_281
timestamp 1688980957
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_293
timestamp 1688980957
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_305
timestamp 1688980957
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_317
timestamp 1688980957
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_329
timestamp 1688980957
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_335
timestamp 1688980957
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_337
timestamp 1688980957
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_349
timestamp 1688980957
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_361
timestamp 1688980957
transform 1 0 34316 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1688980957
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 1688980957
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1688980957
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 1688980957
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_41
timestamp 1688980957
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_53
timestamp 1688980957
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_65
timestamp 1688980957
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_77
timestamp 1688980957
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_83
timestamp 1688980957
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_85
timestamp 1688980957
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_97
timestamp 1688980957
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_109
timestamp 1688980957
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_121
timestamp 1688980957
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_133
timestamp 1688980957
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_139
timestamp 1688980957
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_141
timestamp 1688980957
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_153
timestamp 1688980957
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_165
timestamp 1688980957
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_177
timestamp 1688980957
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_189
timestamp 1688980957
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_195
timestamp 1688980957
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_197
timestamp 1688980957
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_209
timestamp 1688980957
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_221
timestamp 1688980957
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_233
timestamp 1688980957
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_245
timestamp 1688980957
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_251
timestamp 1688980957
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_253
timestamp 1688980957
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_265
timestamp 1688980957
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_277
timestamp 1688980957
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_289
timestamp 1688980957
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_301
timestamp 1688980957
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_307
timestamp 1688980957
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_309
timestamp 1688980957
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_321
timestamp 1688980957
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_333
timestamp 1688980957
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_345
timestamp 1688980957
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_357
timestamp 1688980957
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_363
timestamp 1688980957
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_6
timestamp 1688980957
transform 1 0 1656 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_18
timestamp 1688980957
transform 1 0 2760 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_30
timestamp 1688980957
transform 1 0 3864 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_42
timestamp 1688980957
transform 1 0 4968 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_54
timestamp 1688980957
transform 1 0 6072 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_57
timestamp 1688980957
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_69
timestamp 1688980957
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_81
timestamp 1688980957
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_93
timestamp 1688980957
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_105
timestamp 1688980957
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_111
timestamp 1688980957
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_113
timestamp 1688980957
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_125
timestamp 1688980957
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_137
timestamp 1688980957
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_149
timestamp 1688980957
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_161
timestamp 1688980957
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_167
timestamp 1688980957
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_169
timestamp 1688980957
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_181
timestamp 1688980957
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_193
timestamp 1688980957
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_205
timestamp 1688980957
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_217
timestamp 1688980957
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_223
timestamp 1688980957
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_225
timestamp 1688980957
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_237
timestamp 1688980957
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_249
timestamp 1688980957
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_261
timestamp 1688980957
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_273
timestamp 1688980957
transform 1 0 26220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_279
timestamp 1688980957
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_281
timestamp 1688980957
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_293
timestamp 1688980957
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_305
timestamp 1688980957
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_317
timestamp 1688980957
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_329
timestamp 1688980957
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_335
timestamp 1688980957
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_337
timestamp 1688980957
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_349
timestamp 1688980957
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_361
timestamp 1688980957
transform 1 0 34316 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp 1688980957
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_15
timestamp 1688980957
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 1688980957
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_29
timestamp 1688980957
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_41
timestamp 1688980957
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_53
timestamp 1688980957
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_65
timestamp 1688980957
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_77
timestamp 1688980957
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_83
timestamp 1688980957
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_85
timestamp 1688980957
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_97
timestamp 1688980957
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_109
timestamp 1688980957
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_121
timestamp 1688980957
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_133
timestamp 1688980957
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_139
timestamp 1688980957
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_141
timestamp 1688980957
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_153
timestamp 1688980957
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_165
timestamp 1688980957
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_177
timestamp 1688980957
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_189
timestamp 1688980957
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_195
timestamp 1688980957
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_197
timestamp 1688980957
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_209
timestamp 1688980957
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_221
timestamp 1688980957
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_233
timestamp 1688980957
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_245
timestamp 1688980957
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_251
timestamp 1688980957
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_253
timestamp 1688980957
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_265
timestamp 1688980957
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_277
timestamp 1688980957
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_289
timestamp 1688980957
transform 1 0 27692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_301
timestamp 1688980957
transform 1 0 28796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_307
timestamp 1688980957
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_309
timestamp 1688980957
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_321
timestamp 1688980957
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_333
timestamp 1688980957
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_345
timestamp 1688980957
transform 1 0 32844 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_357
timestamp 1688980957
transform 1 0 33948 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_363
timestamp 1688980957
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_3
timestamp 1688980957
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_15
timestamp 1688980957
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_27
timestamp 1688980957
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_39
timestamp 1688980957
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_51
timestamp 1688980957
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_55
timestamp 1688980957
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_57
timestamp 1688980957
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_69
timestamp 1688980957
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_81
timestamp 1688980957
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_93
timestamp 1688980957
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_105
timestamp 1688980957
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_111
timestamp 1688980957
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_113
timestamp 1688980957
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_125
timestamp 1688980957
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_137
timestamp 1688980957
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_149
timestamp 1688980957
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_161
timestamp 1688980957
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_167
timestamp 1688980957
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_169
timestamp 1688980957
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_181
timestamp 1688980957
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_193
timestamp 1688980957
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_205
timestamp 1688980957
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_217
timestamp 1688980957
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_223
timestamp 1688980957
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_225
timestamp 1688980957
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_237
timestamp 1688980957
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_249
timestamp 1688980957
transform 1 0 24012 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_261
timestamp 1688980957
transform 1 0 25116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_273
timestamp 1688980957
transform 1 0 26220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_279
timestamp 1688980957
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_281
timestamp 1688980957
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_293
timestamp 1688980957
transform 1 0 28060 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_305
timestamp 1688980957
transform 1 0 29164 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_317
timestamp 1688980957
transform 1 0 30268 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_329
timestamp 1688980957
transform 1 0 31372 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_335
timestamp 1688980957
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_337
timestamp 1688980957
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_349
timestamp 1688980957
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_361
timestamp 1688980957
transform 1 0 34316 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_3
timestamp 1688980957
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_15
timestamp 1688980957
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 1688980957
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_29
timestamp 1688980957
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_41
timestamp 1688980957
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_53
timestamp 1688980957
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_65
timestamp 1688980957
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_77
timestamp 1688980957
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_83
timestamp 1688980957
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_85
timestamp 1688980957
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_97
timestamp 1688980957
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_109
timestamp 1688980957
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_121
timestamp 1688980957
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_133
timestamp 1688980957
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_139
timestamp 1688980957
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_141
timestamp 1688980957
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_153
timestamp 1688980957
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_165
timestamp 1688980957
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_177
timestamp 1688980957
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_189
timestamp 1688980957
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_195
timestamp 1688980957
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_197
timestamp 1688980957
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_209
timestamp 1688980957
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_221
timestamp 1688980957
transform 1 0 21436 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_233
timestamp 1688980957
transform 1 0 22540 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_245
timestamp 1688980957
transform 1 0 23644 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_251
timestamp 1688980957
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_253
timestamp 1688980957
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_265
timestamp 1688980957
transform 1 0 25484 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_277
timestamp 1688980957
transform 1 0 26588 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_289
timestamp 1688980957
transform 1 0 27692 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_301
timestamp 1688980957
transform 1 0 28796 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_307
timestamp 1688980957
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_309
timestamp 1688980957
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_321
timestamp 1688980957
transform 1 0 30636 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_333
timestamp 1688980957
transform 1 0 31740 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_345
timestamp 1688980957
transform 1 0 32844 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_357
timestamp 1688980957
transform 1 0 33948 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_363
timestamp 1688980957
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_3
timestamp 1688980957
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_15
timestamp 1688980957
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_27
timestamp 1688980957
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_39
timestamp 1688980957
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_51
timestamp 1688980957
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_55
timestamp 1688980957
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_57
timestamp 1688980957
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_69
timestamp 1688980957
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_81
timestamp 1688980957
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_93
timestamp 1688980957
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_105
timestamp 1688980957
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_111
timestamp 1688980957
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_113
timestamp 1688980957
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_125
timestamp 1688980957
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_137
timestamp 1688980957
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_149
timestamp 1688980957
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_161
timestamp 1688980957
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_167
timestamp 1688980957
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_169
timestamp 1688980957
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_181
timestamp 1688980957
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_193
timestamp 1688980957
transform 1 0 18860 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_205
timestamp 1688980957
transform 1 0 19964 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_217
timestamp 1688980957
transform 1 0 21068 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_223
timestamp 1688980957
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_225
timestamp 1688980957
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_237
timestamp 1688980957
transform 1 0 22908 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_249
timestamp 1688980957
transform 1 0 24012 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_261
timestamp 1688980957
transform 1 0 25116 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_273
timestamp 1688980957
transform 1 0 26220 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_279
timestamp 1688980957
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_281
timestamp 1688980957
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_293
timestamp 1688980957
transform 1 0 28060 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_305
timestamp 1688980957
transform 1 0 29164 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_317
timestamp 1688980957
transform 1 0 30268 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_329
timestamp 1688980957
transform 1 0 31372 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_335
timestamp 1688980957
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_337
timestamp 1688980957
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_349
timestamp 1688980957
transform 1 0 33212 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_361
timestamp 1688980957
transform 1 0 34316 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_3
timestamp 1688980957
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_15
timestamp 1688980957
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_27
timestamp 1688980957
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_29
timestamp 1688980957
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_41
timestamp 1688980957
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_53
timestamp 1688980957
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_65
timestamp 1688980957
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_77
timestamp 1688980957
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_83
timestamp 1688980957
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_85
timestamp 1688980957
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_97
timestamp 1688980957
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_109
timestamp 1688980957
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_121
timestamp 1688980957
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_133
timestamp 1688980957
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_139
timestamp 1688980957
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_141
timestamp 1688980957
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_153
timestamp 1688980957
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_165
timestamp 1688980957
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_177
timestamp 1688980957
transform 1 0 17388 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_189
timestamp 1688980957
transform 1 0 18492 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_195
timestamp 1688980957
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_197
timestamp 1688980957
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_209
timestamp 1688980957
transform 1 0 20332 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_221
timestamp 1688980957
transform 1 0 21436 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_233
timestamp 1688980957
transform 1 0 22540 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_245
timestamp 1688980957
transform 1 0 23644 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_251
timestamp 1688980957
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_253
timestamp 1688980957
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_265
timestamp 1688980957
transform 1 0 25484 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_277
timestamp 1688980957
transform 1 0 26588 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_289
timestamp 1688980957
transform 1 0 27692 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_301
timestamp 1688980957
transform 1 0 28796 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_307
timestamp 1688980957
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_309
timestamp 1688980957
transform 1 0 29532 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_321
timestamp 1688980957
transform 1 0 30636 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_333
timestamp 1688980957
transform 1 0 31740 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_345
timestamp 1688980957
transform 1 0 32844 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_357
timestamp 1688980957
transform 1 0 33948 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_363
timestamp 1688980957
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_3
timestamp 1688980957
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_15
timestamp 1688980957
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_27
timestamp 1688980957
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_39
timestamp 1688980957
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_51
timestamp 1688980957
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_55
timestamp 1688980957
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_57
timestamp 1688980957
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_69
timestamp 1688980957
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_81
timestamp 1688980957
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_93
timestamp 1688980957
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_105
timestamp 1688980957
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_111
timestamp 1688980957
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_113
timestamp 1688980957
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_125
timestamp 1688980957
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_137
timestamp 1688980957
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_149
timestamp 1688980957
transform 1 0 14812 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_161
timestamp 1688980957
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_167
timestamp 1688980957
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_169
timestamp 1688980957
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_181
timestamp 1688980957
transform 1 0 17756 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_193
timestamp 1688980957
transform 1 0 18860 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_205
timestamp 1688980957
transform 1 0 19964 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_217
timestamp 1688980957
transform 1 0 21068 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_223
timestamp 1688980957
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_225
timestamp 1688980957
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_237
timestamp 1688980957
transform 1 0 22908 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_249
timestamp 1688980957
transform 1 0 24012 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_261
timestamp 1688980957
transform 1 0 25116 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_273
timestamp 1688980957
transform 1 0 26220 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_279
timestamp 1688980957
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_281
timestamp 1688980957
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_293
timestamp 1688980957
transform 1 0 28060 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_305
timestamp 1688980957
transform 1 0 29164 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_317
timestamp 1688980957
transform 1 0 30268 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_329
timestamp 1688980957
transform 1 0 31372 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_335
timestamp 1688980957
transform 1 0 31924 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_337
timestamp 1688980957
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_349
timestamp 1688980957
transform 1 0 33212 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_361
timestamp 1688980957
transform 1 0 34316 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_3
timestamp 1688980957
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_15
timestamp 1688980957
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_27
timestamp 1688980957
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_29
timestamp 1688980957
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_41
timestamp 1688980957
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_53
timestamp 1688980957
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_65
timestamp 1688980957
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_77
timestamp 1688980957
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_83
timestamp 1688980957
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_85
timestamp 1688980957
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_97
timestamp 1688980957
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_109
timestamp 1688980957
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_121
timestamp 1688980957
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_133
timestamp 1688980957
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_139
timestamp 1688980957
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_141
timestamp 1688980957
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_153
timestamp 1688980957
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_165
timestamp 1688980957
transform 1 0 16284 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_177
timestamp 1688980957
transform 1 0 17388 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_189
timestamp 1688980957
transform 1 0 18492 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_195
timestamp 1688980957
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_197
timestamp 1688980957
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_209
timestamp 1688980957
transform 1 0 20332 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_221
timestamp 1688980957
transform 1 0 21436 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_233
timestamp 1688980957
transform 1 0 22540 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_245
timestamp 1688980957
transform 1 0 23644 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_251
timestamp 1688980957
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_253
timestamp 1688980957
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_265
timestamp 1688980957
transform 1 0 25484 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_277
timestamp 1688980957
transform 1 0 26588 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_289
timestamp 1688980957
transform 1 0 27692 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_301
timestamp 1688980957
transform 1 0 28796 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_307
timestamp 1688980957
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_309
timestamp 1688980957
transform 1 0 29532 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_321
timestamp 1688980957
transform 1 0 30636 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_333
timestamp 1688980957
transform 1 0 31740 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_345
timestamp 1688980957
transform 1 0 32844 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_357
timestamp 1688980957
transform 1 0 33948 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_363
timestamp 1688980957
transform 1 0 34500 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_3
timestamp 1688980957
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_15
timestamp 1688980957
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_27
timestamp 1688980957
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_39
timestamp 1688980957
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_51
timestamp 1688980957
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_55
timestamp 1688980957
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_57
timestamp 1688980957
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_69
timestamp 1688980957
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_81
timestamp 1688980957
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_93
timestamp 1688980957
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_105
timestamp 1688980957
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_111
timestamp 1688980957
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_113
timestamp 1688980957
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_125
timestamp 1688980957
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_137
timestamp 1688980957
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_149
timestamp 1688980957
transform 1 0 14812 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_161
timestamp 1688980957
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_167
timestamp 1688980957
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_169
timestamp 1688980957
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_181
timestamp 1688980957
transform 1 0 17756 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_193
timestamp 1688980957
transform 1 0 18860 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_205
timestamp 1688980957
transform 1 0 19964 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_217
timestamp 1688980957
transform 1 0 21068 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_223
timestamp 1688980957
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_225
timestamp 1688980957
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_237
timestamp 1688980957
transform 1 0 22908 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_249
timestamp 1688980957
transform 1 0 24012 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_261
timestamp 1688980957
transform 1 0 25116 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_273
timestamp 1688980957
transform 1 0 26220 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_279
timestamp 1688980957
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_281
timestamp 1688980957
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_293
timestamp 1688980957
transform 1 0 28060 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_305
timestamp 1688980957
transform 1 0 29164 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_317
timestamp 1688980957
transform 1 0 30268 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_329
timestamp 1688980957
transform 1 0 31372 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_335
timestamp 1688980957
transform 1 0 31924 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_337
timestamp 1688980957
transform 1 0 32108 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_349
timestamp 1688980957
transform 1 0 33212 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_361
timestamp 1688980957
transform 1 0 34316 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_3
timestamp 1688980957
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_15
timestamp 1688980957
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_27
timestamp 1688980957
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_29
timestamp 1688980957
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_41
timestamp 1688980957
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_53
timestamp 1688980957
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_65
timestamp 1688980957
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_77
timestamp 1688980957
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_83
timestamp 1688980957
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_85
timestamp 1688980957
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_97
timestamp 1688980957
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_109
timestamp 1688980957
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_121
timestamp 1688980957
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_133
timestamp 1688980957
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_139
timestamp 1688980957
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_141
timestamp 1688980957
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_153
timestamp 1688980957
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_165
timestamp 1688980957
transform 1 0 16284 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_177
timestamp 1688980957
transform 1 0 17388 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_189
timestamp 1688980957
transform 1 0 18492 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_195
timestamp 1688980957
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_197
timestamp 1688980957
transform 1 0 19228 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_209
timestamp 1688980957
transform 1 0 20332 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_221
timestamp 1688980957
transform 1 0 21436 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_233
timestamp 1688980957
transform 1 0 22540 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_245
timestamp 1688980957
transform 1 0 23644 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_251
timestamp 1688980957
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_253
timestamp 1688980957
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_265
timestamp 1688980957
transform 1 0 25484 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_277
timestamp 1688980957
transform 1 0 26588 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_289
timestamp 1688980957
transform 1 0 27692 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_301
timestamp 1688980957
transform 1 0 28796 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_307
timestamp 1688980957
transform 1 0 29348 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_309
timestamp 1688980957
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_321
timestamp 1688980957
transform 1 0 30636 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_333
timestamp 1688980957
transform 1 0 31740 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_345
timestamp 1688980957
transform 1 0 32844 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_357
timestamp 1688980957
transform 1 0 33948 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_363
timestamp 1688980957
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_3
timestamp 1688980957
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_15
timestamp 1688980957
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_27
timestamp 1688980957
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_39
timestamp 1688980957
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_51
timestamp 1688980957
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_55
timestamp 1688980957
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_57
timestamp 1688980957
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_69
timestamp 1688980957
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_81
timestamp 1688980957
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_93
timestamp 1688980957
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_105
timestamp 1688980957
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_111
timestamp 1688980957
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_113
timestamp 1688980957
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_125
timestamp 1688980957
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_137
timestamp 1688980957
transform 1 0 13708 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_149
timestamp 1688980957
transform 1 0 14812 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_161
timestamp 1688980957
transform 1 0 15916 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_167
timestamp 1688980957
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_169
timestamp 1688980957
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_181
timestamp 1688980957
transform 1 0 17756 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_193
timestamp 1688980957
transform 1 0 18860 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_205
timestamp 1688980957
transform 1 0 19964 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_217
timestamp 1688980957
transform 1 0 21068 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_223
timestamp 1688980957
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_225
timestamp 1688980957
transform 1 0 21804 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_237
timestamp 1688980957
transform 1 0 22908 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_249
timestamp 1688980957
transform 1 0 24012 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_261
timestamp 1688980957
transform 1 0 25116 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_273
timestamp 1688980957
transform 1 0 26220 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_279
timestamp 1688980957
transform 1 0 26772 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_281
timestamp 1688980957
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_293
timestamp 1688980957
transform 1 0 28060 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_305
timestamp 1688980957
transform 1 0 29164 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_317
timestamp 1688980957
transform 1 0 30268 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_329
timestamp 1688980957
transform 1 0 31372 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_335
timestamp 1688980957
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_337
timestamp 1688980957
transform 1 0 32108 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_349
timestamp 1688980957
transform 1 0 33212 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_361
timestamp 1688980957
transform 1 0 34316 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_3
timestamp 1688980957
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_15
timestamp 1688980957
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_27
timestamp 1688980957
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_29
timestamp 1688980957
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_41
timestamp 1688980957
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_53
timestamp 1688980957
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_65
timestamp 1688980957
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_77
timestamp 1688980957
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_83
timestamp 1688980957
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_85
timestamp 1688980957
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_97
timestamp 1688980957
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_109
timestamp 1688980957
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_121
timestamp 1688980957
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_133
timestamp 1688980957
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_139
timestamp 1688980957
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_141
timestamp 1688980957
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_153
timestamp 1688980957
transform 1 0 15180 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_165
timestamp 1688980957
transform 1 0 16284 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_177
timestamp 1688980957
transform 1 0 17388 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_189
timestamp 1688980957
transform 1 0 18492 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_195
timestamp 1688980957
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_197
timestamp 1688980957
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_209
timestamp 1688980957
transform 1 0 20332 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_221
timestamp 1688980957
transform 1 0 21436 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_233
timestamp 1688980957
transform 1 0 22540 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_245
timestamp 1688980957
transform 1 0 23644 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_251
timestamp 1688980957
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_253
timestamp 1688980957
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_265
timestamp 1688980957
transform 1 0 25484 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_277
timestamp 1688980957
transform 1 0 26588 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_289
timestamp 1688980957
transform 1 0 27692 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_301
timestamp 1688980957
transform 1 0 28796 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_307
timestamp 1688980957
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_309
timestamp 1688980957
transform 1 0 29532 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_321
timestamp 1688980957
transform 1 0 30636 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_333
timestamp 1688980957
transform 1 0 31740 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_345
timestamp 1688980957
transform 1 0 32844 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_357
timestamp 1688980957
transform 1 0 33948 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_3
timestamp 1688980957
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_15
timestamp 1688980957
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_27
timestamp 1688980957
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_39
timestamp 1688980957
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_51
timestamp 1688980957
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_55
timestamp 1688980957
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_57
timestamp 1688980957
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_69
timestamp 1688980957
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_81
timestamp 1688980957
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_93
timestamp 1688980957
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_105
timestamp 1688980957
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_111
timestamp 1688980957
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_113
timestamp 1688980957
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_125
timestamp 1688980957
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_137
timestamp 1688980957
transform 1 0 13708 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_149
timestamp 1688980957
transform 1 0 14812 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_161
timestamp 1688980957
transform 1 0 15916 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_167
timestamp 1688980957
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_169
timestamp 1688980957
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_181
timestamp 1688980957
transform 1 0 17756 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_193
timestamp 1688980957
transform 1 0 18860 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_205
timestamp 1688980957
transform 1 0 19964 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_217
timestamp 1688980957
transform 1 0 21068 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_223
timestamp 1688980957
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_225
timestamp 1688980957
transform 1 0 21804 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_237
timestamp 1688980957
transform 1 0 22908 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_249
timestamp 1688980957
transform 1 0 24012 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_261
timestamp 1688980957
transform 1 0 25116 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_273
timestamp 1688980957
transform 1 0 26220 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_279
timestamp 1688980957
transform 1 0 26772 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_281
timestamp 1688980957
transform 1 0 26956 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_293
timestamp 1688980957
transform 1 0 28060 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_305
timestamp 1688980957
transform 1 0 29164 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_317
timestamp 1688980957
transform 1 0 30268 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_329
timestamp 1688980957
transform 1 0 31372 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_335
timestamp 1688980957
transform 1 0 31924 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_337
timestamp 1688980957
transform 1 0 32108 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_349
timestamp 1688980957
transform 1 0 33212 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_361
timestamp 1688980957
transform 1 0 34316 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_6
timestamp 1688980957
transform 1 0 1656 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_18
timestamp 1688980957
transform 1 0 2760 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_26
timestamp 1688980957
transform 1 0 3496 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_29
timestamp 1688980957
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_41
timestamp 1688980957
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_53
timestamp 1688980957
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_65
timestamp 1688980957
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_77
timestamp 1688980957
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_83
timestamp 1688980957
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_85
timestamp 1688980957
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_97
timestamp 1688980957
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_109
timestamp 1688980957
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_121
timestamp 1688980957
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_133
timestamp 1688980957
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_139
timestamp 1688980957
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_141
timestamp 1688980957
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_153
timestamp 1688980957
transform 1 0 15180 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_165
timestamp 1688980957
transform 1 0 16284 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_177
timestamp 1688980957
transform 1 0 17388 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_189
timestamp 1688980957
transform 1 0 18492 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_195
timestamp 1688980957
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_197
timestamp 1688980957
transform 1 0 19228 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_209
timestamp 1688980957
transform 1 0 20332 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_221
timestamp 1688980957
transform 1 0 21436 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_233
timestamp 1688980957
transform 1 0 22540 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_245
timestamp 1688980957
transform 1 0 23644 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_251
timestamp 1688980957
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_253
timestamp 1688980957
transform 1 0 24380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_265
timestamp 1688980957
transform 1 0 25484 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_277
timestamp 1688980957
transform 1 0 26588 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_289
timestamp 1688980957
transform 1 0 27692 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_301
timestamp 1688980957
transform 1 0 28796 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_307
timestamp 1688980957
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_309
timestamp 1688980957
transform 1 0 29532 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_321
timestamp 1688980957
transform 1 0 30636 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_333
timestamp 1688980957
transform 1 0 31740 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_345
timestamp 1688980957
transform 1 0 32844 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_357
timestamp 1688980957
transform 1 0 33948 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_363
timestamp 1688980957
transform 1 0 34500 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_3
timestamp 1688980957
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_15
timestamp 1688980957
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_27
timestamp 1688980957
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_39
timestamp 1688980957
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_51
timestamp 1688980957
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_55
timestamp 1688980957
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_57
timestamp 1688980957
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_69
timestamp 1688980957
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_81
timestamp 1688980957
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_93
timestamp 1688980957
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_105
timestamp 1688980957
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_111
timestamp 1688980957
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_113
timestamp 1688980957
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_125
timestamp 1688980957
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_137
timestamp 1688980957
transform 1 0 13708 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_149
timestamp 1688980957
transform 1 0 14812 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_161
timestamp 1688980957
transform 1 0 15916 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_167
timestamp 1688980957
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_169
timestamp 1688980957
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_181
timestamp 1688980957
transform 1 0 17756 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_193
timestamp 1688980957
transform 1 0 18860 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_205
timestamp 1688980957
transform 1 0 19964 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_217
timestamp 1688980957
transform 1 0 21068 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_223
timestamp 1688980957
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_225
timestamp 1688980957
transform 1 0 21804 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_237
timestamp 1688980957
transform 1 0 22908 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_249
timestamp 1688980957
transform 1 0 24012 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_261
timestamp 1688980957
transform 1 0 25116 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_273
timestamp 1688980957
transform 1 0 26220 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_279
timestamp 1688980957
transform 1 0 26772 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_281
timestamp 1688980957
transform 1 0 26956 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_293
timestamp 1688980957
transform 1 0 28060 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_305
timestamp 1688980957
transform 1 0 29164 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_317
timestamp 1688980957
transform 1 0 30268 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_329
timestamp 1688980957
transform 1 0 31372 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_335
timestamp 1688980957
transform 1 0 31924 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_337
timestamp 1688980957
transform 1 0 32108 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_349
timestamp 1688980957
transform 1 0 33212 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_361
timestamp 1688980957
transform 1 0 34316 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_3
timestamp 1688980957
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_15
timestamp 1688980957
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_27
timestamp 1688980957
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_29
timestamp 1688980957
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_41
timestamp 1688980957
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_53
timestamp 1688980957
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_65
timestamp 1688980957
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_77
timestamp 1688980957
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_83
timestamp 1688980957
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_85
timestamp 1688980957
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_97
timestamp 1688980957
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_109
timestamp 1688980957
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_121
timestamp 1688980957
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_133
timestamp 1688980957
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_139
timestamp 1688980957
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_141
timestamp 1688980957
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_153
timestamp 1688980957
transform 1 0 15180 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_165
timestamp 1688980957
transform 1 0 16284 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_177
timestamp 1688980957
transform 1 0 17388 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_189
timestamp 1688980957
transform 1 0 18492 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_195
timestamp 1688980957
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_197
timestamp 1688980957
transform 1 0 19228 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_209
timestamp 1688980957
transform 1 0 20332 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_221
timestamp 1688980957
transform 1 0 21436 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_233
timestamp 1688980957
transform 1 0 22540 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_245
timestamp 1688980957
transform 1 0 23644 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_251
timestamp 1688980957
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_253
timestamp 1688980957
transform 1 0 24380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_265
timestamp 1688980957
transform 1 0 25484 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_277
timestamp 1688980957
transform 1 0 26588 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_289
timestamp 1688980957
transform 1 0 27692 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_301
timestamp 1688980957
transform 1 0 28796 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_307
timestamp 1688980957
transform 1 0 29348 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_309
timestamp 1688980957
transform 1 0 29532 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_321
timestamp 1688980957
transform 1 0 30636 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_333
timestamp 1688980957
transform 1 0 31740 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_345
timestamp 1688980957
transform 1 0 32844 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_357
timestamp 1688980957
transform 1 0 33948 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_363
timestamp 1688980957
transform 1 0 34500 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_3
timestamp 1688980957
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_15
timestamp 1688980957
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_27
timestamp 1688980957
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_39
timestamp 1688980957
transform 1 0 4692 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_51
timestamp 1688980957
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_55
timestamp 1688980957
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_57
timestamp 1688980957
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_69
timestamp 1688980957
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_81
timestamp 1688980957
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_93
timestamp 1688980957
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_105
timestamp 1688980957
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_111
timestamp 1688980957
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_113
timestamp 1688980957
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_125
timestamp 1688980957
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_137
timestamp 1688980957
transform 1 0 13708 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_149
timestamp 1688980957
transform 1 0 14812 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_161
timestamp 1688980957
transform 1 0 15916 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_167
timestamp 1688980957
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_169
timestamp 1688980957
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_181
timestamp 1688980957
transform 1 0 17756 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_193
timestamp 1688980957
transform 1 0 18860 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_205
timestamp 1688980957
transform 1 0 19964 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_217
timestamp 1688980957
transform 1 0 21068 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_223
timestamp 1688980957
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_225
timestamp 1688980957
transform 1 0 21804 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_237
timestamp 1688980957
transform 1 0 22908 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_249
timestamp 1688980957
transform 1 0 24012 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_261
timestamp 1688980957
transform 1 0 25116 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_273
timestamp 1688980957
transform 1 0 26220 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_279
timestamp 1688980957
transform 1 0 26772 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_281
timestamp 1688980957
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_293
timestamp 1688980957
transform 1 0 28060 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_305
timestamp 1688980957
transform 1 0 29164 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_317
timestamp 1688980957
transform 1 0 30268 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_329
timestamp 1688980957
transform 1 0 31372 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_335
timestamp 1688980957
transform 1 0 31924 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_337
timestamp 1688980957
transform 1 0 32108 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_349
timestamp 1688980957
transform 1 0 33212 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_361
timestamp 1688980957
transform 1 0 34316 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_3
timestamp 1688980957
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_15
timestamp 1688980957
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_27
timestamp 1688980957
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_29
timestamp 1688980957
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_41
timestamp 1688980957
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_53
timestamp 1688980957
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_65
timestamp 1688980957
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_77
timestamp 1688980957
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_83
timestamp 1688980957
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_85
timestamp 1688980957
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_97
timestamp 1688980957
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_109
timestamp 1688980957
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_121
timestamp 1688980957
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_133
timestamp 1688980957
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_139
timestamp 1688980957
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_141
timestamp 1688980957
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_153
timestamp 1688980957
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_165
timestamp 1688980957
transform 1 0 16284 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_177
timestamp 1688980957
transform 1 0 17388 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_189
timestamp 1688980957
transform 1 0 18492 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_195
timestamp 1688980957
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_197
timestamp 1688980957
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_209
timestamp 1688980957
transform 1 0 20332 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_221
timestamp 1688980957
transform 1 0 21436 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_233
timestamp 1688980957
transform 1 0 22540 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_245
timestamp 1688980957
transform 1 0 23644 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_251
timestamp 1688980957
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_253
timestamp 1688980957
transform 1 0 24380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_265
timestamp 1688980957
transform 1 0 25484 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_277
timestamp 1688980957
transform 1 0 26588 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_289
timestamp 1688980957
transform 1 0 27692 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_301
timestamp 1688980957
transform 1 0 28796 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_307
timestamp 1688980957
transform 1 0 29348 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_309
timestamp 1688980957
transform 1 0 29532 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_321
timestamp 1688980957
transform 1 0 30636 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_333
timestamp 1688980957
transform 1 0 31740 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_345
timestamp 1688980957
transform 1 0 32844 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_357
timestamp 1688980957
transform 1 0 33948 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_363
timestamp 1688980957
transform 1 0 34500 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_3
timestamp 1688980957
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_15
timestamp 1688980957
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_27
timestamp 1688980957
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_39
timestamp 1688980957
transform 1 0 4692 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_51
timestamp 1688980957
transform 1 0 5796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_55
timestamp 1688980957
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_57
timestamp 1688980957
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_69
timestamp 1688980957
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_81
timestamp 1688980957
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_93
timestamp 1688980957
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_105
timestamp 1688980957
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_111
timestamp 1688980957
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_113
timestamp 1688980957
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_125
timestamp 1688980957
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_137
timestamp 1688980957
transform 1 0 13708 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_149
timestamp 1688980957
transform 1 0 14812 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_161
timestamp 1688980957
transform 1 0 15916 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_167
timestamp 1688980957
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_169
timestamp 1688980957
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_181
timestamp 1688980957
transform 1 0 17756 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_193
timestamp 1688980957
transform 1 0 18860 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_205
timestamp 1688980957
transform 1 0 19964 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_217
timestamp 1688980957
transform 1 0 21068 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_223
timestamp 1688980957
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_225
timestamp 1688980957
transform 1 0 21804 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_237
timestamp 1688980957
transform 1 0 22908 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_249
timestamp 1688980957
transform 1 0 24012 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_261
timestamp 1688980957
transform 1 0 25116 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_273
timestamp 1688980957
transform 1 0 26220 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_279
timestamp 1688980957
transform 1 0 26772 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_281
timestamp 1688980957
transform 1 0 26956 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_293
timestamp 1688980957
transform 1 0 28060 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_305
timestamp 1688980957
transform 1 0 29164 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_317
timestamp 1688980957
transform 1 0 30268 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_329
timestamp 1688980957
transform 1 0 31372 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_335
timestamp 1688980957
transform 1 0 31924 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_337
timestamp 1688980957
transform 1 0 32108 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_349
timestamp 1688980957
transform 1 0 33212 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_361
timestamp 1688980957
transform 1 0 34316 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_3
timestamp 1688980957
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_15
timestamp 1688980957
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_27
timestamp 1688980957
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_29
timestamp 1688980957
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_41
timestamp 1688980957
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_53
timestamp 1688980957
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_65
timestamp 1688980957
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_77
timestamp 1688980957
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_83
timestamp 1688980957
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_85
timestamp 1688980957
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_97
timestamp 1688980957
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_109
timestamp 1688980957
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_121
timestamp 1688980957
transform 1 0 12236 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_133
timestamp 1688980957
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_139
timestamp 1688980957
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_141
timestamp 1688980957
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_153
timestamp 1688980957
transform 1 0 15180 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_165
timestamp 1688980957
transform 1 0 16284 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_177
timestamp 1688980957
transform 1 0 17388 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_189
timestamp 1688980957
transform 1 0 18492 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_195
timestamp 1688980957
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_197
timestamp 1688980957
transform 1 0 19228 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_209
timestamp 1688980957
transform 1 0 20332 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_221
timestamp 1688980957
transform 1 0 21436 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_233
timestamp 1688980957
transform 1 0 22540 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_245
timestamp 1688980957
transform 1 0 23644 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_251
timestamp 1688980957
transform 1 0 24196 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_253
timestamp 1688980957
transform 1 0 24380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_265
timestamp 1688980957
transform 1 0 25484 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_277
timestamp 1688980957
transform 1 0 26588 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_289
timestamp 1688980957
transform 1 0 27692 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_301
timestamp 1688980957
transform 1 0 28796 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_307
timestamp 1688980957
transform 1 0 29348 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_309
timestamp 1688980957
transform 1 0 29532 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_321
timestamp 1688980957
transform 1 0 30636 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_333
timestamp 1688980957
transform 1 0 31740 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_345
timestamp 1688980957
transform 1 0 32844 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_357
timestamp 1688980957
transform 1 0 33948 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_363
timestamp 1688980957
transform 1 0 34500 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_3
timestamp 1688980957
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_15
timestamp 1688980957
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_27
timestamp 1688980957
transform 1 0 3588 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_39
timestamp 1688980957
transform 1 0 4692 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_51
timestamp 1688980957
transform 1 0 5796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_55
timestamp 1688980957
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_57
timestamp 1688980957
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_69
timestamp 1688980957
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_81
timestamp 1688980957
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_93
timestamp 1688980957
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_105
timestamp 1688980957
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_111
timestamp 1688980957
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_113
timestamp 1688980957
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_125
timestamp 1688980957
transform 1 0 12604 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_137
timestamp 1688980957
transform 1 0 13708 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_149
timestamp 1688980957
transform 1 0 14812 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_161
timestamp 1688980957
transform 1 0 15916 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_167
timestamp 1688980957
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_169
timestamp 1688980957
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_181
timestamp 1688980957
transform 1 0 17756 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_193
timestamp 1688980957
transform 1 0 18860 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_205
timestamp 1688980957
transform 1 0 19964 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_217
timestamp 1688980957
transform 1 0 21068 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_223
timestamp 1688980957
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_225
timestamp 1688980957
transform 1 0 21804 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_237
timestamp 1688980957
transform 1 0 22908 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_249
timestamp 1688980957
transform 1 0 24012 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_261
timestamp 1688980957
transform 1 0 25116 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_273
timestamp 1688980957
transform 1 0 26220 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_279
timestamp 1688980957
transform 1 0 26772 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_281
timestamp 1688980957
transform 1 0 26956 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_293
timestamp 1688980957
transform 1 0 28060 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_305
timestamp 1688980957
transform 1 0 29164 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_317
timestamp 1688980957
transform 1 0 30268 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_329
timestamp 1688980957
transform 1 0 31372 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_335
timestamp 1688980957
transform 1 0 31924 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_337
timestamp 1688980957
transform 1 0 32108 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_349
timestamp 1688980957
transform 1 0 33212 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_361
timestamp 1688980957
transform 1 0 34316 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_3
timestamp 1688980957
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_15
timestamp 1688980957
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_27
timestamp 1688980957
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_29
timestamp 1688980957
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_41
timestamp 1688980957
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_53
timestamp 1688980957
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_65
timestamp 1688980957
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_77
timestamp 1688980957
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_83
timestamp 1688980957
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_85
timestamp 1688980957
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_97
timestamp 1688980957
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_109
timestamp 1688980957
transform 1 0 11132 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_121
timestamp 1688980957
transform 1 0 12236 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_133
timestamp 1688980957
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_139
timestamp 1688980957
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_141
timestamp 1688980957
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_153
timestamp 1688980957
transform 1 0 15180 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_165
timestamp 1688980957
transform 1 0 16284 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_177
timestamp 1688980957
transform 1 0 17388 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_189
timestamp 1688980957
transform 1 0 18492 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_195
timestamp 1688980957
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_197
timestamp 1688980957
transform 1 0 19228 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_209
timestamp 1688980957
transform 1 0 20332 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_221
timestamp 1688980957
transform 1 0 21436 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_233
timestamp 1688980957
transform 1 0 22540 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_245
timestamp 1688980957
transform 1 0 23644 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_251
timestamp 1688980957
transform 1 0 24196 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_253
timestamp 1688980957
transform 1 0 24380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_265
timestamp 1688980957
transform 1 0 25484 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_277
timestamp 1688980957
transform 1 0 26588 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_289
timestamp 1688980957
transform 1 0 27692 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_301
timestamp 1688980957
transform 1 0 28796 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_307
timestamp 1688980957
transform 1 0 29348 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_309
timestamp 1688980957
transform 1 0 29532 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_321
timestamp 1688980957
transform 1 0 30636 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_333
timestamp 1688980957
transform 1 0 31740 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_345
timestamp 1688980957
transform 1 0 32844 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_357
timestamp 1688980957
transform 1 0 33948 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_363
timestamp 1688980957
transform 1 0 34500 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_3
timestamp 1688980957
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_15
timestamp 1688980957
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_27
timestamp 1688980957
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_39
timestamp 1688980957
transform 1 0 4692 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_51
timestamp 1688980957
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_55
timestamp 1688980957
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_57
timestamp 1688980957
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_69
timestamp 1688980957
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_81
timestamp 1688980957
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_93
timestamp 1688980957
transform 1 0 9660 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_101
timestamp 1688980957
transform 1 0 10396 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_111
timestamp 1688980957
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_126
timestamp 1688980957
transform 1 0 12696 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_138
timestamp 1688980957
transform 1 0 13800 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_142
timestamp 1688980957
transform 1 0 14168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_147
timestamp 1688980957
transform 1 0 14628 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_155
timestamp 1688980957
transform 1 0 15364 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_166
timestamp 1688980957
transform 1 0 16376 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_169
timestamp 1688980957
transform 1 0 16652 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_181
timestamp 1688980957
transform 1 0 17756 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_187
timestamp 1688980957
transform 1 0 18308 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_202
timestamp 1688980957
transform 1 0 19688 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_210
timestamp 1688980957
transform 1 0 20424 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_215
timestamp 1688980957
transform 1 0 20884 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_225
timestamp 1688980957
transform 1 0 21804 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_237
timestamp 1688980957
transform 1 0 22908 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_249
timestamp 1688980957
transform 1 0 24012 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_261
timestamp 1688980957
transform 1 0 25116 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_273
timestamp 1688980957
transform 1 0 26220 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_279
timestamp 1688980957
transform 1 0 26772 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_281
timestamp 1688980957
transform 1 0 26956 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_293
timestamp 1688980957
transform 1 0 28060 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_305
timestamp 1688980957
transform 1 0 29164 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_317
timestamp 1688980957
transform 1 0 30268 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_329
timestamp 1688980957
transform 1 0 31372 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_335
timestamp 1688980957
transform 1 0 31924 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_337
timestamp 1688980957
transform 1 0 32108 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_349
timestamp 1688980957
transform 1 0 33212 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_361
timestamp 1688980957
transform 1 0 34316 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_3
timestamp 1688980957
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_15
timestamp 1688980957
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_27
timestamp 1688980957
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_29
timestamp 1688980957
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_41
timestamp 1688980957
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_53
timestamp 1688980957
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_65
timestamp 1688980957
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_77
timestamp 1688980957
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_83
timestamp 1688980957
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_85
timestamp 1688980957
transform 1 0 8924 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_91
timestamp 1688980957
transform 1 0 9476 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_95
timestamp 1688980957
transform 1 0 9844 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_133
timestamp 1688980957
transform 1 0 13340 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_139
timestamp 1688980957
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_141
timestamp 1688980957
transform 1 0 14076 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_169
timestamp 1688980957
transform 1 0 16652 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_177
timestamp 1688980957
transform 1 0 17388 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_197
timestamp 1688980957
transform 1 0 19228 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_223
timestamp 1688980957
transform 1 0 21620 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_235
timestamp 1688980957
transform 1 0 22724 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_247
timestamp 1688980957
transform 1 0 23828 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_251
timestamp 1688980957
transform 1 0 24196 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_253
timestamp 1688980957
transform 1 0 24380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_265
timestamp 1688980957
transform 1 0 25484 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_277
timestamp 1688980957
transform 1 0 26588 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_289
timestamp 1688980957
transform 1 0 27692 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_301
timestamp 1688980957
transform 1 0 28796 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_307
timestamp 1688980957
transform 1 0 29348 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_309
timestamp 1688980957
transform 1 0 29532 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_321
timestamp 1688980957
transform 1 0 30636 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_333
timestamp 1688980957
transform 1 0 31740 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_345
timestamp 1688980957
transform 1 0 32844 0 1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_3
timestamp 1688980957
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_15
timestamp 1688980957
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_27
timestamp 1688980957
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_39
timestamp 1688980957
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_51
timestamp 1688980957
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_55
timestamp 1688980957
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_57
timestamp 1688980957
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_69
timestamp 1688980957
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_81
timestamp 1688980957
transform 1 0 8556 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_85
timestamp 1688980957
transform 1 0 8924 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_111
timestamp 1688980957
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_113
timestamp 1688980957
transform 1 0 11500 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_143
timestamp 1688980957
transform 1 0 14260 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_177
timestamp 1688980957
transform 1 0 17388 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_185
timestamp 1688980957
transform 1 0 18124 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_212
timestamp 1688980957
transform 1 0 20608 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_217
timestamp 1688980957
transform 1 0 21068 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_223
timestamp 1688980957
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_246
timestamp 1688980957
transform 1 0 23736 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_258
timestamp 1688980957
transform 1 0 24840 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_270
timestamp 1688980957
transform 1 0 25944 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_278
timestamp 1688980957
transform 1 0 26680 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_281
timestamp 1688980957
transform 1 0 26956 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_293
timestamp 1688980957
transform 1 0 28060 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_305
timestamp 1688980957
transform 1 0 29164 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_317
timestamp 1688980957
transform 1 0 30268 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_329
timestamp 1688980957
transform 1 0 31372 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_335
timestamp 1688980957
transform 1 0 31924 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_337
timestamp 1688980957
transform 1 0 32108 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_349
timestamp 1688980957
transform 1 0 33212 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_361
timestamp 1688980957
transform 1 0 34316 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_3
timestamp 1688980957
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_15
timestamp 1688980957
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_27
timestamp 1688980957
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_29
timestamp 1688980957
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_41
timestamp 1688980957
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_53
timestamp 1688980957
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_65
timestamp 1688980957
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_77
timestamp 1688980957
transform 1 0 8188 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_141
timestamp 1688980957
transform 1 0 14076 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_157
timestamp 1688980957
transform 1 0 15548 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_174
timestamp 1688980957
transform 1 0 17112 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_185
timestamp 1688980957
transform 1 0 18124 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_195
timestamp 1688980957
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_197
timestamp 1688980957
transform 1 0 19228 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_203
timestamp 1688980957
transform 1 0 19780 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_220
timestamp 1688980957
transform 1 0 21344 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_247
timestamp 1688980957
transform 1 0 23828 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_251
timestamp 1688980957
transform 1 0 24196 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_253
timestamp 1688980957
transform 1 0 24380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_265
timestamp 1688980957
transform 1 0 25484 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_277
timestamp 1688980957
transform 1 0 26588 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_289
timestamp 1688980957
transform 1 0 27692 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_301
timestamp 1688980957
transform 1 0 28796 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_307
timestamp 1688980957
transform 1 0 29348 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_309
timestamp 1688980957
transform 1 0 29532 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_321
timestamp 1688980957
transform 1 0 30636 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_333
timestamp 1688980957
transform 1 0 31740 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_345
timestamp 1688980957
transform 1 0 32844 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_357
timestamp 1688980957
transform 1 0 33948 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_363
timestamp 1688980957
transform 1 0 34500 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_3
timestamp 1688980957
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_15
timestamp 1688980957
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_27
timestamp 1688980957
transform 1 0 3588 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_39
timestamp 1688980957
transform 1 0 4692 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_51
timestamp 1688980957
transform 1 0 5796 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_55
timestamp 1688980957
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_57
timestamp 1688980957
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_69
timestamp 1688980957
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_81
timestamp 1688980957
transform 1 0 8556 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_99
timestamp 1688980957
transform 1 0 10212 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_110
timestamp 1688980957
transform 1 0 11224 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_121
timestamp 1688980957
transform 1 0 12236 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_146
timestamp 1688980957
transform 1 0 14536 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_201
timestamp 1688980957
transform 1 0 19596 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_213
timestamp 1688980957
transform 1 0 20700 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_222
timestamp 1688980957
transform 1 0 21528 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_235
timestamp 1688980957
transform 1 0 22724 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_245
timestamp 1688980957
transform 1 0 23644 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_257
timestamp 1688980957
transform 1 0 24748 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_269
timestamp 1688980957
transform 1 0 25852 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_277
timestamp 1688980957
transform 1 0 26588 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_281
timestamp 1688980957
transform 1 0 26956 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_293
timestamp 1688980957
transform 1 0 28060 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_305
timestamp 1688980957
transform 1 0 29164 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_317
timestamp 1688980957
transform 1 0 30268 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_329
timestamp 1688980957
transform 1 0 31372 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_335
timestamp 1688980957
transform 1 0 31924 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_337
timestamp 1688980957
transform 1 0 32108 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_349
timestamp 1688980957
transform 1 0 33212 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_361
timestamp 1688980957
transform 1 0 34316 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_19
timestamp 1688980957
transform 1 0 2852 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_27
timestamp 1688980957
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_29
timestamp 1688980957
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_41
timestamp 1688980957
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_53
timestamp 1688980957
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_65
timestamp 1688980957
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_77
timestamp 1688980957
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_83
timestamp 1688980957
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_111
timestamp 1688980957
transform 1 0 11316 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_116
timestamp 1688980957
transform 1 0 11776 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_126
timestamp 1688980957
transform 1 0 12696 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_134
timestamp 1688980957
transform 1 0 13432 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_156
timestamp 1688980957
transform 1 0 15456 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_171
timestamp 1688980957
transform 1 0 16836 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_210
timestamp 1688980957
transform 1 0 20424 0 1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_220
timestamp 1688980957
transform 1 0 21344 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_232
timestamp 1688980957
transform 1 0 22448 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_240
timestamp 1688980957
transform 1 0 23184 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_245
timestamp 1688980957
transform 1 0 23644 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_251
timestamp 1688980957
transform 1 0 24196 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_253
timestamp 1688980957
transform 1 0 24380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_265
timestamp 1688980957
transform 1 0 25484 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_277
timestamp 1688980957
transform 1 0 26588 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_289
timestamp 1688980957
transform 1 0 27692 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_301
timestamp 1688980957
transform 1 0 28796 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_307
timestamp 1688980957
transform 1 0 29348 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_309
timestamp 1688980957
transform 1 0 29532 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_321
timestamp 1688980957
transform 1 0 30636 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_333
timestamp 1688980957
transform 1 0 31740 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_345
timestamp 1688980957
transform 1 0 32844 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_357
timestamp 1688980957
transform 1 0 33948 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_363
timestamp 1688980957
transform 1 0 34500 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_3
timestamp 1688980957
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_15
timestamp 1688980957
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_27
timestamp 1688980957
transform 1 0 3588 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_39
timestamp 1688980957
transform 1 0 4692 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_51
timestamp 1688980957
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_55
timestamp 1688980957
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_57
timestamp 1688980957
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_69
timestamp 1688980957
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_81
timestamp 1688980957
transform 1 0 8556 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_93
timestamp 1688980957
transform 1 0 9660 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_107
timestamp 1688980957
transform 1 0 10948 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_111
timestamp 1688980957
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_113
timestamp 1688980957
transform 1 0 11500 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_121
timestamp 1688980957
transform 1 0 12236 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_126
timestamp 1688980957
transform 1 0 12696 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_130
timestamp 1688980957
transform 1 0 13064 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_138
timestamp 1688980957
transform 1 0 13800 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_169
timestamp 1688980957
transform 1 0 16652 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_208
timestamp 1688980957
transform 1 0 20240 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_212
timestamp 1688980957
transform 1 0 20608 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_220
timestamp 1688980957
transform 1 0 21344 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_225
timestamp 1688980957
transform 1 0 21804 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_255
timestamp 1688980957
transform 1 0 24564 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_267
timestamp 1688980957
transform 1 0 25668 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_279
timestamp 1688980957
transform 1 0 26772 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_281
timestamp 1688980957
transform 1 0 26956 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_293
timestamp 1688980957
transform 1 0 28060 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_305
timestamp 1688980957
transform 1 0 29164 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_317
timestamp 1688980957
transform 1 0 30268 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_329
timestamp 1688980957
transform 1 0 31372 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_335
timestamp 1688980957
transform 1 0 31924 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_337
timestamp 1688980957
transform 1 0 32108 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_349
timestamp 1688980957
transform 1 0 33212 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_361
timestamp 1688980957
transform 1 0 34316 0 -1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_3
timestamp 1688980957
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_15
timestamp 1688980957
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_27
timestamp 1688980957
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_29
timestamp 1688980957
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_41
timestamp 1688980957
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_53
timestamp 1688980957
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_65
timestamp 1688980957
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_77
timestamp 1688980957
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_83
timestamp 1688980957
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_85
timestamp 1688980957
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_97
timestamp 1688980957
transform 1 0 10028 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_101
timestamp 1688980957
transform 1 0 10396 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_105
timestamp 1688980957
transform 1 0 10764 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_141
timestamp 1688980957
transform 1 0 14076 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_158
timestamp 1688980957
transform 1 0 15640 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_167
timestamp 1688980957
transform 1 0 16468 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_184
timestamp 1688980957
transform 1 0 18032 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_202
timestamp 1688980957
transform 1 0 19688 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_208
timestamp 1688980957
transform 1 0 20240 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_212
timestamp 1688980957
transform 1 0 20608 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_236
timestamp 1688980957
transform 1 0 22816 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_250
timestamp 1688980957
transform 1 0 24104 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_253
timestamp 1688980957
transform 1 0 24380 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_257
timestamp 1688980957
transform 1 0 24748 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_261
timestamp 1688980957
transform 1 0 25116 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_273
timestamp 1688980957
transform 1 0 26220 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_285
timestamp 1688980957
transform 1 0 27324 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_297
timestamp 1688980957
transform 1 0 28428 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_305
timestamp 1688980957
transform 1 0 29164 0 1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_309
timestamp 1688980957
transform 1 0 29532 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_321
timestamp 1688980957
transform 1 0 30636 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_333
timestamp 1688980957
transform 1 0 31740 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_345
timestamp 1688980957
transform 1 0 32844 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_357
timestamp 1688980957
transform 1 0 33948 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_363
timestamp 1688980957
transform 1 0 34500 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_3
timestamp 1688980957
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_15
timestamp 1688980957
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_27
timestamp 1688980957
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_39
timestamp 1688980957
transform 1 0 4692 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_51
timestamp 1688980957
transform 1 0 5796 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_55
timestamp 1688980957
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_57
timestamp 1688980957
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_69
timestamp 1688980957
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_81
timestamp 1688980957
transform 1 0 8556 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_96
timestamp 1688980957
transform 1 0 9936 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_122
timestamp 1688980957
transform 1 0 12328 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_126
timestamp 1688980957
transform 1 0 12696 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_167
timestamp 1688980957
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_169
timestamp 1688980957
transform 1 0 16652 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_209
timestamp 1688980957
transform 1 0 20332 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_221
timestamp 1688980957
transform 1 0 21436 0 -1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_255
timestamp 1688980957
transform 1 0 24564 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_267
timestamp 1688980957
transform 1 0 25668 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_279
timestamp 1688980957
transform 1 0 26772 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_281
timestamp 1688980957
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_293
timestamp 1688980957
transform 1 0 28060 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_305
timestamp 1688980957
transform 1 0 29164 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_317
timestamp 1688980957
transform 1 0 30268 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_329
timestamp 1688980957
transform 1 0 31372 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_335
timestamp 1688980957
transform 1 0 31924 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_337
timestamp 1688980957
transform 1 0 32108 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_349
timestamp 1688980957
transform 1 0 33212 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_361
timestamp 1688980957
transform 1 0 34316 0 -1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_3
timestamp 1688980957
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_15
timestamp 1688980957
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_27
timestamp 1688980957
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_29
timestamp 1688980957
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_41
timestamp 1688980957
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_53
timestamp 1688980957
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_65
timestamp 1688980957
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_77
timestamp 1688980957
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_83
timestamp 1688980957
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_101
timestamp 1688980957
transform 1 0 10396 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_105
timestamp 1688980957
transform 1 0 10764 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_109
timestamp 1688980957
transform 1 0 11132 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_118
timestamp 1688980957
transform 1 0 11960 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_147
timestamp 1688980957
transform 1 0 14628 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_159
timestamp 1688980957
transform 1 0 15732 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_185
timestamp 1688980957
transform 1 0 18124 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_195
timestamp 1688980957
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_197
timestamp 1688980957
transform 1 0 19228 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_206
timestamp 1688980957
transform 1 0 20056 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_223
timestamp 1688980957
transform 1 0 21620 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_238
timestamp 1688980957
transform 1 0 23000 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_248
timestamp 1688980957
transform 1 0 23920 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_253
timestamp 1688980957
transform 1 0 24380 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_257
timestamp 1688980957
transform 1 0 24748 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_261
timestamp 1688980957
transform 1 0 25116 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_273
timestamp 1688980957
transform 1 0 26220 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_285
timestamp 1688980957
transform 1 0 27324 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_297
timestamp 1688980957
transform 1 0 28428 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_305
timestamp 1688980957
transform 1 0 29164 0 1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_309
timestamp 1688980957
transform 1 0 29532 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_321
timestamp 1688980957
transform 1 0 30636 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_333
timestamp 1688980957
transform 1 0 31740 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_345
timestamp 1688980957
transform 1 0 32844 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_357
timestamp 1688980957
transform 1 0 33948 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_363
timestamp 1688980957
transform 1 0 34500 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_3
timestamp 1688980957
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_15
timestamp 1688980957
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_27
timestamp 1688980957
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_39
timestamp 1688980957
transform 1 0 4692 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_51
timestamp 1688980957
transform 1 0 5796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_55
timestamp 1688980957
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_57
timestamp 1688980957
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_69
timestamp 1688980957
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_81
timestamp 1688980957
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_93
timestamp 1688980957
transform 1 0 9660 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_113
timestamp 1688980957
transform 1 0 11500 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_125
timestamp 1688980957
transform 1 0 12604 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_144
timestamp 1688980957
transform 1 0 14352 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_150
timestamp 1688980957
transform 1 0 14904 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_161
timestamp 1688980957
transform 1 0 15916 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_167
timestamp 1688980957
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_186
timestamp 1688980957
transform 1 0 18216 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_194
timestamp 1688980957
transform 1 0 18952 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_204
timestamp 1688980957
transform 1 0 19872 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_221
timestamp 1688980957
transform 1 0 21436 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_233
timestamp 1688980957
transform 1 0 22540 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_242
timestamp 1688980957
transform 1 0 23368 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_254
timestamp 1688980957
transform 1 0 24472 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_266
timestamp 1688980957
transform 1 0 25576 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_278
timestamp 1688980957
transform 1 0 26680 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_281
timestamp 1688980957
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_293
timestamp 1688980957
transform 1 0 28060 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_305
timestamp 1688980957
transform 1 0 29164 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_317
timestamp 1688980957
transform 1 0 30268 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_329
timestamp 1688980957
transform 1 0 31372 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_335
timestamp 1688980957
transform 1 0 31924 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_337
timestamp 1688980957
transform 1 0 32108 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_349
timestamp 1688980957
transform 1 0 33212 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_361
timestamp 1688980957
transform 1 0 34316 0 -1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_3
timestamp 1688980957
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_15
timestamp 1688980957
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_27
timestamp 1688980957
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_29
timestamp 1688980957
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_41
timestamp 1688980957
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_53
timestamp 1688980957
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_65
timestamp 1688980957
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_77
timestamp 1688980957
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_83
timestamp 1688980957
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_85
timestamp 1688980957
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_97
timestamp 1688980957
transform 1 0 10028 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_130
timestamp 1688980957
transform 1 0 13064 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_141
timestamp 1688980957
transform 1 0 14076 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_151
timestamp 1688980957
transform 1 0 14996 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_155
timestamp 1688980957
transform 1 0 15364 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_159
timestamp 1688980957
transform 1 0 15732 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_163
timestamp 1688980957
transform 1 0 16100 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_195
timestamp 1688980957
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_205
timestamp 1688980957
transform 1 0 19964 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_216
timestamp 1688980957
transform 1 0 20976 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_224
timestamp 1688980957
transform 1 0 21712 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_232
timestamp 1688980957
transform 1 0 22448 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_253
timestamp 1688980957
transform 1 0 24380 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_257
timestamp 1688980957
transform 1 0 24748 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_261
timestamp 1688980957
transform 1 0 25116 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_273
timestamp 1688980957
transform 1 0 26220 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_285
timestamp 1688980957
transform 1 0 27324 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_297
timestamp 1688980957
transform 1 0 28428 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_305
timestamp 1688980957
transform 1 0 29164 0 1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_309
timestamp 1688980957
transform 1 0 29532 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_321
timestamp 1688980957
transform 1 0 30636 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_333
timestamp 1688980957
transform 1 0 31740 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_345
timestamp 1688980957
transform 1 0 32844 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_357
timestamp 1688980957
transform 1 0 33948 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_363
timestamp 1688980957
transform 1 0 34500 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_3
timestamp 1688980957
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_15
timestamp 1688980957
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_27
timestamp 1688980957
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_39
timestamp 1688980957
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_51
timestamp 1688980957
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_55
timestamp 1688980957
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_57
timestamp 1688980957
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_69
timestamp 1688980957
transform 1 0 7452 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_93
timestamp 1688980957
transform 1 0 9660 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_101
timestamp 1688980957
transform 1 0 10396 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_116
timestamp 1688980957
transform 1 0 11776 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_120
timestamp 1688980957
transform 1 0 12144 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_133
timestamp 1688980957
transform 1 0 13340 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_140
timestamp 1688980957
transform 1 0 13984 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_185
timestamp 1688980957
transform 1 0 18124 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_218
timestamp 1688980957
transform 1 0 21160 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_225
timestamp 1688980957
transform 1 0 21804 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_252
timestamp 1688980957
transform 1 0 24288 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_264
timestamp 1688980957
transform 1 0 25392 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_276
timestamp 1688980957
transform 1 0 26496 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_281
timestamp 1688980957
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_293
timestamp 1688980957
transform 1 0 28060 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_305
timestamp 1688980957
transform 1 0 29164 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_317
timestamp 1688980957
transform 1 0 30268 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_329
timestamp 1688980957
transform 1 0 31372 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_335
timestamp 1688980957
transform 1 0 31924 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_337
timestamp 1688980957
transform 1 0 32108 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_349
timestamp 1688980957
transform 1 0 33212 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_361
timestamp 1688980957
transform 1 0 34316 0 -1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_3
timestamp 1688980957
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_15
timestamp 1688980957
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_27
timestamp 1688980957
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_29
timestamp 1688980957
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_41
timestamp 1688980957
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_53
timestamp 1688980957
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_65
timestamp 1688980957
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_77
timestamp 1688980957
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_83
timestamp 1688980957
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_85
timestamp 1688980957
transform 1 0 8924 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_93
timestamp 1688980957
transform 1 0 9660 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_125
timestamp 1688980957
transform 1 0 12604 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_138
timestamp 1688980957
transform 1 0 13800 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_141
timestamp 1688980957
transform 1 0 14076 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_147
timestamp 1688980957
transform 1 0 14628 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_164
timestamp 1688980957
transform 1 0 16192 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_178
timestamp 1688980957
transform 1 0 17480 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_244
timestamp 1688980957
transform 1 0 23552 0 1 26112
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_253
timestamp 1688980957
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_265
timestamp 1688980957
transform 1 0 25484 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_277
timestamp 1688980957
transform 1 0 26588 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_289
timestamp 1688980957
transform 1 0 27692 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_301
timestamp 1688980957
transform 1 0 28796 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_307
timestamp 1688980957
transform 1 0 29348 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_309
timestamp 1688980957
transform 1 0 29532 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_321
timestamp 1688980957
transform 1 0 30636 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_333
timestamp 1688980957
transform 1 0 31740 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_345
timestamp 1688980957
transform 1 0 32844 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_357
timestamp 1688980957
transform 1 0 33948 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_363
timestamp 1688980957
transform 1 0 34500 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_3
timestamp 1688980957
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_15
timestamp 1688980957
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_27
timestamp 1688980957
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_39
timestamp 1688980957
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_51
timestamp 1688980957
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_55
timestamp 1688980957
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_57
timestamp 1688980957
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_69
timestamp 1688980957
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_81
timestamp 1688980957
transform 1 0 8556 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_85
timestamp 1688980957
transform 1 0 8924 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_91
timestamp 1688980957
transform 1 0 9476 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_103
timestamp 1688980957
transform 1 0 10580 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_111
timestamp 1688980957
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_119
timestamp 1688980957
transform 1 0 12052 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_125
timestamp 1688980957
transform 1 0 12604 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_142
timestamp 1688980957
transform 1 0 14168 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_146
timestamp 1688980957
transform 1 0 14536 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_169
timestamp 1688980957
transform 1 0 16652 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_190
timestamp 1688980957
transform 1 0 18584 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_200
timestamp 1688980957
transform 1 0 19504 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_256
timestamp 1688980957
transform 1 0 24656 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_268
timestamp 1688980957
transform 1 0 25760 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_281
timestamp 1688980957
transform 1 0 26956 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_293
timestamp 1688980957
transform 1 0 28060 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_305
timestamp 1688980957
transform 1 0 29164 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_317
timestamp 1688980957
transform 1 0 30268 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_329
timestamp 1688980957
transform 1 0 31372 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_335
timestamp 1688980957
transform 1 0 31924 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_337
timestamp 1688980957
transform 1 0 32108 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_349
timestamp 1688980957
transform 1 0 33212 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_361
timestamp 1688980957
transform 1 0 34316 0 -1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_3
timestamp 1688980957
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_15
timestamp 1688980957
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_27
timestamp 1688980957
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_29
timestamp 1688980957
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_41
timestamp 1688980957
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_53
timestamp 1688980957
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_65
timestamp 1688980957
transform 1 0 7084 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_85
timestamp 1688980957
transform 1 0 8924 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_104
timestamp 1688980957
transform 1 0 10672 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_116
timestamp 1688980957
transform 1 0 11776 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_123
timestamp 1688980957
transform 1 0 12420 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_127
timestamp 1688980957
transform 1 0 12788 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_136
timestamp 1688980957
transform 1 0 13616 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_141
timestamp 1688980957
transform 1 0 14076 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_150
timestamp 1688980957
transform 1 0 14904 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_154
timestamp 1688980957
transform 1 0 15272 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_178
timestamp 1688980957
transform 1 0 17480 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_205
timestamp 1688980957
transform 1 0 19964 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_232
timestamp 1688980957
transform 1 0 22448 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_236
timestamp 1688980957
transform 1 0 22816 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_240
timestamp 1688980957
transform 1 0 23184 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_249
timestamp 1688980957
transform 1 0 24012 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_253
timestamp 1688980957
transform 1 0 24380 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_257
timestamp 1688980957
transform 1 0 24748 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_261
timestamp 1688980957
transform 1 0 25116 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_273
timestamp 1688980957
transform 1 0 26220 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_285
timestamp 1688980957
transform 1 0 27324 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_297
timestamp 1688980957
transform 1 0 28428 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_305
timestamp 1688980957
transform 1 0 29164 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_309
timestamp 1688980957
transform 1 0 29532 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_321
timestamp 1688980957
transform 1 0 30636 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_333
timestamp 1688980957
transform 1 0 31740 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_345
timestamp 1688980957
transform 1 0 32844 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_357
timestamp 1688980957
transform 1 0 33948 0 1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_3
timestamp 1688980957
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_15
timestamp 1688980957
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_27
timestamp 1688980957
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_39
timestamp 1688980957
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_51
timestamp 1688980957
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_55
timestamp 1688980957
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_57
timestamp 1688980957
transform 1 0 6348 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_63
timestamp 1688980957
transform 1 0 6900 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_94
timestamp 1688980957
transform 1 0 9752 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_111
timestamp 1688980957
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_118
timestamp 1688980957
transform 1 0 11960 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47_136
timestamp 1688980957
transform 1 0 13616 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_155
timestamp 1688980957
transform 1 0 15364 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_185
timestamp 1688980957
transform 1 0 18124 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_211
timestamp 1688980957
transform 1 0 20516 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_222
timestamp 1688980957
transform 1 0 21528 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_230
timestamp 1688980957
transform 1 0 22264 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_242
timestamp 1688980957
transform 1 0 23368 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_254
timestamp 1688980957
transform 1 0 24472 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_266
timestamp 1688980957
transform 1 0 25576 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_278
timestamp 1688980957
transform 1 0 26680 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_281
timestamp 1688980957
transform 1 0 26956 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_293
timestamp 1688980957
transform 1 0 28060 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_305
timestamp 1688980957
transform 1 0 29164 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_317
timestamp 1688980957
transform 1 0 30268 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_329
timestamp 1688980957
transform 1 0 31372 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_335
timestamp 1688980957
transform 1 0 31924 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_337
timestamp 1688980957
transform 1 0 32108 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_349
timestamp 1688980957
transform 1 0 33212 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47_361
timestamp 1688980957
transform 1 0 34316 0 -1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_3
timestamp 1688980957
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_15
timestamp 1688980957
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_27
timestamp 1688980957
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_29
timestamp 1688980957
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_41
timestamp 1688980957
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_53
timestamp 1688980957
transform 1 0 5980 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_60
timestamp 1688980957
transform 1 0 6624 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_85
timestamp 1688980957
transform 1 0 8924 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_97
timestamp 1688980957
transform 1 0 10028 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_114
timestamp 1688980957
transform 1 0 11592 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_141
timestamp 1688980957
transform 1 0 14076 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_178
timestamp 1688980957
transform 1 0 17480 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_187
timestamp 1688980957
transform 1 0 18308 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_197
timestamp 1688980957
transform 1 0 19228 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_221
timestamp 1688980957
transform 1 0 21436 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_244
timestamp 1688980957
transform 1 0 23552 0 1 28288
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_253
timestamp 1688980957
transform 1 0 24380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_265
timestamp 1688980957
transform 1 0 25484 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_277
timestamp 1688980957
transform 1 0 26588 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_289
timestamp 1688980957
transform 1 0 27692 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_301
timestamp 1688980957
transform 1 0 28796 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_307
timestamp 1688980957
transform 1 0 29348 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_309
timestamp 1688980957
transform 1 0 29532 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_321
timestamp 1688980957
transform 1 0 30636 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_333
timestamp 1688980957
transform 1 0 31740 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_345
timestamp 1688980957
transform 1 0 32844 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_357
timestamp 1688980957
transform 1 0 33948 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_363
timestamp 1688980957
transform 1 0 34500 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_6
timestamp 1688980957
transform 1 0 1656 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_18
timestamp 1688980957
transform 1 0 2760 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_30
timestamp 1688980957
transform 1 0 3864 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_42
timestamp 1688980957
transform 1 0 4968 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_50
timestamp 1688980957
transform 1 0 5704 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_57
timestamp 1688980957
transform 1 0 6348 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_127
timestamp 1688980957
transform 1 0 12788 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_133
timestamp 1688980957
transform 1 0 13340 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_137
timestamp 1688980957
transform 1 0 13708 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_220
timestamp 1688980957
transform 1 0 21344 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_254
timestamp 1688980957
transform 1 0 24472 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_266
timestamp 1688980957
transform 1 0 25576 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_278
timestamp 1688980957
transform 1 0 26680 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_281
timestamp 1688980957
transform 1 0 26956 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_293
timestamp 1688980957
transform 1 0 28060 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_305
timestamp 1688980957
transform 1 0 29164 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_317
timestamp 1688980957
transform 1 0 30268 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_329
timestamp 1688980957
transform 1 0 31372 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_335
timestamp 1688980957
transform 1 0 31924 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_337
timestamp 1688980957
transform 1 0 32108 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_349
timestamp 1688980957
transform 1 0 33212 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_361
timestamp 1688980957
transform 1 0 34316 0 -1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_3
timestamp 1688980957
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_15
timestamp 1688980957
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_27
timestamp 1688980957
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_29
timestamp 1688980957
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_41
timestamp 1688980957
transform 1 0 4876 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_50_49
timestamp 1688980957
transform 1 0 5612 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_57
timestamp 1688980957
transform 1 0 6348 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_50_65
timestamp 1688980957
transform 1 0 7084 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_93
timestamp 1688980957
transform 1 0 9660 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_135
timestamp 1688980957
transform 1 0 13524 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_139
timestamp 1688980957
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_192
timestamp 1688980957
transform 1 0 18768 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_202
timestamp 1688980957
transform 1 0 19688 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_250
timestamp 1688980957
transform 1 0 24104 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_253
timestamp 1688980957
transform 1 0 24380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_265
timestamp 1688980957
transform 1 0 25484 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_277
timestamp 1688980957
transform 1 0 26588 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_289
timestamp 1688980957
transform 1 0 27692 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_301
timestamp 1688980957
transform 1 0 28796 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_307
timestamp 1688980957
transform 1 0 29348 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_309
timestamp 1688980957
transform 1 0 29532 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_321
timestamp 1688980957
transform 1 0 30636 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_333
timestamp 1688980957
transform 1 0 31740 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_345
timestamp 1688980957
transform 1 0 32844 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_357
timestamp 1688980957
transform 1 0 33948 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_363
timestamp 1688980957
transform 1 0 34500 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_3
timestamp 1688980957
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_15
timestamp 1688980957
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_27
timestamp 1688980957
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_39
timestamp 1688980957
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_51
timestamp 1688980957
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_55
timestamp 1688980957
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_57
timestamp 1688980957
transform 1 0 6348 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_62
timestamp 1688980957
transform 1 0 6808 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_77
timestamp 1688980957
transform 1 0 8188 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_85
timestamp 1688980957
transform 1 0 8924 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_108
timestamp 1688980957
transform 1 0 11040 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_116
timestamp 1688980957
transform 1 0 11776 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_133
timestamp 1688980957
transform 1 0 13340 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_160
timestamp 1688980957
transform 1 0 15824 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_169
timestamp 1688980957
transform 1 0 16652 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_182
timestamp 1688980957
transform 1 0 17848 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_203
timestamp 1688980957
transform 1 0 19780 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_209
timestamp 1688980957
transform 1 0 20332 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_213
timestamp 1688980957
transform 1 0 20700 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_51_221
timestamp 1688980957
transform 1 0 21436 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_234
timestamp 1688980957
transform 1 0 22632 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_240
timestamp 1688980957
transform 1 0 23184 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_257
timestamp 1688980957
transform 1 0 24748 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_269
timestamp 1688980957
transform 1 0 25852 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_51_277
timestamp 1688980957
transform 1 0 26588 0 -1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_281
timestamp 1688980957
transform 1 0 26956 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_293
timestamp 1688980957
transform 1 0 28060 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_305
timestamp 1688980957
transform 1 0 29164 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_317
timestamp 1688980957
transform 1 0 30268 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_329
timestamp 1688980957
transform 1 0 31372 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_335
timestamp 1688980957
transform 1 0 31924 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_337
timestamp 1688980957
transform 1 0 32108 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_349
timestamp 1688980957
transform 1 0 33212 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_51_361
timestamp 1688980957
transform 1 0 34316 0 -1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_3
timestamp 1688980957
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_15
timestamp 1688980957
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_27
timestamp 1688980957
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_29
timestamp 1688980957
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_41
timestamp 1688980957
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_52_53
timestamp 1688980957
transform 1 0 5980 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_61
timestamp 1688980957
transform 1 0 6716 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_78
timestamp 1688980957
transform 1 0 8280 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52_129
timestamp 1688980957
transform 1 0 12972 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_133
timestamp 1688980957
transform 1 0 13340 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_151
timestamp 1688980957
transform 1 0 14996 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_176
timestamp 1688980957
transform 1 0 17296 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_197
timestamp 1688980957
transform 1 0 19228 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_239
timestamp 1688980957
transform 1 0 23092 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_52_249
timestamp 1688980957
transform 1 0 24012 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_253
timestamp 1688980957
transform 1 0 24380 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_260
timestamp 1688980957
transform 1 0 25024 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_272
timestamp 1688980957
transform 1 0 26128 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_284
timestamp 1688980957
transform 1 0 27232 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_296
timestamp 1688980957
transform 1 0 28336 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_309
timestamp 1688980957
transform 1 0 29532 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_321
timestamp 1688980957
transform 1 0 30636 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_333
timestamp 1688980957
transform 1 0 31740 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_345
timestamp 1688980957
transform 1 0 32844 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_357
timestamp 1688980957
transform 1 0 33948 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_363
timestamp 1688980957
transform 1 0 34500 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_3
timestamp 1688980957
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_15
timestamp 1688980957
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_27
timestamp 1688980957
transform 1 0 3588 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_39
timestamp 1688980957
transform 1 0 4692 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_51
timestamp 1688980957
transform 1 0 5796 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_55
timestamp 1688980957
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_57
timestamp 1688980957
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_69
timestamp 1688980957
transform 1 0 7452 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_96
timestamp 1688980957
transform 1 0 9936 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53_100
timestamp 1688980957
transform 1 0 10304 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53_110
timestamp 1688980957
transform 1 0 11224 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_163
timestamp 1688980957
transform 1 0 16100 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_167
timestamp 1688980957
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_169
timestamp 1688980957
transform 1 0 16652 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_173
timestamp 1688980957
transform 1 0 17020 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53_177
timestamp 1688980957
transform 1 0 17388 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_53_196
timestamp 1688980957
transform 1 0 19136 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_220
timestamp 1688980957
transform 1 0 21344 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_241
timestamp 1688980957
transform 1 0 23276 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53_255
timestamp 1688980957
transform 1 0 24564 0 -1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_266
timestamp 1688980957
transform 1 0 25576 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53_278
timestamp 1688980957
transform 1 0 26680 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_281
timestamp 1688980957
transform 1 0 26956 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_293
timestamp 1688980957
transform 1 0 28060 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_305
timestamp 1688980957
transform 1 0 29164 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_317
timestamp 1688980957
transform 1 0 30268 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_329
timestamp 1688980957
transform 1 0 31372 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_335
timestamp 1688980957
transform 1 0 31924 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_337
timestamp 1688980957
transform 1 0 32108 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_349
timestamp 1688980957
transform 1 0 33212 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53_361
timestamp 1688980957
transform 1 0 34316 0 -1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_3
timestamp 1688980957
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_15
timestamp 1688980957
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_27
timestamp 1688980957
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_29
timestamp 1688980957
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_41
timestamp 1688980957
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_53
timestamp 1688980957
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_54_65
timestamp 1688980957
transform 1 0 7084 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_54_101
timestamp 1688980957
transform 1 0 10396 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_105
timestamp 1688980957
transform 1 0 10764 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_130
timestamp 1688980957
transform 1 0 13064 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_54_141
timestamp 1688980957
transform 1 0 14076 0 1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_147
timestamp 1688980957
transform 1 0 14628 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_54_166
timestamp 1688980957
transform 1 0 16376 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_176
timestamp 1688980957
transform 1 0 17296 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_54_184
timestamp 1688980957
transform 1 0 18032 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_188
timestamp 1688980957
transform 1 0 18400 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_195
timestamp 1688980957
transform 1 0 19044 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_54_197
timestamp 1688980957
transform 1 0 19228 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_217
timestamp 1688980957
transform 1 0 21068 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_269
timestamp 1688980957
transform 1 0 25852 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_281
timestamp 1688980957
transform 1 0 26956 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_293
timestamp 1688980957
transform 1 0 28060 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_54_305
timestamp 1688980957
transform 1 0 29164 0 1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_309
timestamp 1688980957
transform 1 0 29532 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_321
timestamp 1688980957
transform 1 0 30636 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_333
timestamp 1688980957
transform 1 0 31740 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_345
timestamp 1688980957
transform 1 0 32844 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_357
timestamp 1688980957
transform 1 0 33948 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_363
timestamp 1688980957
transform 1 0 34500 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_3
timestamp 1688980957
transform 1 0 1380 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_15
timestamp 1688980957
transform 1 0 2484 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_27
timestamp 1688980957
transform 1 0 3588 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_39
timestamp 1688980957
transform 1 0 4692 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_55_51
timestamp 1688980957
transform 1 0 5796 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_55
timestamp 1688980957
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_55_57
timestamp 1688980957
transform 1 0 6348 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_55_65
timestamp 1688980957
transform 1 0 7084 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_111
timestamp 1688980957
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_55_129
timestamp 1688980957
transform 1 0 12972 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_55_152
timestamp 1688980957
transform 1 0 15088 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_55_166
timestamp 1688980957
transform 1 0 16376 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_55_219
timestamp 1688980957
transform 1 0 21252 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_223
timestamp 1688980957
transform 1 0 21620 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_273
timestamp 1688980957
transform 1 0 26220 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_279
timestamp 1688980957
transform 1 0 26772 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_281
timestamp 1688980957
transform 1 0 26956 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_293
timestamp 1688980957
transform 1 0 28060 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_305
timestamp 1688980957
transform 1 0 29164 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_317
timestamp 1688980957
transform 1 0 30268 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_329
timestamp 1688980957
transform 1 0 31372 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_335
timestamp 1688980957
transform 1 0 31924 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_337
timestamp 1688980957
transform 1 0 32108 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_349
timestamp 1688980957
transform 1 0 33212 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_55_361
timestamp 1688980957
transform 1 0 34316 0 -1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_3
timestamp 1688980957
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_15
timestamp 1688980957
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_27
timestamp 1688980957
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_29
timestamp 1688980957
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_41
timestamp 1688980957
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_53
timestamp 1688980957
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_65
timestamp 1688980957
transform 1 0 7084 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_101
timestamp 1688980957
transform 1 0 10396 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_110
timestamp 1688980957
transform 1 0 11224 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_56_122
timestamp 1688980957
transform 1 0 12328 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_56_157
timestamp 1688980957
transform 1 0 15548 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_56_170
timestamp 1688980957
transform 1 0 16744 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_56_194
timestamp 1688980957
transform 1 0 18952 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_56_221
timestamp 1688980957
transform 1 0 21436 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_56_233
timestamp 1688980957
transform 1 0 22540 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_237
timestamp 1688980957
transform 1 0 22908 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_251
timestamp 1688980957
transform 1 0 24196 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_264
timestamp 1688980957
transform 1 0 25392 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_276
timestamp 1688980957
transform 1 0 26496 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_288
timestamp 1688980957
transform 1 0 27600 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_56_300
timestamp 1688980957
transform 1 0 28704 0 1 32640
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_309
timestamp 1688980957
transform 1 0 29532 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_321
timestamp 1688980957
transform 1 0 30636 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_333
timestamp 1688980957
transform 1 0 31740 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_345
timestamp 1688980957
transform 1 0 32844 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_357
timestamp 1688980957
transform 1 0 33948 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_363
timestamp 1688980957
transform 1 0 34500 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_3
timestamp 1688980957
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_15
timestamp 1688980957
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_27
timestamp 1688980957
transform 1 0 3588 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_39
timestamp 1688980957
transform 1 0 4692 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57_51
timestamp 1688980957
transform 1 0 5796 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_55
timestamp 1688980957
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57_57
timestamp 1688980957
transform 1 0 6348 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_57_65
timestamp 1688980957
transform 1 0 7084 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_84
timestamp 1688980957
transform 1 0 8832 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_129
timestamp 1688980957
transform 1 0 12972 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57_164
timestamp 1688980957
transform 1 0 16192 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_175
timestamp 1688980957
transform 1 0 17204 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57_185
timestamp 1688980957
transform 1 0 18124 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_193
timestamp 1688980957
transform 1 0 18860 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57_216
timestamp 1688980957
transform 1 0 20976 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_233
timestamp 1688980957
transform 1 0 22540 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_258
timestamp 1688980957
transform 1 0 24840 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57_270
timestamp 1688980957
transform 1 0 25944 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57_278
timestamp 1688980957
transform 1 0 26680 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_281
timestamp 1688980957
transform 1 0 26956 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_293
timestamp 1688980957
transform 1 0 28060 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_305
timestamp 1688980957
transform 1 0 29164 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_317
timestamp 1688980957
transform 1 0 30268 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_329
timestamp 1688980957
transform 1 0 31372 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_335
timestamp 1688980957
transform 1 0 31924 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_337
timestamp 1688980957
transform 1 0 32108 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_349
timestamp 1688980957
transform 1 0 33212 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_57_361
timestamp 1688980957
transform 1 0 34316 0 -1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_3
timestamp 1688980957
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_15
timestamp 1688980957
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_27
timestamp 1688980957
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_29
timestamp 1688980957
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_41
timestamp 1688980957
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_53
timestamp 1688980957
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_65
timestamp 1688980957
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_77
timestamp 1688980957
transform 1 0 8188 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58_99
timestamp 1688980957
transform 1 0 10212 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_130
timestamp 1688980957
transform 1 0 13064 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58_146
timestamp 1688980957
transform 1 0 14536 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_58_164
timestamp 1688980957
transform 1 0 16192 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_168
timestamp 1688980957
transform 1 0 16560 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_58_172
timestamp 1688980957
transform 1 0 16928 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58_188
timestamp 1688980957
transform 1 0 18400 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58_194
timestamp 1688980957
transform 1 0 18952 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_197
timestamp 1688980957
transform 1 0 19228 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_251
timestamp 1688980957
transform 1 0 24196 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_258
timestamp 1688980957
transform 1 0 24840 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_270
timestamp 1688980957
transform 1 0 25944 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_282
timestamp 1688980957
transform 1 0 27048 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_294
timestamp 1688980957
transform 1 0 28152 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58_306
timestamp 1688980957
transform 1 0 29256 0 1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_309
timestamp 1688980957
transform 1 0 29532 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_321
timestamp 1688980957
transform 1 0 30636 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_333
timestamp 1688980957
transform 1 0 31740 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_345
timestamp 1688980957
transform 1 0 32844 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_357
timestamp 1688980957
transform 1 0 33948 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_363
timestamp 1688980957
transform 1 0 34500 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_3
timestamp 1688980957
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_15
timestamp 1688980957
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_27
timestamp 1688980957
transform 1 0 3588 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_39
timestamp 1688980957
transform 1 0 4692 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_59_51
timestamp 1688980957
transform 1 0 5796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_55
timestamp 1688980957
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_57
timestamp 1688980957
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_69
timestamp 1688980957
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_59_81
timestamp 1688980957
transform 1 0 8556 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_113
timestamp 1688980957
transform 1 0 11500 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_59_146
timestamp 1688980957
transform 1 0 14536 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_150
timestamp 1688980957
transform 1 0 14904 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_169
timestamp 1688980957
transform 1 0 16652 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_59_176
timestamp 1688980957
transform 1 0 17296 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_59_195
timestamp 1688980957
transform 1 0 19044 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_59_221
timestamp 1688980957
transform 1 0 21436 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_59_225
timestamp 1688980957
transform 1 0 21804 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_59_240
timestamp 1688980957
transform 1 0 23184 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_266
timestamp 1688980957
transform 1 0 25576 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_59_278
timestamp 1688980957
transform 1 0 26680 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_281
timestamp 1688980957
transform 1 0 26956 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_293
timestamp 1688980957
transform 1 0 28060 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_305
timestamp 1688980957
transform 1 0 29164 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_317
timestamp 1688980957
transform 1 0 30268 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_329
timestamp 1688980957
transform 1 0 31372 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_335
timestamp 1688980957
transform 1 0 31924 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_337
timestamp 1688980957
transform 1 0 32108 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_349
timestamp 1688980957
transform 1 0 33212 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_59_361
timestamp 1688980957
transform 1 0 34316 0 -1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_3
timestamp 1688980957
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_15
timestamp 1688980957
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_27
timestamp 1688980957
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_29
timestamp 1688980957
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_41
timestamp 1688980957
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_53
timestamp 1688980957
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_65
timestamp 1688980957
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_77
timestamp 1688980957
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_83
timestamp 1688980957
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_60_85
timestamp 1688980957
transform 1 0 8924 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_89
timestamp 1688980957
transform 1 0 9292 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_118
timestamp 1688980957
transform 1 0 11960 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_60_144
timestamp 1688980957
transform 1 0 14352 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_175
timestamp 1688980957
transform 1 0 17204 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_60_197
timestamp 1688980957
transform 1 0 19228 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_201
timestamp 1688980957
transform 1 0 19596 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_60_205
timestamp 1688980957
transform 1 0 19964 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_232
timestamp 1688980957
transform 1 0 22448 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_236
timestamp 1688980957
transform 1 0 22816 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_242
timestamp 1688980957
transform 1 0 23368 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_60_248
timestamp 1688980957
transform 1 0 23920 0 1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_253
timestamp 1688980957
transform 1 0 24380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_265
timestamp 1688980957
transform 1 0 25484 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_277
timestamp 1688980957
transform 1 0 26588 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_289
timestamp 1688980957
transform 1 0 27692 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_301
timestamp 1688980957
transform 1 0 28796 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_307
timestamp 1688980957
transform 1 0 29348 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_309
timestamp 1688980957
transform 1 0 29532 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_321
timestamp 1688980957
transform 1 0 30636 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_333
timestamp 1688980957
transform 1 0 31740 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_345
timestamp 1688980957
transform 1 0 32844 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_60_357
timestamp 1688980957
transform 1 0 33948 0 1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_3
timestamp 1688980957
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_15
timestamp 1688980957
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_27
timestamp 1688980957
transform 1 0 3588 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_39
timestamp 1688980957
transform 1 0 4692 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_61_51
timestamp 1688980957
transform 1 0 5796 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_55
timestamp 1688980957
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_57
timestamp 1688980957
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_69
timestamp 1688980957
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_61_81
timestamp 1688980957
transform 1 0 8556 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_108
timestamp 1688980957
transform 1 0 11040 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_61_113
timestamp 1688980957
transform 1 0 11500 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_61_118
timestamp 1688980957
transform 1 0 11960 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_61_141
timestamp 1688980957
transform 1 0 14076 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_61_165
timestamp 1688980957
transform 1 0 16284 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_169
timestamp 1688980957
transform 1 0 16652 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_176
timestamp 1688980957
transform 1 0 17296 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_223
timestamp 1688980957
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_253
timestamp 1688980957
transform 1 0 24380 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_265
timestamp 1688980957
transform 1 0 25484 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_61_277
timestamp 1688980957
transform 1 0 26588 0 -1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_281
timestamp 1688980957
transform 1 0 26956 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_293
timestamp 1688980957
transform 1 0 28060 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_305
timestamp 1688980957
transform 1 0 29164 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_317
timestamp 1688980957
transform 1 0 30268 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_329
timestamp 1688980957
transform 1 0 31372 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_335
timestamp 1688980957
transform 1 0 31924 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_337
timestamp 1688980957
transform 1 0 32108 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_349
timestamp 1688980957
transform 1 0 33212 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_61_361
timestamp 1688980957
transform 1 0 34316 0 -1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_6
timestamp 1688980957
transform 1 0 1656 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_62_18
timestamp 1688980957
transform 1 0 2760 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_62_26
timestamp 1688980957
transform 1 0 3496 0 1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_29
timestamp 1688980957
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_41
timestamp 1688980957
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_53
timestamp 1688980957
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_62_65
timestamp 1688980957
transform 1 0 7084 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_62_76
timestamp 1688980957
transform 1 0 8096 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_62_85
timestamp 1688980957
transform 1 0 8924 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_95
timestamp 1688980957
transform 1 0 9844 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_127
timestamp 1688980957
transform 1 0 12788 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_62_137
timestamp 1688980957
transform 1 0 13708 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_62_157
timestamp 1688980957
transform 1 0 15548 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_178
timestamp 1688980957
transform 1 0 17480 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_192
timestamp 1688980957
transform 1 0 18768 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_205
timestamp 1688980957
transform 1 0 19964 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_230
timestamp 1688980957
transform 1 0 22264 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_62_247
timestamp 1688980957
transform 1 0 23828 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_251
timestamp 1688980957
transform 1 0 24196 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_253
timestamp 1688980957
transform 1 0 24380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_265
timestamp 1688980957
transform 1 0 25484 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_277
timestamp 1688980957
transform 1 0 26588 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_289
timestamp 1688980957
transform 1 0 27692 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_301
timestamp 1688980957
transform 1 0 28796 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_307
timestamp 1688980957
transform 1 0 29348 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_309
timestamp 1688980957
transform 1 0 29532 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_321
timestamp 1688980957
transform 1 0 30636 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_333
timestamp 1688980957
transform 1 0 31740 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_345
timestamp 1688980957
transform 1 0 32844 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_357
timestamp 1688980957
transform 1 0 33948 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_363
timestamp 1688980957
transform 1 0 34500 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_3
timestamp 1688980957
transform 1 0 1380 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_15
timestamp 1688980957
transform 1 0 2484 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_27
timestamp 1688980957
transform 1 0 3588 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_39
timestamp 1688980957
transform 1 0 4692 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_63_51
timestamp 1688980957
transform 1 0 5796 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_55
timestamp 1688980957
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_57
timestamp 1688980957
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_63_73
timestamp 1688980957
transform 1 0 7820 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_63_113
timestamp 1688980957
transform 1 0 11500 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_63_148
timestamp 1688980957
transform 1 0 14720 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_156
timestamp 1688980957
transform 1 0 15456 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_185
timestamp 1688980957
transform 1 0 18124 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_209
timestamp 1688980957
transform 1 0 20332 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_223
timestamp 1688980957
transform 1 0 21620 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_225
timestamp 1688980957
transform 1 0 21804 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_258
timestamp 1688980957
transform 1 0 24840 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_63_270
timestamp 1688980957
transform 1 0 25944 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_63_278
timestamp 1688980957
transform 1 0 26680 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_281
timestamp 1688980957
transform 1 0 26956 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_293
timestamp 1688980957
transform 1 0 28060 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_305
timestamp 1688980957
transform 1 0 29164 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_317
timestamp 1688980957
transform 1 0 30268 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_329
timestamp 1688980957
transform 1 0 31372 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_335
timestamp 1688980957
transform 1 0 31924 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_337
timestamp 1688980957
transform 1 0 32108 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_349
timestamp 1688980957
transform 1 0 33212 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_63_361
timestamp 1688980957
transform 1 0 34316 0 -1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_3
timestamp 1688980957
transform 1 0 1380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_15
timestamp 1688980957
transform 1 0 2484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_27
timestamp 1688980957
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_29
timestamp 1688980957
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_41
timestamp 1688980957
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_64_53
timestamp 1688980957
transform 1 0 5980 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_64_61
timestamp 1688980957
transform 1 0 6716 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_85
timestamp 1688980957
transform 1 0 8924 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_91
timestamp 1688980957
transform 1 0 9476 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_64_146
timestamp 1688980957
transform 1 0 14536 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_150
timestamp 1688980957
transform 1 0 14904 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_64_218
timestamp 1688980957
transform 1 0 21160 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_222
timestamp 1688980957
transform 1 0 21528 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_239
timestamp 1688980957
transform 1 0 23092 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_251
timestamp 1688980957
transform 1 0 24196 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_253
timestamp 1688980957
transform 1 0 24380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_265
timestamp 1688980957
transform 1 0 25484 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_277
timestamp 1688980957
transform 1 0 26588 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_289
timestamp 1688980957
transform 1 0 27692 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_301
timestamp 1688980957
transform 1 0 28796 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_307
timestamp 1688980957
transform 1 0 29348 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_309
timestamp 1688980957
transform 1 0 29532 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_321
timestamp 1688980957
transform 1 0 30636 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_333
timestamp 1688980957
transform 1 0 31740 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_345
timestamp 1688980957
transform 1 0 32844 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_357
timestamp 1688980957
transform 1 0 33948 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_363
timestamp 1688980957
transform 1 0 34500 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_3
timestamp 1688980957
transform 1 0 1380 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_15
timestamp 1688980957
transform 1 0 2484 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_27
timestamp 1688980957
transform 1 0 3588 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_39
timestamp 1688980957
transform 1 0 4692 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_65_51
timestamp 1688980957
transform 1 0 5796 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_55
timestamp 1688980957
transform 1 0 6164 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_65_57
timestamp 1688980957
transform 1 0 6348 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_65_65
timestamp 1688980957
transform 1 0 7084 0 -1 38080
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_71
timestamp 1688980957
transform 1 0 7636 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_83
timestamp 1688980957
transform 1 0 8740 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_65_87
timestamp 1688980957
transform 1 0 9108 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_65_95
timestamp 1688980957
transform 1 0 9844 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_65_124
timestamp 1688980957
transform 1 0 12512 0 -1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_131
timestamp 1688980957
transform 1 0 13156 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_65_143
timestamp 1688980957
transform 1 0 14260 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_65_164
timestamp 1688980957
transform 1 0 16192 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_65_169
timestamp 1688980957
transform 1 0 16652 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_65_204
timestamp 1688980957
transform 1 0 19872 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_65_216
timestamp 1688980957
transform 1 0 20976 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_232
timestamp 1688980957
transform 1 0 22448 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_241
timestamp 1688980957
transform 1 0 23276 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_253
timestamp 1688980957
transform 1 0 24380 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_265
timestamp 1688980957
transform 1 0 25484 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_65_277
timestamp 1688980957
transform 1 0 26588 0 -1 38080
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_281
timestamp 1688980957
transform 1 0 26956 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_293
timestamp 1688980957
transform 1 0 28060 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_305
timestamp 1688980957
transform 1 0 29164 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_317
timestamp 1688980957
transform 1 0 30268 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_65_329
timestamp 1688980957
transform 1 0 31372 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_335
timestamp 1688980957
transform 1 0 31924 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_337
timestamp 1688980957
transform 1 0 32108 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_349
timestamp 1688980957
transform 1 0 33212 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_65_361
timestamp 1688980957
transform 1 0 34316 0 -1 38080
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_3
timestamp 1688980957
transform 1 0 1380 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_15
timestamp 1688980957
transform 1 0 2484 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_27
timestamp 1688980957
transform 1 0 3588 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_66_29
timestamp 1688980957
transform 1 0 3772 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_66_37
timestamp 1688980957
transform 1 0 4508 0 1 38080
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_48
timestamp 1688980957
transform 1 0 5520 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_60
timestamp 1688980957
transform 1 0 6624 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_72
timestamp 1688980957
transform 1 0 7728 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_83
timestamp 1688980957
transform 1 0 8740 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_85
timestamp 1688980957
transform 1 0 8924 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_97
timestamp 1688980957
transform 1 0 10028 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_109
timestamp 1688980957
transform 1 0 11132 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_121
timestamp 1688980957
transform 1 0 12236 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_66_133
timestamp 1688980957
transform 1 0 13340 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_141
timestamp 1688980957
transform 1 0 14076 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_66_158
timestamp 1688980957
transform 1 0 15640 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_66_176
timestamp 1688980957
transform 1 0 17296 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_66_186
timestamp 1688980957
transform 1 0 18216 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_66_197
timestamp 1688980957
transform 1 0 19228 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_66_217
timestamp 1688980957
transform 1 0 21068 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_245
timestamp 1688980957
transform 1 0 23644 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_251
timestamp 1688980957
transform 1 0 24196 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_253
timestamp 1688980957
transform 1 0 24380 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_265
timestamp 1688980957
transform 1 0 25484 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_277
timestamp 1688980957
transform 1 0 26588 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_289
timestamp 1688980957
transform 1 0 27692 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_301
timestamp 1688980957
transform 1 0 28796 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_307
timestamp 1688980957
transform 1 0 29348 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_309
timestamp 1688980957
transform 1 0 29532 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_321
timestamp 1688980957
transform 1 0 30636 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_333
timestamp 1688980957
transform 1 0 31740 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_345
timestamp 1688980957
transform 1 0 32844 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_357
timestamp 1688980957
transform 1 0 33948 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_363
timestamp 1688980957
transform 1 0 34500 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_11
timestamp 1688980957
transform 1 0 2116 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_23
timestamp 1688980957
transform 1 0 3220 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_35
timestamp 1688980957
transform 1 0 4324 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_67_47
timestamp 1688980957
transform 1 0 5428 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_55
timestamp 1688980957
transform 1 0 6164 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_57
timestamp 1688980957
transform 1 0 6348 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_69
timestamp 1688980957
transform 1 0 7452 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_81
timestamp 1688980957
transform 1 0 8556 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_93
timestamp 1688980957
transform 1 0 9660 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_105
timestamp 1688980957
transform 1 0 10764 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_111
timestamp 1688980957
transform 1 0 11316 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_113
timestamp 1688980957
transform 1 0 11500 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_125
timestamp 1688980957
transform 1 0 12604 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_137
timestamp 1688980957
transform 1 0 13708 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_190
timestamp 1688980957
transform 1 0 18584 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_67_202
timestamp 1688980957
transform 1 0 19688 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_206
timestamp 1688980957
transform 1 0 20056 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_223
timestamp 1688980957
transform 1 0 21620 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_249
timestamp 1688980957
transform 1 0 24012 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_261
timestamp 1688980957
transform 1 0 25116 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_273
timestamp 1688980957
transform 1 0 26220 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_279
timestamp 1688980957
transform 1 0 26772 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_281
timestamp 1688980957
transform 1 0 26956 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_293
timestamp 1688980957
transform 1 0 28060 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_305
timestamp 1688980957
transform 1 0 29164 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_317
timestamp 1688980957
transform 1 0 30268 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_329
timestamp 1688980957
transform 1 0 31372 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_335
timestamp 1688980957
transform 1 0 31924 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_337
timestamp 1688980957
transform 1 0 32108 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_349
timestamp 1688980957
transform 1 0 33212 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_67_361
timestamp 1688980957
transform 1 0 34316 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_6
timestamp 1688980957
transform 1 0 1656 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_68_23
timestamp 1688980957
transform 1 0 3220 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_27
timestamp 1688980957
transform 1 0 3588 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_29
timestamp 1688980957
transform 1 0 3772 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_41
timestamp 1688980957
transform 1 0 4876 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_68_53
timestamp 1688980957
transform 1 0 5980 0 1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_57
timestamp 1688980957
transform 1 0 6348 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_68_69
timestamp 1688980957
transform 1 0 7452 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_68_77
timestamp 1688980957
transform 1 0 8188 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_83
timestamp 1688980957
transform 1 0 8740 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_85
timestamp 1688980957
transform 1 0 8924 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_97
timestamp 1688980957
transform 1 0 10028 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_68_109
timestamp 1688980957
transform 1 0 11132 0 1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_113
timestamp 1688980957
transform 1 0 11500 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_125
timestamp 1688980957
transform 1 0 12604 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_68_137
timestamp 1688980957
transform 1 0 13708 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_68_141
timestamp 1688980957
transform 1 0 14076 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_68_148
timestamp 1688980957
transform 1 0 14720 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_153
timestamp 1688980957
transform 1 0 15180 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_167
timestamp 1688980957
transform 1 0 16468 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_68_169
timestamp 1688980957
transform 1 0 16652 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_68_174
timestamp 1688980957
transform 1 0 17112 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_68_187
timestamp 1688980957
transform 1 0 18308 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_195
timestamp 1688980957
transform 1 0 19044 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_197
timestamp 1688980957
transform 1 0 19228 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_68_209
timestamp 1688980957
transform 1 0 20332 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_68_214
timestamp 1688980957
transform 1 0 20792 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_218
timestamp 1688980957
transform 1 0 21160 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_68_222
timestamp 1688980957
transform 1 0 21528 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_68_225
timestamp 1688980957
transform 1 0 21804 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_68_243
timestamp 1688980957
transform 1 0 23460 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_251
timestamp 1688980957
transform 1 0 24196 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_253
timestamp 1688980957
transform 1 0 24380 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_265
timestamp 1688980957
transform 1 0 25484 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_68_277
timestamp 1688980957
transform 1 0 26588 0 1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_281
timestamp 1688980957
transform 1 0 26956 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_293
timestamp 1688980957
transform 1 0 28060 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_68_305
timestamp 1688980957
transform 1 0 29164 0 1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_309
timestamp 1688980957
transform 1 0 29532 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_321
timestamp 1688980957
transform 1 0 30636 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_68_333
timestamp 1688980957
transform 1 0 31740 0 1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_337
timestamp 1688980957
transform 1 0 32108 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_349
timestamp 1688980957
transform 1 0 33212 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 3220 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1688980957
transform 1 0 4784 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1688980957
transform -1 0 8740 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  hold4 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 15364 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1688980957
transform -1 0 14904 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  hold6 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 15456 0 -1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 1688980957
transform -1 0 17388 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 1688980957
transform 1 0 21804 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 1688980957
transform 1 0 21804 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp 1688980957
transform 1 0 20424 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp 1688980957
transform 1 0 20608 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold12
timestamp 1688980957
transform 1 0 10488 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp 1688980957
transform -1 0 12972 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold14
timestamp 1688980957
transform -1 0 18768 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold15
timestamp 1688980957
transform 1 0 15824 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold16
timestamp 1688980957
transform -1 0 14076 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold17
timestamp 1688980957
transform 1 0 13984 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  hold18
timestamp 1688980957
transform 1 0 17664 0 1 25024
box -38 -48 958 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold19
timestamp 1688980957
transform 1 0 15824 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold20
timestamp 1688980957
transform -1 0 9660 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold21
timestamp 1688980957
transform 1 0 10488 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold22
timestamp 1688980957
transform -1 0 20148 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold23
timestamp 1688980957
transform -1 0 19136 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold24
timestamp 1688980957
transform -1 0 18308 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold25
timestamp 1688980957
transform 1 0 16744 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold26
timestamp 1688980957
transform -1 0 19412 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold27
timestamp 1688980957
transform -1 0 18676 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold28
timestamp 1688980957
transform 1 0 12788 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold29
timestamp 1688980957
transform 1 0 12052 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold30
timestamp 1688980957
transform -1 0 10396 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold31
timestamp 1688980957
transform 1 0 8924 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  hold32
timestamp 1688980957
transform 1 0 15548 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold33
timestamp 1688980957
transform 1 0 14076 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold34
timestamp 1688980957
transform -1 0 21436 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold35
timestamp 1688980957
transform -1 0 20608 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold36
timestamp 1688980957
transform 1 0 15088 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold37
timestamp 1688980957
transform -1 0 16192 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  hold38
timestamp 1688980957
transform -1 0 16928 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold39
timestamp 1688980957
transform 1 0 18124 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold40
timestamp 1688980957
transform -1 0 18032 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  hold41
timestamp 1688980957
transform -1 0 17664 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold42
timestamp 1688980957
transform -1 0 16376 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold43
timestamp 1688980957
transform 1 0 14352 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold44
timestamp 1688980957
transform -1 0 19504 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold45
timestamp 1688980957
transform 1 0 17112 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold46
timestamp 1688980957
transform 1 0 9108 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold47
timestamp 1688980957
transform -1 0 19964 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold48
timestamp 1688980957
transform -1 0 20516 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold49
timestamp 1688980957
transform -1 0 12236 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold50
timestamp 1688980957
transform -1 0 11316 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold51
timestamp 1688980957
transform -1 0 19136 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold52
timestamp 1688980957
transform 1 0 16928 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold53
timestamp 1688980957
transform -1 0 10948 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold54
timestamp 1688980957
transform -1 0 10212 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold55
timestamp 1688980957
transform 1 0 15824 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold56
timestamp 1688980957
transform -1 0 11592 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold57
timestamp 1688980957
transform -1 0 9752 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold58
timestamp 1688980957
transform -1 0 9752 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold59
timestamp 1688980957
transform -1 0 20056 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold60
timestamp 1688980957
transform 1 0 21988 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold61
timestamp 1688980957
transform 1 0 11592 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold62
timestamp 1688980957
transform -1 0 9660 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold63
timestamp 1688980957
transform -1 0 14536 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold64
timestamp 1688980957
transform -1 0 11684 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold65
timestamp 1688980957
transform -1 0 9200 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold66
timestamp 1688980957
transform -1 0 9660 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold67
timestamp 1688980957
transform 1 0 17480 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold68
timestamp 1688980957
transform 1 0 21252 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold69
timestamp 1688980957
transform -1 0 26220 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold70
timestamp 1688980957
transform -1 0 25576 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold71
timestamp 1688980957
transform -1 0 8832 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold72
timestamp 1688980957
transform 1 0 24840 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold73
timestamp 1688980957
transform -1 0 25392 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold74
timestamp 1688980957
transform 1 0 11776 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold75
timestamp 1688980957
transform 1 0 23276 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold76
timestamp 1688980957
transform -1 0 10948 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold77
timestamp 1688980957
transform 1 0 16008 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold78
timestamp 1688980957
transform -1 0 16192 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold79
timestamp 1688980957
transform -1 0 14536 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold80
timestamp 1688980957
transform -1 0 13800 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold81
timestamp 1688980957
transform 1 0 8740 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold82
timestamp 1688980957
transform -1 0 17388 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold83
timestamp 1688980957
transform -1 0 18124 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold84
timestamp 1688980957
transform 1 0 8280 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold85
timestamp 1688980957
transform 1 0 21712 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold86
timestamp 1688980957
transform 1 0 20240 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold87
timestamp 1688980957
transform 1 0 22632 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold88
timestamp 1688980957
transform -1 0 16468 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold89
timestamp 1688980957
transform 1 0 10672 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold90
timestamp 1688980957
transform -1 0 12236 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold91
timestamp 1688980957
transform -1 0 12512 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold92
timestamp 1688980957
transform -1 0 11408 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold93
timestamp 1688980957
transform -1 0 12880 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold94
timestamp 1688980957
transform -1 0 23184 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold95
timestamp 1688980957
transform -1 0 19136 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold96
timestamp 1688980957
transform -1 0 23276 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold97
timestamp 1688980957
transform -1 0 23644 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold98
timestamp 1688980957
transform 1 0 22448 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold99
timestamp 1688980957
transform -1 0 22356 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold100
timestamp 1688980957
transform -1 0 10948 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold101
timestamp 1688980957
transform 1 0 13248 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold102
timestamp 1688980957
transform -1 0 21252 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold103
timestamp 1688980957
transform 1 0 20332 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold104
timestamp 1688980957
transform -1 0 24196 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold105 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 14260 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold106
timestamp 1688980957
transform -1 0 13616 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  hold107
timestamp 1688980957
transform 1 0 14352 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold108
timestamp 1688980957
transform -1 0 13984 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  hold109
timestamp 1688980957
transform -1 0 25116 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold110
timestamp 1688980957
transform 1 0 23276 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  hold111
timestamp 1688980957
transform -1 0 25116 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold112
timestamp 1688980957
transform 1 0 23184 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  hold113
timestamp 1688980957
transform -1 0 15180 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold114
timestamp 1688980957
transform -1 0 16560 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold115
timestamp 1688980957
transform 1 0 18400 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold116
timestamp 1688980957
transform -1 0 19688 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  hold117
timestamp 1688980957
transform -1 0 14904 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold118
timestamp 1688980957
transform 1 0 12880 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  hold119
timestamp 1688980957
transform -1 0 16928 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold120
timestamp 1688980957
transform -1 0 16008 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  hold121
timestamp 1688980957
transform -1 0 17388 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold122
timestamp 1688980957
transform 1 0 15088 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  hold123
timestamp 1688980957
transform -1 0 25116 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold124
timestamp 1688980957
transform -1 0 23920 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold125
timestamp 1688980957
transform -1 0 16468 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold126
timestamp 1688980957
transform 1 0 14904 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  hold127
timestamp 1688980957
transform -1 0 25116 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold128
timestamp 1688980957
transform 1 0 22908 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold129
timestamp 1688980957
transform -1 0 22540 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold130
timestamp 1688980957
transform -1 0 21068 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  hold131
timestamp 1688980957
transform 1 0 20792 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold132
timestamp 1688980957
transform -1 0 21528 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold133
timestamp 1688980957
transform -1 0 16928 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold134
timestamp 1688980957
transform 1 0 12236 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  hold135
timestamp 1688980957
transform 1 0 11500 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold136
timestamp 1688980957
transform -1 0 11408 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  hold137
timestamp 1688980957
transform 1 0 10488 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold138
timestamp 1688980957
transform -1 0 11960 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  hold139
timestamp 1688980957
transform 1 0 17756 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold140
timestamp 1688980957
transform 1 0 18400 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold141
timestamp 1688980957
transform -1 0 19964 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold142
timestamp 1688980957
transform 1 0 23276 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  hold143
timestamp 1688980957
transform -1 0 19964 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold144
timestamp 1688980957
transform 1 0 17756 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold145
timestamp 1688980957
transform -1 0 13064 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold146
timestamp 1688980957
transform 1 0 18216 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold147
timestamp 1688980957
transform 1 0 20700 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold148
timestamp 1688980957
transform 1 0 19780 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold149
timestamp 1688980957
transform 1 0 1380 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold150
timestamp 1688980957
transform -1 0 2484 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold151
timestamp 1688980957
transform 1 0 16100 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold152
timestamp 1688980957
transform 1 0 15824 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold153
timestamp 1688980957
transform -1 0 18584 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold154
timestamp 1688980957
transform 1 0 16376 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1688980957
transform 1 0 14904 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1688980957
transform 1 0 34316 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input3
timestamp 1688980957
transform -1 0 34592 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1688980957
transform 1 0 8464 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1688980957
transform -1 0 1656 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input6
timestamp 1688980957
transform 1 0 1380 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input7
timestamp 1688980957
transform 1 0 1380 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__buf_12  output8 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 21988 0 1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output9
timestamp 1688980957
transform 1 0 20240 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output10
timestamp 1688980957
transform -1 0 2852 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output11
timestamp 1688980957
transform 1 0 33120 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1688980957
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1688980957
transform -1 0 34868 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1688980957
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1688980957
transform -1 0 34868 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1688980957
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1688980957
transform -1 0 34868 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1688980957
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1688980957
transform -1 0 34868 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1688980957
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1688980957
transform -1 0 34868 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1688980957
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1688980957
transform -1 0 34868 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1688980957
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1688980957
transform -1 0 34868 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1688980957
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1688980957
transform -1 0 34868 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1688980957
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1688980957
transform -1 0 34868 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1688980957
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1688980957
transform -1 0 34868 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1688980957
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1688980957
transform -1 0 34868 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1688980957
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1688980957
transform -1 0 34868 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1688980957
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1688980957
transform -1 0 34868 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1688980957
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1688980957
transform -1 0 34868 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1688980957
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1688980957
transform -1 0 34868 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1688980957
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1688980957
transform -1 0 34868 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1688980957
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1688980957
transform -1 0 34868 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1688980957
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1688980957
transform -1 0 34868 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1688980957
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1688980957
transform -1 0 34868 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1688980957
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1688980957
transform -1 0 34868 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1688980957
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1688980957
transform -1 0 34868 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1688980957
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1688980957
transform -1 0 34868 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1688980957
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1688980957
transform -1 0 34868 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1688980957
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1688980957
transform -1 0 34868 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1688980957
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1688980957
transform -1 0 34868 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1688980957
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1688980957
transform -1 0 34868 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1688980957
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1688980957
transform -1 0 34868 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1688980957
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1688980957
transform -1 0 34868 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1688980957
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1688980957
transform -1 0 34868 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1688980957
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1688980957
transform -1 0 34868 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1688980957
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1688980957
transform -1 0 34868 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1688980957
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1688980957
transform -1 0 34868 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1688980957
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1688980957
transform -1 0 34868 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1688980957
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1688980957
transform -1 0 34868 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1688980957
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1688980957
transform -1 0 34868 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1688980957
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1688980957
transform -1 0 34868 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1688980957
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1688980957
transform -1 0 34868 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1688980957
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1688980957
transform -1 0 34868 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1688980957
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1688980957
transform -1 0 34868 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1688980957
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1688980957
transform -1 0 34868 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1688980957
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1688980957
transform -1 0 34868 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1688980957
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1688980957
transform -1 0 34868 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1688980957
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1688980957
transform -1 0 34868 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1688980957
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1688980957
transform -1 0 34868 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1688980957
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1688980957
transform -1 0 34868 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1688980957
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1688980957
transform -1 0 34868 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1688980957
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1688980957
transform -1 0 34868 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1688980957
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1688980957
transform -1 0 34868 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1688980957
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1688980957
transform -1 0 34868 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1688980957
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1688980957
transform -1 0 34868 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1688980957
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1688980957
transform -1 0 34868 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1688980957
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1688980957
transform -1 0 34868 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1688980957
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1688980957
transform -1 0 34868 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1688980957
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1688980957
transform -1 0 34868 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1688980957
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1688980957
transform -1 0 34868 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1688980957
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1688980957
transform -1 0 34868 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1688980957
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1688980957
transform -1 0 34868 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1688980957
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1688980957
transform -1 0 34868 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1688980957
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1688980957
transform -1 0 34868 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1688980957
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1688980957
transform -1 0 34868 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1688980957
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1688980957
transform -1 0 34868 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1688980957
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1688980957
transform -1 0 34868 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1688980957
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1688980957
transform -1 0 34868 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1688980957
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1688980957
transform -1 0 34868 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1688980957
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1688980957
transform -1 0 34868 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1688980957
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1688980957
transform -1 0 34868 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1688980957
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1688980957
transform -1 0 34868 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1688980957
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1688980957
transform -1 0 34868 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1688980957
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1688980957
transform -1 0 34868 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rgb_mixer_13
timestamp 1688980957
transform -1 0 13892 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rgb_mixer_14
timestamp 1688980957
transform -1 0 1656 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rgb_mixer_15
timestamp 1688980957
transform 1 0 34316 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rgb_mixer_16
timestamp 1688980957
transform -1 0 1656 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rgb_mixer_17
timestamp 1688980957
transform -1 0 34592 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rgb_mixer_18
timestamp 1688980957
transform 1 0 27140 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rgb_mixer_19
timestamp 1688980957
transform 1 0 1380 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rgb_mixer_20
timestamp 1688980957
transform -1 0 34592 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rgb_mixer_21
timestamp 1688980957
transform 1 0 6532 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rgb_mixer_22
timestamp 1688980957
transform 1 0 34224 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1688980957
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1688980957
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1688980957
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1688980957
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1688980957
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1688980957
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1688980957
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1688980957
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1688980957
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1688980957
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1688980957
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1688980957
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1688980957
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1688980957
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1688980957
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1688980957
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1688980957
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1688980957
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1688980957
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1688980957
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1688980957
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1688980957
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1688980957
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1688980957
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1688980957
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1688980957
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1688980957
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1688980957
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1688980957
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1688980957
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1688980957
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1688980957
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1688980957
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1688980957
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1688980957
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1688980957
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1688980957
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1688980957
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1688980957
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1688980957
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1688980957
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1688980957
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1688980957
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1688980957
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1688980957
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1688980957
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1688980957
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1688980957
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1688980957
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1688980957
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1688980957
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1688980957
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1688980957
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1688980957
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1688980957
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1688980957
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1688980957
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1688980957
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1688980957
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1688980957
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1688980957
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1688980957
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1688980957
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1688980957
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1688980957
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1688980957
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1688980957
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1688980957
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1688980957
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1688980957
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1688980957
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1688980957
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1688980957
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1688980957
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1688980957
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1688980957
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1688980957
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1688980957
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1688980957
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1688980957
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1688980957
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1688980957
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1688980957
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1688980957
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1688980957
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1688980957
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1688980957
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1688980957
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1688980957
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1688980957
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1688980957
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1688980957
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1688980957
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1688980957
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1688980957
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1688980957
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1688980957
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1688980957
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1688980957
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1688980957
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1688980957
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1688980957
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1688980957
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1688980957
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1688980957
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1688980957
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1688980957
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1688980957
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1688980957
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1688980957
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1688980957
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1688980957
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1688980957
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1688980957
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1688980957
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1688980957
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1688980957
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1688980957
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1688980957
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1688980957
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1688980957
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1688980957
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1688980957
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1688980957
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1688980957
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1688980957
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1688980957
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1688980957
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1688980957
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1688980957
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1688980957
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1688980957
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1688980957
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1688980957
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1688980957
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1688980957
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1688980957
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1688980957
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1688980957
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1688980957
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1688980957
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1688980957
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1688980957
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1688980957
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1688980957
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1688980957
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1688980957
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1688980957
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1688980957
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1688980957
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1688980957
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1688980957
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1688980957
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1688980957
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1688980957
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1688980957
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1688980957
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1688980957
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1688980957
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1688980957
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1688980957
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1688980957
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1688980957
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1688980957
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1688980957
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1688980957
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1688980957
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1688980957
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1688980957
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1688980957
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1688980957
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1688980957
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1688980957
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1688980957
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1688980957
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1688980957
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1688980957
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1688980957
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1688980957
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1688980957
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1688980957
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1688980957
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1688980957
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1688980957
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1688980957
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1688980957
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1688980957
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1688980957
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1688980957
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1688980957
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1688980957
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1688980957
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1688980957
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1688980957
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1688980957
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1688980957
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1688980957
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1688980957
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1688980957
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1688980957
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1688980957
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1688980957
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1688980957
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1688980957
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1688980957
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1688980957
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1688980957
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1688980957
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1688980957
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1688980957
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1688980957
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1688980957
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1688980957
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1688980957
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1688980957
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1688980957
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1688980957
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1688980957
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1688980957
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1688980957
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1688980957
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1688980957
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1688980957
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1688980957
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1688980957
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1688980957
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1688980957
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1688980957
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1688980957
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1688980957
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1688980957
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1688980957
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1688980957
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1688980957
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1688980957
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1688980957
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1688980957
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1688980957
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1688980957
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1688980957
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1688980957
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1688980957
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1688980957
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1688980957
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1688980957
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1688980957
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1688980957
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1688980957
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1688980957
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1688980957
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1688980957
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1688980957
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1688980957
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1688980957
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1688980957
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1688980957
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1688980957
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1688980957
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1688980957
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1688980957
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1688980957
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1688980957
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1688980957
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1688980957
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1688980957
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1688980957
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1688980957
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1688980957
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1688980957
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1688980957
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1688980957
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1688980957
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1688980957
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1688980957
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1688980957
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1688980957
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1688980957
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1688980957
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1688980957
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1688980957
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1688980957
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1688980957
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1688980957
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1688980957
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1688980957
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1688980957
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1688980957
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1688980957
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1688980957
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1688980957
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1688980957
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1688980957
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1688980957
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1688980957
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1688980957
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1688980957
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1688980957
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1688980957
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1688980957
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1688980957
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1688980957
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1688980957
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1688980957
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1688980957
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1688980957
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1688980957
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1688980957
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1688980957
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1688980957
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1688980957
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1688980957
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1688980957
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1688980957
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1688980957
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1688980957
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1688980957
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1688980957
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1688980957
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1688980957
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1688980957
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1688980957
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1688980957
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1688980957
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1688980957
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1688980957
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1688980957
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1688980957
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1688980957
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1688980957
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1688980957
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1688980957
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1688980957
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1688980957
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1688980957
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1688980957
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1688980957
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1688980957
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1688980957
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1688980957
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1688980957
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1688980957
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1688980957
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1688980957
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1688980957
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1688980957
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1688980957
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1688980957
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1688980957
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1688980957
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1688980957
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1688980957
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1688980957
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1688980957
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1688980957
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1688980957
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1688980957
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1688980957
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1688980957
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1688980957
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1688980957
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1688980957
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1688980957
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1688980957
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1688980957
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1688980957
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1688980957
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1688980957
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1688980957
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1688980957
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1688980957
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1688980957
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1688980957
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1688980957
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1688980957
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1688980957
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1688980957
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1688980957
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1688980957
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1688980957
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1688980957
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1688980957
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1688980957
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1688980957
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1688980957
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1688980957
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1688980957
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1688980957
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1688980957
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1688980957
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1688980957
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1688980957
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1688980957
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1688980957
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1688980957
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1688980957
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1688980957
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1688980957
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1688980957
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1688980957
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1688980957
transform 1 0 26864 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1688980957
transform 1 0 32016 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1688980957
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1688980957
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1688980957
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1688980957
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1688980957
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1688980957
transform 1 0 29440 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1688980957
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1688980957
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1688980957
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1688980957
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1688980957
transform 1 0 26864 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1688980957
transform 1 0 32016 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1688980957
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1688980957
transform 1 0 6256 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1688980957
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1688980957
transform 1 0 11408 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1688980957
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1688980957
transform 1 0 16560 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1688980957
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1688980957
transform 1 0 21712 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1688980957
transform 1 0 24288 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1688980957
transform 1 0 26864 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1688980957
transform 1 0 29440 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1688980957
transform 1 0 32016 0 1 39168
box -38 -48 130 592
<< labels >>
flabel metal2 s 28970 41200 29082 42000 0 FreeSans 448 90 0 0 clk
port 0 nsew signal input
flabel metal2 s 14802 41200 14914 42000 0 FreeSans 448 90 0 0 enc0_a
port 1 nsew signal input
flabel metal3 s 35200 34628 36000 34868 0 FreeSans 960 0 0 0 enc0_b
port 2 nsew signal input
flabel metal3 s 35200 12868 36000 13108 0 FreeSans 960 0 0 0 enc1_a
port 3 nsew signal input
flabel metal2 s 8362 41200 8474 42000 0 FreeSans 448 90 0 0 enc1_b
port 4 nsew signal input
flabel metal3 s 0 28508 800 28748 0 FreeSans 960 0 0 0 enc2_a
port 5 nsew signal input
flabel metal3 s 0 14228 800 14468 0 FreeSans 960 0 0 0 enc2_b
port 6 nsew signal input
flabel metal3 s 35200 5388 36000 5628 0 FreeSans 960 0 0 0 io_oeb_high[0]
port 7 nsew signal tristate
flabel metal2 s 27038 0 27150 800 0 FreeSans 448 90 0 0 io_oeb_high[1]
port 8 nsew signal tristate
flabel metal2 s -10 0 102 800 0 FreeSans 448 90 0 0 io_oeb_high[2]
port 9 nsew signal tristate
flabel metal2 s 35410 41200 35522 42000 0 FreeSans 448 90 0 0 io_oeb_high[3]
port 10 nsew signal tristate
flabel metal2 s 6430 0 6542 800 0 FreeSans 448 90 0 0 io_oeb_high[4]
port 11 nsew signal tristate
flabel metal2 s 34122 0 34234 800 0 FreeSans 448 90 0 0 io_oeb_high[5]
port 12 nsew signal tristate
flabel metal2 s 13514 0 13626 800 0 FreeSans 448 90 0 0 io_oeb_low[0]
port 13 nsew signal tristate
flabel metal3 s 0 6748 800 6988 0 FreeSans 960 0 0 0 io_oeb_low[1]
port 14 nsew signal tristate
flabel metal3 s 35200 27148 36000 27388 0 FreeSans 960 0 0 0 io_oeb_low[2]
port 15 nsew signal tristate
flabel metal3 s 0 35988 800 36228 0 FreeSans 960 0 0 0 io_oeb_low[3]
port 16 nsew signal tristate
flabel metal2 s 21886 41200 21998 42000 0 FreeSans 448 90 0 0 pwm0_out
port 17 nsew signal tristate
flabel metal2 s 20598 0 20710 800 0 FreeSans 448 90 0 0 pwm1_out
port 18 nsew signal tristate
flabel metal3 s 0 21708 800 21948 0 FreeSans 960 0 0 0 pwm2_out
port 19 nsew signal tristate
flabel metal2 s 1278 41200 1390 42000 0 FreeSans 448 90 0 0 reset
port 20 nsew signal input
flabel metal3 s 35200 19668 36000 19908 0 FreeSans 960 0 0 0 sync
port 21 nsew signal tristate
flabel metal4 s 5164 2128 5484 39760 0 FreeSans 1920 90 0 0 vccd1
port 22 nsew power bidirectional
flabel metal4 s 13605 2128 13925 39760 0 FreeSans 1920 90 0 0 vccd1
port 22 nsew power bidirectional
flabel metal4 s 22046 2128 22366 39760 0 FreeSans 1920 90 0 0 vccd1
port 22 nsew power bidirectional
flabel metal4 s 30487 2128 30807 39760 0 FreeSans 1920 90 0 0 vccd1
port 22 nsew power bidirectional
flabel metal4 s 9384 2128 9704 39760 0 FreeSans 1920 90 0 0 vssd1
port 23 nsew ground bidirectional
flabel metal4 s 17825 2128 18145 39760 0 FreeSans 1920 90 0 0 vssd1
port 23 nsew ground bidirectional
flabel metal4 s 26266 2128 26586 39760 0 FreeSans 1920 90 0 0 vssd1
port 23 nsew ground bidirectional
flabel metal4 s 34707 2128 35027 39760 0 FreeSans 1920 90 0 0 vssd1
port 23 nsew ground bidirectional
rlabel metal1 17986 39712 17986 39712 0 vccd1
rlabel via1 18065 39168 18065 39168 0 vssd1
rlabel metal1 8280 36346 8280 36346 0 _000_
rlabel metal1 16376 36346 16376 36346 0 _001_
rlabel metal1 14209 38998 14209 38998 0 _002_
rlabel metal1 14198 38250 14198 38250 0 _003_
rlabel metal1 14842 37910 14842 37910 0 _004_
rlabel metal1 15946 38250 15946 38250 0 _005_
rlabel metal1 17234 38998 17234 38998 0 _006_
rlabel metal1 17884 35666 17884 35666 0 _007_
rlabel metal2 19090 36754 19090 36754 0 _008_
rlabel metal1 16514 36890 16514 36890 0 _009_
rlabel metal1 20562 35666 20562 35666 0 _010_
rlabel metal1 24426 35802 24426 35802 0 _011_
rlabel metal2 20746 38114 20746 38114 0 _012_
rlabel metal1 20511 38998 20511 38998 0 _013_
rlabel metal1 21482 39032 21482 39032 0 _014_
rlabel metal2 23046 36958 23046 36958 0 _015_
rlabel metal1 19775 35734 19775 35734 0 _016_
rlabel metal2 21390 35938 21390 35938 0 _017_
rlabel metal2 23874 35938 23874 35938 0 _018_
rlabel metal1 22264 32334 22264 32334 0 _019_
rlabel metal2 23874 30022 23874 30022 0 _020_
rlabel metal2 23874 31552 23874 31552 0 _021_
rlabel metal1 24375 32470 24375 32470 0 _022_
rlabel metal1 24564 33626 24564 33626 0 _023_
rlabel metal1 23889 33558 23889 33558 0 _024_
rlabel metal1 22356 33082 22356 33082 0 _025_
rlabel via1 22765 33898 22765 33898 0 _026_
rlabel metal1 21758 31994 21758 31994 0 _027_
rlabel metal1 13386 35802 13386 35802 0 _028_
rlabel via1 9057 36822 9057 36822 0 _029_
rlabel metal1 9420 35666 9420 35666 0 _030_
rlabel metal1 9839 35054 9839 35054 0 _031_
rlabel metal1 10023 37162 10023 37162 0 _032_
rlabel metal1 11449 37162 11449 37162 0 _033_
rlabel viali 12267 34578 12267 34578 0 _034_
rlabel metal1 13769 34986 13769 34986 0 _035_
rlabel metal1 12875 37162 12875 37162 0 _036_
rlabel metal1 9108 32470 9108 32470 0 _037_
rlabel metal1 6762 30124 6762 30124 0 _038_
rlabel metal2 8050 31586 8050 31586 0 _039_
rlabel via1 9241 31790 9241 31790 0 _040_
rlabel metal1 7999 33558 7999 33558 0 _041_
rlabel via1 9241 32878 9241 32878 0 _042_
rlabel metal1 11009 33558 11009 33558 0 _043_
rlabel via1 12654 33490 12654 33490 0 _044_
rlabel metal1 12539 32402 12539 32402 0 _045_
rlabel metal2 12558 30906 12558 30906 0 _046_
rlabel metal1 16836 20026 16836 20026 0 _047_
rlabel metal1 15226 21386 15226 21386 0 _048_
rlabel metal1 14352 19482 14352 19482 0 _049_
rlabel metal1 13202 20026 13202 20026 0 _050_
rlabel metal1 12236 20434 12236 20434 0 _051_
rlabel metal1 11178 19312 11178 19312 0 _052_
rlabel metal1 8648 20978 8648 20978 0 _053_
rlabel metal1 9752 21454 9752 21454 0 _054_
rlabel metal2 15042 34850 15042 34850 0 _055_
rlabel metal1 6624 28730 6624 28730 0 _056_
rlabel metal1 7815 29614 7815 29614 0 _057_
rlabel metal1 7436 27370 7436 27370 0 _058_
rlabel metal1 7666 28118 7666 28118 0 _059_
rlabel metal1 9655 27370 9655 27370 0 _060_
rlabel metal1 10212 29818 10212 29818 0 _061_
rlabel metal1 9977 30294 9977 30294 0 _062_
rlabel metal1 10058 28118 10058 28118 0 _063_
rlabel metal1 14030 31450 14030 31450 0 _064_
rlabel metal2 13386 32980 13386 32980 0 _065_
rlabel metal1 15686 33626 15686 33626 0 _066_
rlabel metal1 14996 30362 14996 30362 0 _067_
rlabel metal2 17710 34612 17710 34612 0 _068_
rlabel metal1 18400 31246 18400 31246 0 _069_
rlabel metal1 19182 33456 19182 33456 0 _070_
rlabel metal1 20332 31790 20332 31790 0 _071_
rlabel metal1 21850 29580 21850 29580 0 _072_
rlabel metal2 16054 35190 16054 35190 0 _073_
rlabel metal1 21068 24174 21068 24174 0 _074_
rlabel metal1 20700 27506 20700 27506 0 _075_
rlabel metal1 23230 27098 23230 27098 0 _076_
rlabel metal1 23552 24718 23552 24718 0 _077_
rlabel metal1 23138 23834 23138 23834 0 _078_
rlabel metal1 22862 22746 22862 22746 0 _079_
rlabel metal1 20005 19754 20005 19754 0 _080_
rlabel metal1 22402 20434 22402 20434 0 _081_
rlabel metal2 14122 30430 14122 30430 0 _082_
rlabel metal1 21942 29104 21942 29104 0 _083_
rlabel metal1 14904 23086 14904 23086 0 _084_
rlabel metal1 16974 23834 16974 23834 0 _085_
rlabel metal1 15686 25670 15686 25670 0 _086_
rlabel metal1 13156 23834 13156 23834 0 _087_
rlabel metal1 12834 26554 12834 26554 0 _088_
rlabel metal2 11270 26044 11270 26044 0 _089_
rlabel metal1 9568 23834 9568 23834 0 _090_
rlabel metal2 12742 24004 12742 24004 0 _091_
rlabel metal1 11898 28458 11898 28458 0 _092_
rlabel metal1 14306 27506 14306 27506 0 _093_
rlabel metal1 14122 30124 14122 30124 0 _094_
rlabel metal1 16192 27982 16192 27982 0 _095_
rlabel via1 17162 27438 17162 27438 0 _096_
rlabel metal2 16790 28730 16790 28730 0 _097_
rlabel metal2 20378 28492 20378 28492 0 _098_
rlabel metal1 18814 28594 18814 28594 0 _099_
rlabel metal1 20332 28730 20332 28730 0 _100_
rlabel metal1 15640 25806 15640 25806 0 _101_
rlabel metal1 15962 25738 15962 25738 0 _102_
rlabel metal2 17158 26724 17158 26724 0 _103_
rlabel metal1 18430 23766 18430 23766 0 _104_
rlabel metal1 17342 23154 17342 23154 0 _105_
rlabel metal1 16767 22066 16767 22066 0 _106_
rlabel metal1 18538 22610 18538 22610 0 _107_
rlabel metal2 18446 19618 18446 19618 0 _108_
rlabel metal1 20424 30702 20424 30702 0 _109_
rlabel metal1 19642 30158 19642 30158 0 _110_
rlabel metal1 20194 30634 20194 30634 0 _111_
rlabel metal1 19182 30260 19182 30260 0 _112_
rlabel metal1 17480 30226 17480 30226 0 _113_
rlabel metal1 17250 30158 17250 30158 0 _114_
rlabel metal1 15962 29580 15962 29580 0 _115_
rlabel metal1 17664 31994 17664 31994 0 _116_
rlabel via1 14030 30141 14030 30141 0 _117_
rlabel metal1 15732 29614 15732 29614 0 _118_
rlabel metal2 14582 31042 14582 31042 0 _119_
rlabel metal1 15456 29614 15456 29614 0 _120_
rlabel metal1 16422 29818 16422 29818 0 _121_
rlabel metal1 17204 31926 17204 31926 0 _122_
rlabel metal1 17894 30226 17894 30226 0 _123_
rlabel metal1 18998 30192 18998 30192 0 _124_
rlabel metal1 20010 30362 20010 30362 0 _125_
rlabel metal1 17388 20842 17388 20842 0 _126_
rlabel metal1 11638 34544 11638 34544 0 _127_
rlabel metal1 19780 33898 19780 33898 0 _128_
rlabel metal1 15686 23698 15686 23698 0 _129_
rlabel metal1 20470 21488 20470 21488 0 _130_
rlabel metal1 20194 21420 20194 21420 0 _131_
rlabel via1 20285 21998 20285 21998 0 _132_
rlabel metal1 20194 22950 20194 22950 0 _133_
rlabel metal1 19642 24854 19642 24854 0 _134_
rlabel metal1 19964 23766 19964 23766 0 _135_
rlabel metal1 19752 25262 19752 25262 0 _136_
rlabel metal1 20654 25806 20654 25806 0 _137_
rlabel metal1 19550 26384 19550 26384 0 _138_
rlabel metal1 20424 25874 20424 25874 0 _139_
rlabel metal1 20056 25874 20056 25874 0 _140_
rlabel metal1 20010 25262 20010 25262 0 _141_
rlabel metal1 20240 23698 20240 23698 0 _142_
rlabel metal1 19458 22644 19458 22644 0 _143_
rlabel metal1 20286 22406 20286 22406 0 _144_
rlabel metal1 19826 21862 19826 21862 0 _145_
rlabel metal1 20615 20978 20615 20978 0 _146_
rlabel metal2 14582 19856 14582 19856 0 _147_
rlabel metal1 10810 22032 10810 22032 0 _148_
rlabel metal1 10810 21454 10810 21454 0 _149_
rlabel metal1 11868 21998 11868 21998 0 _150_
rlabel metal1 12512 21522 12512 21522 0 _151_
rlabel metal1 13202 22032 13202 22032 0 _152_
rlabel metal1 12926 21590 12926 21590 0 _153_
rlabel via1 14673 21998 14673 21998 0 _154_
rlabel metal1 14444 20978 14444 20978 0 _155_
rlabel metal2 15134 21828 15134 21828 0 _156_
rlabel metal1 14720 21114 14720 21114 0 _157_
rlabel metal1 15134 20910 15134 20910 0 _158_
rlabel metal1 14950 21114 14950 21114 0 _159_
rlabel metal1 13110 21522 13110 21522 0 _160_
rlabel metal1 12558 21658 12558 21658 0 _161_
rlabel metal1 12190 21556 12190 21556 0 _162_
rlabel metal1 11362 21522 11362 21522 0 _163_
rlabel metal1 10718 21658 10718 21658 0 _164_
rlabel metal2 17342 38352 17342 38352 0 _165_
rlabel metal1 17158 36176 17158 36176 0 _166_
rlabel metal1 18124 37434 18124 37434 0 _167_
rlabel metal2 17250 36890 17250 36890 0 _168_
rlabel metal1 18584 33966 18584 33966 0 _169_
rlabel metal2 15594 32300 15594 32300 0 _170_
rlabel metal1 13892 38930 13892 38930 0 _171_
rlabel metal1 13754 38420 13754 38420 0 _172_
rlabel metal1 14766 37434 14766 37434 0 _173_
rlabel metal1 16146 38930 16146 38930 0 _174_
rlabel metal1 18630 39338 18630 39338 0 _175_
rlabel metal1 16882 39440 16882 39440 0 _176_
rlabel metal1 17066 35666 17066 35666 0 _177_
rlabel metal1 18906 36108 18906 36108 0 _178_
rlabel metal1 16008 36754 16008 36754 0 _179_
rlabel metal2 21206 37536 21206 37536 0 _180_
rlabel metal2 21850 35904 21850 35904 0 _181_
rlabel metal2 22402 36380 22402 36380 0 _182_
rlabel metal1 21344 35258 21344 35258 0 _183_
rlabel metal1 24012 35258 24012 35258 0 _184_
rlabel metal1 20792 37842 20792 37842 0 _185_
rlabel metal1 20746 39372 20746 39372 0 _186_
rlabel metal1 21298 39474 21298 39474 0 _187_
rlabel metal1 22816 37230 22816 37230 0 _188_
rlabel metal1 20746 36754 20746 36754 0 _189_
rlabel metal1 21344 35666 21344 35666 0 _190_
rlabel metal1 22034 32844 22034 32844 0 _191_
rlabel metal1 23920 35666 23920 35666 0 _192_
rlabel metal1 23552 31926 23552 31926 0 _193_
rlabel metal2 22954 32198 22954 32198 0 _194_
rlabel metal2 23966 31892 23966 31892 0 _195_
rlabel metal1 23046 32436 23046 32436 0 _196_
rlabel metal1 24104 29274 24104 29274 0 _197_
rlabel metal1 24150 30906 24150 30906 0 _198_
rlabel metal1 24610 32912 24610 32912 0 _199_
rlabel metal1 24656 33490 24656 33490 0 _200_
rlabel metal1 24288 33966 24288 33966 0 _201_
rlabel metal2 22494 33762 22494 33762 0 _202_
rlabel metal1 22402 33014 22402 33014 0 _203_
rlabel metal1 21482 31790 21482 31790 0 _204_
rlabel metal1 13156 36210 13156 36210 0 _205_
rlabel metal1 12926 35700 12926 35700 0 _206_
rlabel metal2 12558 36516 12558 36516 0 _207_
rlabel metal1 12834 35734 12834 35734 0 _208_
rlabel metal1 8786 37842 8786 37842 0 _209_
rlabel metal1 9844 35258 9844 35258 0 _210_
rlabel metal1 10212 36142 10212 36142 0 _211_
rlabel metal1 12558 36074 12558 36074 0 _212_
rlabel metal1 10396 37842 10396 37842 0 _213_
rlabel metal1 12052 36278 12052 36278 0 _214_
rlabel metal1 11178 35700 11178 35700 0 _215_
rlabel metal1 14306 35156 14306 35156 0 _216_
rlabel metal1 14076 37434 14076 37434 0 _217_
rlabel metal2 10902 33116 10902 33116 0 _218_
rlabel metal1 9430 32368 9430 32368 0 _219_
rlabel metal1 9338 32266 9338 32266 0 _220_
rlabel metal1 9522 32436 9522 32436 0 _221_
rlabel metal1 6440 29818 6440 29818 0 _222_
rlabel metal1 8280 31314 8280 31314 0 _223_
rlabel metal1 7958 32470 7958 32470 0 _224_
rlabel metal1 8280 33082 8280 33082 0 _225_
rlabel metal1 8786 33966 8786 33966 0 _226_
rlabel metal1 11316 33490 11316 33490 0 _227_
rlabel metal1 9384 30226 9384 30226 0 _228_
rlabel metal2 11362 34884 11362 34884 0 _229_
rlabel metal1 11362 32912 11362 32912 0 _230_
rlabel metal1 8326 28696 8326 28696 0 _231_
rlabel metal1 11362 29206 11362 29206 0 _232_
rlabel metal1 10074 28526 10074 28526 0 _233_
rlabel metal1 11224 28730 11224 28730 0 _234_
rlabel metal2 21712 21522 21712 21522 0 _235_
rlabel metal1 14720 21862 14720 21862 0 _236_
rlabel metal2 13248 21522 13248 21522 0 _237_
rlabel metal1 14398 19346 14398 19346 0 _238_
rlabel metal1 12880 21114 12880 21114 0 _239_
rlabel metal2 13340 21420 13340 21420 0 _240_
rlabel metal1 18722 20944 18722 20944 0 _241_
rlabel metal1 13524 21114 13524 21114 0 _242_
rlabel metal1 12466 20978 12466 20978 0 _243_
rlabel metal1 10258 19822 10258 19822 0 _244_
rlabel metal1 9936 20026 9936 20026 0 _245_
rlabel metal1 9154 21318 9154 21318 0 _246_
rlabel metal1 8832 20570 8832 20570 0 _247_
rlabel metal1 9568 21522 9568 21522 0 _248_
rlabel metal1 14996 34578 14996 34578 0 _249_
rlabel metal1 6302 28526 6302 28526 0 _250_
rlabel metal1 8096 29274 8096 29274 0 _251_
rlabel metal1 7130 28050 7130 28050 0 _252_
rlabel metal1 7406 28050 7406 28050 0 _253_
rlabel metal1 9752 27098 9752 27098 0 _254_
rlabel metal1 10580 29614 10580 29614 0 _255_
rlabel metal1 9660 30294 9660 30294 0 _256_
rlabel metal2 11546 28322 11546 28322 0 _257_
rlabel metal1 17848 35122 17848 35122 0 _258_
rlabel metal1 17940 35190 17940 35190 0 _259_
rlabel metal1 16790 35088 16790 35088 0 _260_
rlabel metal1 16882 34986 16882 34986 0 _261_
rlabel metal1 15364 32334 15364 32334 0 _262_
rlabel metal1 19872 31790 19872 31790 0 _263_
rlabel metal2 14398 31756 14398 31756 0 _264_
rlabel metal1 16376 32878 16376 32878 0 _265_
rlabel metal1 13938 34170 13938 34170 0 _266_
rlabel metal1 14214 32878 14214 32878 0 _267_
rlabel metal1 14536 32198 14536 32198 0 _268_
rlabel metal1 13432 34102 13432 34102 0 _269_
rlabel metal1 13846 32436 13846 32436 0 _270_
rlabel metal1 15548 32878 15548 32878 0 _271_
rlabel metal2 16146 33286 16146 33286 0 _272_
rlabel metal1 16330 32742 16330 32742 0 _273_
rlabel metal1 16008 33490 16008 33490 0 _274_
rlabel metal1 15870 33354 15870 33354 0 _275_
rlabel metal1 14904 33082 14904 33082 0 _276_
rlabel metal1 15042 33456 15042 33456 0 _277_
rlabel metal1 16468 32334 16468 32334 0 _278_
rlabel metal2 15594 32844 15594 32844 0 _279_
rlabel metal1 16928 32402 16928 32402 0 _280_
rlabel metal1 17020 32198 17020 32198 0 _281_
rlabel metal1 16238 32436 16238 32436 0 _282_
rlabel metal1 16652 33490 16652 33490 0 _283_
rlabel metal1 17894 32844 17894 32844 0 _284_
rlabel metal1 18676 33082 18676 33082 0 _285_
rlabel metal1 17434 33286 17434 33286 0 _286_
rlabel metal1 18032 33626 18032 33626 0 _287_
rlabel metal1 17802 32402 17802 32402 0 _288_
rlabel metal1 17710 31824 17710 31824 0 _289_
rlabel metal1 17802 31348 17802 31348 0 _290_
rlabel metal2 17618 31969 17618 31969 0 _291_
rlabel metal1 19274 33388 19274 33388 0 _292_
rlabel metal1 21114 32810 21114 32810 0 _293_
rlabel metal1 19964 32742 19964 32742 0 _294_
rlabel metal1 20654 33456 20654 33456 0 _295_
rlabel metal2 19182 32351 19182 32351 0 _296_
rlabel metal2 20194 33388 20194 33388 0 _297_
rlabel metal1 20516 33082 20516 33082 0 _298_
rlabel metal1 19458 33456 19458 33456 0 _299_
rlabel metal1 19699 33558 19699 33558 0 _300_
rlabel metal1 18998 33558 18998 33558 0 _301_
rlabel metal1 20148 32538 20148 32538 0 _302_
rlabel metal2 19734 31892 19734 31892 0 _303_
rlabel metal1 19642 31858 19642 31858 0 _304_
rlabel metal2 21666 30022 21666 30022 0 _305_
rlabel metal1 16238 34646 16238 34646 0 _306_
rlabel metal1 22770 28526 22770 28526 0 _307_
rlabel metal2 22770 29104 22770 29104 0 _308_
rlabel metal1 23184 28730 23184 28730 0 _309_
rlabel metal1 23782 28526 23782 28526 0 _310_
rlabel metal1 23920 25806 23920 25806 0 _311_
rlabel metal1 21896 21318 21896 21318 0 _312_
rlabel metal2 21298 24786 21298 24786 0 _313_
rlabel metal2 21758 25840 21758 25840 0 _314_
rlabel metal1 21574 27846 21574 27846 0 _315_
rlabel viali 21391 26984 21391 26984 0 _316_
rlabel metal1 20470 26418 20470 26418 0 _317_
rlabel metal1 20838 26554 20838 26554 0 _318_
rlabel metal2 20746 26928 20746 26928 0 _319_
rlabel viali 22109 26962 22109 26962 0 _320_
rlabel metal1 23322 26316 23322 26316 0 _321_
rlabel metal2 21942 21216 21942 21216 0 _322_
rlabel metal1 23046 26418 23046 26418 0 _323_
rlabel metal1 22586 26554 22586 26554 0 _324_
rlabel metal1 22540 27098 22540 27098 0 _325_
rlabel metal1 22678 26996 22678 26996 0 _326_
rlabel metal1 23644 26010 23644 26010 0 _327_
rlabel metal2 23138 26044 23138 26044 0 _328_
rlabel metal1 22862 25908 22862 25908 0 _329_
rlabel metal1 22862 24820 22862 24820 0 _330_
rlabel metal1 21970 25874 21970 25874 0 _331_
rlabel metal1 21850 23018 21850 23018 0 _332_
rlabel metal1 21804 22746 21804 22746 0 _333_
rlabel metal1 22816 23086 22816 23086 0 _334_
rlabel metal2 21942 23375 21942 23375 0 _335_
rlabel metal1 22632 24174 22632 24174 0 _336_
rlabel metal1 22011 23562 22011 23562 0 _337_
rlabel metal1 22586 23732 22586 23732 0 _338_
rlabel metal2 22494 23460 22494 23460 0 _339_
rlabel metal1 22218 22678 22218 22678 0 _340_
rlabel metal1 22310 22678 22310 22678 0 _341_
rlabel metal1 22494 19890 22494 19890 0 _342_
rlabel metal1 22770 19754 22770 19754 0 _343_
rlabel metal2 22678 20774 22678 20774 0 _344_
rlabel metal1 22678 22202 22678 22202 0 _345_
rlabel metal1 22494 21556 22494 21556 0 _346_
rlabel metal1 22540 21658 22540 21658 0 _347_
rlabel metal1 20976 20026 20976 20026 0 _348_
rlabel metal1 21344 21522 21344 21522 0 _349_
rlabel metal1 22954 20298 22954 20298 0 _350_
rlabel metal2 21758 20468 21758 20468 0 _351_
rlabel metal2 23598 20638 23598 20638 0 _352_
rlabel metal1 13892 30702 13892 30702 0 _353_
rlabel metal1 21160 29138 21160 29138 0 _354_
rlabel metal2 12742 28492 12742 28492 0 _355_
rlabel metal1 13018 28118 13018 28118 0 _356_
rlabel metal1 12880 27982 12880 27982 0 _357_
rlabel metal1 13524 28186 13524 28186 0 _358_
rlabel metal2 14306 27370 14306 27370 0 _359_
rlabel metal1 13110 26282 13110 26282 0 _360_
rlabel metal2 14674 23290 14674 23290 0 _361_
rlabel metal2 13570 26163 13570 26163 0 _362_
rlabel metal1 15134 24718 15134 24718 0 _363_
rlabel metal1 14904 24242 14904 24242 0 _364_
rlabel metal1 15088 24650 15088 24650 0 _365_
rlabel metal2 15686 24208 15686 24208 0 _366_
rlabel metal1 15962 23732 15962 23732 0 _367_
rlabel metal1 13524 24786 13524 24786 0 _368_
rlabel metal1 14720 25262 14720 25262 0 _369_
rlabel metal1 10074 24786 10074 24786 0 _370_
rlabel metal1 14628 24922 14628 24922 0 _371_
rlabel metal1 14628 25806 14628 25806 0 _372_
rlabel metal1 15502 25296 15502 25296 0 _373_
rlabel metal1 14950 25840 14950 25840 0 _374_
rlabel metal1 13616 24650 13616 24650 0 _375_
rlabel metal1 14490 24174 14490 24174 0 _376_
rlabel metal2 14306 24004 14306 24004 0 _377_
rlabel metal1 13294 23732 13294 23732 0 _378_
rlabel metal1 13938 24378 13938 24378 0 _379_
rlabel metal2 12466 25619 12466 25619 0 _380_
rlabel metal2 13386 26214 13386 26214 0 _381_
rlabel metal1 12466 26418 12466 26418 0 _382_
rlabel metal2 12558 27268 12558 27268 0 _383_
rlabel metal1 13064 25398 13064 25398 0 _384_
rlabel metal1 12604 26350 12604 26350 0 _385_
rlabel metal1 13248 26350 13248 26350 0 _386_
rlabel metal1 12650 25704 12650 25704 0 _387_
rlabel metal1 11822 26316 11822 26316 0 _388_
rlabel metal1 11684 26418 11684 26418 0 _389_
rlabel metal1 10534 24650 10534 24650 0 _390_
rlabel metal1 11960 25262 11960 25262 0 _391_
rlabel metal2 10994 24990 10994 24990 0 _392_
rlabel metal1 12834 25466 12834 25466 0 _393_
rlabel metal1 10580 25262 10580 25262 0 _394_
rlabel metal1 11776 25330 11776 25330 0 _395_
rlabel metal1 10350 24752 10350 24752 0 _396_
rlabel metal1 11132 24242 11132 24242 0 _397_
rlabel metal1 11822 24616 11822 24616 0 _398_
rlabel metal1 11684 23698 11684 23698 0 _399_
rlabel viali 11822 23699 11822 23699 0 _400_
rlabel metal1 11454 29274 11454 29274 0 _401_
rlabel metal1 14306 30226 14306 30226 0 _402_
rlabel metal1 16284 29138 16284 29138 0 _403_
rlabel metal1 16100 28050 16100 28050 0 _404_
rlabel metal1 16652 29274 16652 29274 0 _405_
rlabel metal1 17480 29274 17480 29274 0 _406_
rlabel metal1 17572 28934 17572 28934 0 _407_
rlabel metal1 16422 28730 16422 28730 0 _408_
rlabel metal1 19090 29274 19090 29274 0 _409_
rlabel metal1 18492 29138 18492 29138 0 _410_
rlabel metal1 20010 30192 20010 30192 0 _411_
rlabel metal1 18860 29138 18860 29138 0 _412_
rlabel metal1 20332 28526 20332 28526 0 _413_
rlabel metal1 15548 25942 15548 25942 0 _414_
rlabel metal2 18630 25670 18630 25670 0 _415_
rlabel metal1 17112 26350 17112 26350 0 _416_
rlabel metal2 18262 23885 18262 23885 0 _417_
rlabel metal1 18492 24378 18492 24378 0 _418_
rlabel metal1 19401 21862 19401 21862 0 _419_
rlabel metal1 17020 23086 17020 23086 0 _420_
rlabel metal1 17894 20944 17894 20944 0 _421_
rlabel metal1 17296 20774 17296 20774 0 _422_
rlabel metal1 18906 20910 18906 20910 0 _423_
rlabel metal1 17940 22610 17940 22610 0 _424_
rlabel metal1 18676 19346 18676 19346 0 _425_
rlabel metal1 22034 29648 22034 29648 0 clk
rlabel metal1 19688 20502 19688 20502 0 clknet_0_clk
rlabel metal1 13616 19890 13616 19890 0 clknet_3_0__leaf_clk
rlabel metal2 13938 28254 13938 28254 0 clknet_3_1__leaf_clk
rlabel metal1 22632 20910 22632 20910 0 clknet_3_2__leaf_clk
rlabel metal1 19642 29172 19642 29172 0 clknet_3_3__leaf_clk
rlabel metal2 7406 32640 7406 32640 0 clknet_3_4__leaf_clk
rlabel metal1 12926 33524 12926 33524 0 clknet_3_5__leaf_clk
rlabel metal1 20562 31314 20562 31314 0 clknet_3_6__leaf_clk
rlabel metal1 17158 38828 17158 38828 0 clknet_3_7__leaf_clk
rlabel metal1 18078 39610 18078 39610 0 debounce0_a.button_hist\[0\]
rlabel metal2 17802 37536 17802 37536 0 debounce0_a.button_hist\[1\]
rlabel metal1 16744 37706 16744 37706 0 debounce0_a.button_hist\[2\]
rlabel metal1 17940 38318 17940 38318 0 debounce0_a.button_hist\[3\]
rlabel metal1 18768 38386 18768 38386 0 debounce0_a.button_hist\[4\]
rlabel metal1 18906 35802 18906 35802 0 debounce0_a.button_hist\[5\]
rlabel metal1 18584 37230 18584 37230 0 debounce0_a.button_hist\[6\]
rlabel metal1 17848 37978 17848 37978 0 debounce0_a.button_hist\[7\]
rlabel metal1 17296 37230 17296 37230 0 debounce0_a.debounced
rlabel metal1 9154 36278 9154 36278 0 debounce0_a.reset
rlabel metal1 21873 37638 21873 37638 0 debounce0_b.button_hist\[0\]
rlabel metal1 21298 38420 21298 38420 0 debounce0_b.button_hist\[1\]
rlabel metal2 21666 38454 21666 38454 0 debounce0_b.button_hist\[2\]
rlabel metal1 21942 38318 21942 38318 0 debounce0_b.button_hist\[3\]
rlabel metal2 21942 37060 21942 37060 0 debounce0_b.button_hist\[4\]
rlabel metal2 20562 36244 20562 36244 0 debounce0_b.button_hist\[5\]
rlabel metal1 22264 35530 22264 35530 0 debounce0_b.button_hist\[6\]
rlabel metal1 22356 35666 22356 35666 0 debounce0_b.button_hist\[7\]
rlabel metal1 20102 35258 20102 35258 0 debounce0_b.debounced
rlabel metal1 24288 31994 24288 31994 0 debounce1_a.button_hist\[0\]
rlabel metal1 25300 31994 25300 31994 0 debounce1_a.button_hist\[1\]
rlabel metal1 25392 32538 25392 32538 0 debounce1_a.button_hist\[2\]
rlabel metal1 24426 34714 24426 34714 0 debounce1_a.button_hist\[3\]
rlabel metal1 22862 33626 22862 33626 0 debounce1_a.button_hist\[4\]
rlabel metal1 21436 33490 21436 33490 0 debounce1_a.button_hist\[5\]
rlabel metal1 23966 32878 23966 32878 0 debounce1_a.button_hist\[6\]
rlabel metal1 23598 31994 23598 31994 0 debounce1_a.button_hist\[7\]
rlabel metal2 21482 32096 21482 32096 0 debounce1_a.debounced
rlabel metal1 10856 36686 10856 36686 0 debounce1_b.button_hist\[0\]
rlabel metal1 11362 36210 11362 36210 0 debounce1_b.button_hist\[1\]
rlabel metal2 10810 37026 10810 37026 0 debounce1_b.button_hist\[2\]
rlabel metal1 11960 37774 11960 37774 0 debounce1_b.button_hist\[3\]
rlabel metal1 12466 36822 12466 36822 0 debounce1_b.button_hist\[4\]
rlabel metal2 13386 35156 13386 35156 0 debounce1_b.button_hist\[5\]
rlabel metal1 12696 36686 12696 36686 0 debounce1_b.button_hist\[6\]
rlabel metal1 13064 36890 13064 36890 0 debounce1_b.button_hist\[7\]
rlabel metal1 18492 32878 18492 32878 0 debounce1_b.debounced
rlabel metal2 8418 33218 8418 33218 0 debounce2_a.button_hist\[0\]
rlabel metal1 8832 31994 8832 31994 0 debounce2_a.button_hist\[1\]
rlabel metal1 8786 32810 8786 32810 0 debounce2_a.button_hist\[2\]
rlabel metal2 8786 33150 8786 33150 0 debounce2_a.button_hist\[3\]
rlabel metal1 10580 33082 10580 33082 0 debounce2_a.button_hist\[4\]
rlabel metal1 9614 33388 9614 33388 0 debounce2_a.button_hist\[5\]
rlabel metal1 11592 32878 11592 32878 0 debounce2_a.button_hist\[6\]
rlabel metal1 10902 32334 10902 32334 0 debounce2_a.button_hist\[7\]
rlabel metal1 12374 27914 12374 27914 0 debounce2_a.debounced
rlabel metal1 9384 29274 9384 29274 0 debounce2_b.button_hist\[0\]
rlabel metal1 8786 29070 8786 29070 0 debounce2_b.button_hist\[1\]
rlabel metal1 9430 28050 9430 28050 0 debounce2_b.button_hist\[2\]
rlabel metal1 9568 28594 9568 28594 0 debounce2_b.button_hist\[3\]
rlabel metal1 10442 28526 10442 28526 0 debounce2_b.button_hist\[4\]
rlabel metal1 10442 30906 10442 30906 0 debounce2_b.button_hist\[5\]
rlabel metal1 10350 28934 10350 28934 0 debounce2_b.button_hist\[6\]
rlabel metal1 10534 28390 10534 28390 0 debounce2_b.button_hist\[7\]
rlabel metal1 11546 29478 11546 29478 0 debounce2_b.debounced
rlabel metal1 14996 39406 14996 39406 0 enc0_a
rlabel metal1 34868 35054 34868 35054 0 enc0_b
rlabel metal1 34868 13294 34868 13294 0 enc1_a
rlabel metal1 8556 39406 8556 39406 0 enc1_b
rlabel metal3 751 28628 751 28628 0 enc2_a
rlabel metal3 820 14348 820 14348 0 enc2_b
rlabel metal1 16100 35054 16100 35054 0 encoder0.old_a
rlabel metal1 16100 35122 16100 35122 0 encoder0.old_b
rlabel metal1 14352 32470 14352 32470 0 encoder0.value\[0\]
rlabel metal1 13938 32980 13938 32980 0 encoder0.value\[1\]
rlabel via1 15870 29597 15870 29597 0 encoder0.value\[2\]
rlabel metal1 17342 31348 17342 31348 0 encoder0.value\[3\]
rlabel metal1 18354 34714 18354 34714 0 encoder0.value\[4\]
rlabel metal1 17618 30906 17618 30906 0 encoder0.value\[5\]
rlabel metal1 19734 32844 19734 32844 0 encoder0.value\[6\]
rlabel metal1 20516 31450 20516 31450 0 encoder0.value\[7\]
rlabel metal1 23414 29138 23414 29138 0 encoder1.old_a
rlabel metal1 23460 29070 23460 29070 0 encoder1.old_b
rlabel metal1 21436 24650 21436 24650 0 encoder1.value\[0\]
rlabel metal1 19872 27098 19872 27098 0 encoder1.value\[1\]
rlabel metal2 24610 26605 24610 26605 0 encoder1.value\[2\]
rlabel metal1 20010 24616 20010 24616 0 encoder1.value\[3\]
rlabel metal2 20562 23137 20562 23137 0 encoder1.value\[4\]
rlabel metal1 20562 22508 20562 22508 0 encoder1.value\[5\]
rlabel metal2 20838 20162 20838 20162 0 encoder1.value\[6\]
rlabel metal1 22954 21454 22954 21454 0 encoder1.value\[7\]
rlabel metal1 13110 29172 13110 29172 0 encoder2.old_a
rlabel metal2 13202 28934 13202 28934 0 encoder2.old_b
rlabel metal1 15134 24174 15134 24174 0 encoder2.value\[0\]
rlabel metal1 15732 24038 15732 24038 0 encoder2.value\[1\]
rlabel metal1 14904 26486 14904 26486 0 encoder2.value\[2\]
rlabel metal1 14076 23290 14076 23290 0 encoder2.value\[3\]
rlabel metal1 12788 26758 12788 26758 0 encoder2.value\[4\]
rlabel metal2 11546 22039 11546 22039 0 encoder2.value\[5\]
rlabel metal1 10442 24174 10442 24174 0 encoder2.value\[6\]
rlabel metal1 11178 23290 11178 23290 0 encoder2.value\[7\]
rlabel metal1 14490 39372 14490 39372 0 net1
rlabel metal1 9430 21964 9430 21964 0 net10
rlabel metal1 15456 37230 15456 37230 0 net100
rlabel metal1 13662 32368 13662 32368 0 net101
rlabel metal1 12967 32878 12967 32878 0 net102
rlabel metal1 9660 31246 9660 31246 0 net103
rlabel metal1 15410 24786 15410 24786 0 net104
rlabel metal1 17265 24106 17265 24106 0 net105
rlabel metal1 8832 31382 8832 31382 0 net106
rlabel metal1 21252 27438 21252 27438 0 net107
rlabel metal1 20980 27030 20980 27030 0 net108
rlabel metal1 23368 35598 23368 35598 0 net109
rlabel metal1 26220 20400 26220 20400 0 net11
rlabel metal1 15732 39406 15732 39406 0 net110
rlabel metal2 11270 35802 11270 35802 0 net111
rlabel metal2 11822 28492 11822 28492 0 net112
rlabel metal1 12512 35598 12512 35598 0 net113
rlabel metal1 11454 23562 11454 23562 0 net114
rlabel via1 12194 23086 12194 23086 0 net115
rlabel metal1 22264 34510 22264 34510 0 net116
rlabel metal1 16422 36108 16422 36108 0 net117
rlabel metal1 21574 37740 21574 37740 0 net118
rlabel metal1 22218 20910 22218 20910 0 net119
rlabel metal2 7314 37468 7314 37468 0 net12
rlabel metal1 22954 20502 22954 20502 0 net120
rlabel metal1 21620 36754 21620 36754 0 net121
rlabel metal1 10028 34510 10028 34510 0 net122
rlabel metal1 14168 36890 14168 36890 0 net123
rlabel metal1 20424 32402 20424 32402 0 net124
rlabel via1 21026 31382 21026 31382 0 net125
rlabel metal1 23276 30770 23276 30770 0 net126
rlabel metal1 13294 23562 13294 23562 0 net127
rlabel metal1 12875 23018 12875 23018 0 net128
rlabel metal1 14628 31926 14628 31926 0 net129
rlabel metal2 13570 1027 13570 1027 0 net13
rlabel metal1 13151 31382 13151 31382 0 net130
rlabel metal1 23874 26962 23874 26962 0 net131
rlabel metal1 23731 27030 23731 27030 0 net132
rlabel metal1 21528 22610 21528 22610 0 net133
rlabel metal1 23639 23766 23639 23766 0 net134
rlabel metal2 15134 26316 15134 26316 0 net135
rlabel via1 15874 26350 15874 26350 0 net136
rlabel metal1 19182 37434 19182 37434 0 net137
rlabel metal1 18952 19482 18952 19482 0 net138
rlabel metal2 13018 26554 13018 26554 0 net139
rlabel metal3 1050 6868 1050 6868 0 net14
rlabel metal1 13712 27030 13712 27030 0 net140
rlabel metal1 16974 33456 16974 33456 0 net141
rlabel metal1 15175 33966 15175 33966 0 net142
rlabel metal1 16054 31790 16054 31790 0 net143
rlabel metal1 16038 30634 16038 30634 0 net144
rlabel metal1 23966 24786 23966 24786 0 net145
rlabel via1 23133 25262 23133 25262 0 net146
rlabel metal1 15088 23154 15088 23154 0 net147
rlabel metal1 15313 22678 15313 22678 0 net148
rlabel metal1 23966 21998 23966 21998 0 net149
rlabel via2 34546 27421 34546 27421 0 net15
rlabel metal1 23225 22678 23225 22678 0 net150
rlabel metal1 21298 24922 21298 24922 0 net151
rlabel metal1 20332 24378 20332 24378 0 net152
rlabel metal1 20700 20570 20700 20570 0 net153
rlabel metal1 20286 20400 20286 20400 0 net154
rlabel metal1 16698 35530 16698 35530 0 net155
rlabel metal1 10994 29036 10994 29036 0 net156
rlabel metal1 12742 25296 12742 25296 0 net157
rlabel metal2 10718 26112 10718 26112 0 net158
rlabel metal2 12558 24548 12558 24548 0 net159
rlabel metal3 820 36108 820 36108 0 net16
rlabel metal1 9706 23732 9706 23732 0 net160
rlabel metal1 18860 32402 18860 32402 0 net161
rlabel metal1 18916 30702 18916 30702 0 net162
rlabel metal1 17066 35734 17066 35734 0 net163
rlabel metal1 23874 29614 23874 29614 0 net164
rlabel metal1 17986 34000 17986 34000 0 net165
rlabel metal1 18588 34646 18588 34646 0 net166
rlabel metal2 12374 31484 12374 31484 0 net167
rlabel metal1 20884 29614 20884 29614 0 net168
rlabel metal2 21390 33626 21390 33626 0 net169
rlabel via2 34546 5627 34546 5627 0 net17
rlabel metal1 20608 33966 20608 33966 0 net170
rlabel metal2 3082 39236 3082 39236 0 net171
rlabel metal1 1610 39406 1610 39406 0 net172
rlabel metal1 16836 21522 16836 21522 0 net173
rlabel metal1 16656 20910 16656 20910 0 net174
rlabel metal2 17618 25806 17618 25806 0 net175
rlabel via1 16969 25874 16969 25874 0 net176
rlabel metal2 27094 959 27094 959 0 net18
rlabel metal2 46 1520 46 1520 0 net19
rlabel metal1 33051 34918 33051 34918 0 net2
rlabel metal1 35006 39474 35006 39474 0 net20
rlabel metal2 6486 959 6486 959 0 net21
rlabel metal2 34178 959 34178 959 0 net22
rlabel metal1 2484 39406 2484 39406 0 net23
rlabel metal1 7406 36142 7406 36142 0 net24
rlabel metal2 8050 37026 8050 37026 0 net25
rlabel metal1 14820 29206 14820 29206 0 net26
rlabel metal2 14214 27846 14214 27846 0 net27
rlabel metal1 14168 20910 14168 20910 0 net28
rlabel metal1 16483 20502 16483 20502 0 net29
rlabel metal1 29210 13158 29210 13158 0 net3
rlabel metal1 22678 33354 22678 33354 0 net30
rlabel metal2 22494 31969 22494 31969 0 net31
rlabel metal1 20930 36550 20930 36550 0 net32
rlabel metal1 21348 34986 21348 34986 0 net33
rlabel metal2 11178 30600 11178 30600 0 net34
rlabel metal1 12016 29614 12016 29614 0 net35
rlabel metal1 17710 36108 17710 36108 0 net36
rlabel metal1 16872 36754 16872 36754 0 net37
rlabel metal2 13018 35394 13018 35394 0 net38
rlabel metal1 14531 36142 14531 36142 0 net39
rlabel metal2 8510 38794 8510 38794 0 net4
rlabel metal1 18354 25262 18354 25262 0 net40
rlabel via1 16509 25262 16509 25262 0 net41
rlabel metal1 9522 33626 9522 33626 0 net42
rlabel metal1 11270 32742 11270 32742 0 net43
rlabel metal1 19412 29070 19412 29070 0 net44
rlabel metal1 18528 28050 18528 28050 0 net45
rlabel metal1 17388 29070 17388 29070 0 net46
rlabel metal1 17199 28050 17199 28050 0 net47
rlabel metal1 19182 22406 19182 22406 0 net48
rlabel via1 17981 21998 17981 21998 0 net49
rlabel metal2 6118 29444 6118 29444 0 net5
rlabel metal1 13110 20978 13110 20978 0 net50
rlabel via1 12746 19822 12746 19822 0 net51
rlabel metal1 10396 20774 10396 20774 0 net52
rlabel metal1 9460 20502 9460 20502 0 net53
rlabel metal1 14858 28968 14858 28968 0 net54
rlabel metal1 14577 29614 14577 29614 0 net55
rlabel metal1 20470 28594 20470 28594 0 net56
rlabel via1 19913 29138 19913 29138 0 net57
rlabel metal2 15778 28220 15778 28220 0 net58
rlabel metal1 15456 28186 15456 28186 0 net59
rlabel metal2 1610 21862 1610 21862 0 net6
rlabel metal1 16606 21658 16606 21658 0 net60
rlabel metal1 18032 23018 18032 23018 0 net61
rlabel metal2 17342 23494 17342 23494 0 net62
rlabel metal2 17434 25194 17434 25194 0 net63
rlabel metal1 15594 20842 15594 20842 0 net64
rlabel metal1 14761 19822 14761 19822 0 net65
rlabel metal1 17940 26962 17940 26962 0 net66
rlabel metal1 17884 26350 17884 26350 0 net67
rlabel metal1 9430 35768 9430 35768 0 net68
rlabel metal1 19458 29206 19458 29206 0 net69
rlabel metal1 6210 38318 6210 38318 0 net7
rlabel metal1 18441 27438 18441 27438 0 net70
rlabel metal2 12466 19856 12466 19856 0 net71
rlabel metal2 10626 19618 10626 19618 0 net72
rlabel metal1 17940 21658 17940 21658 0 net73
rlabel metal1 17291 21590 17291 21590 0 net74
rlabel metal1 9614 21590 9614 21590 0 net75
rlabel metal1 9430 21658 9430 21658 0 net76
rlabel metal1 16790 38862 16790 38862 0 net77
rlabel metal1 10810 28662 10810 28662 0 net78
rlabel metal2 9062 27676 9062 27676 0 net79
rlabel metal1 22678 39406 22678 39406 0 net8
rlabel metal1 8648 28186 8648 28186 0 net80
rlabel metal1 19412 24038 19412 24038 0 net81
rlabel metal1 22540 37298 22540 37298 0 net82
rlabel metal2 12558 33524 12558 33524 0 net83
rlabel metal1 8694 29138 8694 29138 0 net84
rlabel metal1 13662 21454 13662 21454 0 net85
rlabel metal1 10810 36346 10810 36346 0 net86
rlabel metal1 8050 28594 8050 28594 0 net87
rlabel metal1 9108 34170 9108 34170 0 net88
rlabel metal1 18216 38522 18216 38522 0 net89
rlabel metal2 20286 7417 20286 7417 0 net9
rlabel metal1 22540 38386 22540 38386 0 net90
rlabel metal2 25530 32674 25530 32674 0 net91
rlabel metal1 24840 34034 24840 34034 0 net92
rlabel metal1 7912 32946 7912 32946 0 net93
rlabel metal1 25254 30770 25254 30770 0 net94
rlabel metal1 24472 33082 24472 33082 0 net95
rlabel metal1 12696 36210 12696 36210 0 net96
rlabel metal1 23782 38386 23782 38386 0 net97
rlabel metal1 10488 36074 10488 36074 0 net98
rlabel metal1 17204 28662 17204 28662 0 net99
rlabel metal1 15364 27438 15364 27438 0 pwm0.count\[0\]
rlabel metal1 15548 29818 15548 29818 0 pwm0.count\[1\]
rlabel metal1 14766 29138 14766 29138 0 pwm0.count\[2\]
rlabel metal2 16054 28084 16054 28084 0 pwm0.count\[3\]
rlabel metal2 18262 29648 18262 29648 0 pwm0.count\[4\]
rlabel metal1 19458 27302 19458 27302 0 pwm0.count\[5\]
rlabel metal1 20102 28628 20102 28628 0 pwm0.count\[6\]
rlabel metal2 21022 29750 21022 29750 0 pwm0.count\[7\]
rlabel metal2 21942 40368 21942 40368 0 pwm0_out
rlabel metal1 17710 25364 17710 25364 0 pwm1.count\[0\]
rlabel metal2 18446 26316 18446 26316 0 pwm1.count\[1\]
rlabel metal1 19504 26486 19504 26486 0 pwm1.count\[2\]
rlabel metal2 19458 25058 19458 25058 0 pwm1.count\[3\]
rlabel via1 19642 23154 19642 23154 0 pwm1.count\[4\]
rlabel metal1 20148 21930 20148 21930 0 pwm1.count\[5\]
rlabel metal1 20007 21998 20007 21998 0 pwm1.count\[6\]
rlabel metal1 20332 21454 20332 21454 0 pwm1.count\[7\]
rlabel metal2 20654 1095 20654 1095 0 pwm1_out
rlabel metal1 15042 20570 15042 20570 0 pwm2.count\[0\]
rlabel metal1 15226 22032 15226 22032 0 pwm2.count\[1\]
rlabel metal1 15456 19958 15456 19958 0 pwm2.count\[2\]
rlabel metal1 13984 21114 13984 21114 0 pwm2.count\[3\]
rlabel metal2 12834 20298 12834 20298 0 pwm2.count\[4\]
rlabel metal2 11960 21522 11960 21522 0 pwm2.count\[5\]
rlabel metal1 11040 21522 11040 21522 0 pwm2.count\[6\]
rlabel metal1 10626 22134 10626 22134 0 pwm2.count\[7\]
rlabel metal3 820 21828 820 21828 0 pwm2_out
rlabel metal1 1380 38930 1380 38930 0 reset
rlabel metal3 34922 19788 34922 19788 0 sync
<< properties >>
string FIXED_BBOX 0 0 36000 42000
<< end >>
