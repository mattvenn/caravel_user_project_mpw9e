magic
tech sky130A
magscale 1 2
timestamp 1696494446
<< obsli1 >>
rect 1104 2159 34868 39729
<< obsm1 >>
rect 14 2128 35498 39760
<< metal2 >>
rect 1278 41200 1390 42000
rect 8362 41200 8474 42000
rect 14802 41200 14914 42000
rect 21886 41200 21998 42000
rect 28970 41200 29082 42000
rect 35410 41200 35522 42000
rect -10 0 102 800
rect 6430 0 6542 800
rect 13514 0 13626 800
rect 20598 0 20710 800
rect 27038 0 27150 800
rect 34122 0 34234 800
<< obsm2 >>
rect 20 41144 1222 41200
rect 1446 41144 8306 41200
rect 8530 41144 14746 41200
rect 14970 41144 21830 41200
rect 22054 41144 28914 41200
rect 29138 41144 35354 41200
rect 20 856 35492 41144
rect 158 800 6374 856
rect 6598 800 13458 856
rect 13682 800 20542 856
rect 20766 800 26982 856
rect 27206 800 34066 856
rect 34290 800 35492 856
<< metal3 >>
rect 0 35988 800 36228
rect 35200 34628 36000 34868
rect 0 28508 800 28748
rect 35200 27148 36000 27388
rect 0 21708 800 21948
rect 35200 19668 36000 19908
rect 0 14228 800 14468
rect 35200 12868 36000 13108
rect 0 6748 800 6988
rect 35200 5388 36000 5628
<< obsm3 >>
rect 798 36308 35220 39745
rect 880 35908 35220 36308
rect 798 34948 35220 35908
rect 798 34548 35120 34948
rect 798 28828 35220 34548
rect 880 28428 35220 28828
rect 798 27468 35220 28428
rect 798 27068 35120 27468
rect 798 22028 35220 27068
rect 880 21628 35220 22028
rect 798 19988 35220 21628
rect 798 19588 35120 19988
rect 798 14548 35220 19588
rect 880 14148 35220 14548
rect 798 13188 35220 14148
rect 798 12788 35120 13188
rect 798 7068 35220 12788
rect 880 6668 35220 7068
rect 798 5708 35220 6668
rect 798 5308 35120 5708
rect 798 2143 35220 5308
<< metal4 >>
rect 5164 2128 5484 39760
rect 9384 2128 9704 39760
rect 13605 2128 13925 39760
rect 17825 2128 18145 39760
rect 22046 2128 22366 39760
rect 26266 2128 26586 39760
rect 30487 2128 30807 39760
rect 34707 2128 35027 39760
<< labels >>
rlabel metal2 s 28970 41200 29082 42000 6 clk
port 1 nsew signal input
rlabel metal2 s 14802 41200 14914 42000 6 enc0_a
port 2 nsew signal input
rlabel metal3 s 35200 34628 36000 34868 6 enc0_b
port 3 nsew signal input
rlabel metal3 s 35200 12868 36000 13108 6 enc1_a
port 4 nsew signal input
rlabel metal2 s 8362 41200 8474 42000 6 enc1_b
port 5 nsew signal input
rlabel metal3 s 0 28508 800 28748 6 enc2_a
port 6 nsew signal input
rlabel metal3 s 0 14228 800 14468 6 enc2_b
port 7 nsew signal input
rlabel metal3 s 35200 5388 36000 5628 6 io_oeb_high[0]
port 8 nsew signal output
rlabel metal2 s 27038 0 27150 800 6 io_oeb_high[1]
port 9 nsew signal output
rlabel metal2 s -10 0 102 800 6 io_oeb_high[2]
port 10 nsew signal output
rlabel metal2 s 35410 41200 35522 42000 6 io_oeb_high[3]
port 11 nsew signal output
rlabel metal2 s 6430 0 6542 800 6 io_oeb_high[4]
port 12 nsew signal output
rlabel metal2 s 34122 0 34234 800 6 io_oeb_high[5]
port 13 nsew signal output
rlabel metal2 s 13514 0 13626 800 6 io_oeb_low[0]
port 14 nsew signal output
rlabel metal3 s 0 6748 800 6988 6 io_oeb_low[1]
port 15 nsew signal output
rlabel metal3 s 35200 27148 36000 27388 6 io_oeb_low[2]
port 16 nsew signal output
rlabel metal3 s 0 35988 800 36228 6 io_oeb_low[3]
port 17 nsew signal output
rlabel metal2 s 21886 41200 21998 42000 6 pwm0_out
port 18 nsew signal output
rlabel metal2 s 20598 0 20710 800 6 pwm1_out
port 19 nsew signal output
rlabel metal3 s 0 21708 800 21948 6 pwm2_out
port 20 nsew signal output
rlabel metal2 s 1278 41200 1390 42000 6 reset
port 21 nsew signal input
rlabel metal3 s 35200 19668 36000 19908 6 sync
port 22 nsew signal output
rlabel metal4 s 5164 2128 5484 39760 6 vccd1
port 23 nsew power bidirectional
rlabel metal4 s 13605 2128 13925 39760 6 vccd1
port 23 nsew power bidirectional
rlabel metal4 s 22046 2128 22366 39760 6 vccd1
port 23 nsew power bidirectional
rlabel metal4 s 30487 2128 30807 39760 6 vccd1
port 23 nsew power bidirectional
rlabel metal4 s 9384 2128 9704 39760 6 vssd1
port 24 nsew ground bidirectional
rlabel metal4 s 17825 2128 18145 39760 6 vssd1
port 24 nsew ground bidirectional
rlabel metal4 s 26266 2128 26586 39760 6 vssd1
port 24 nsew ground bidirectional
rlabel metal4 s 34707 2128 35027 39760 6 vssd1
port 24 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 36000 42000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 2114130
string GDS_FILE /home/zerotoasic/asic_tools/caravel_user_project/openlane/rgb_mixer/runs/23_10_05_10_25/results/signoff/rgb_mixer.magic.gds
string GDS_START 307968
<< end >>

