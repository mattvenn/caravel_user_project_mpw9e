magic
tech sky130A
magscale 1 2
timestamp 1696431772
<< obsli1 >>
rect 1104 2159 34868 39729
<< obsm1 >>
rect 14 2128 35498 39760
<< metal2 >>
rect 7074 41200 7186 42000
rect 16734 41200 16846 42000
rect 26394 41200 26506 42000
rect 35410 41200 35522 42000
rect -10 0 102 800
rect 9006 0 9118 800
rect 18666 0 18778 800
rect 28326 0 28438 800
<< obsm2 >>
rect 20 41144 7018 41200
rect 7242 41144 16678 41200
rect 16902 41144 26338 41200
rect 26562 41144 35354 41200
rect 20 856 35492 41144
rect 158 800 8950 856
rect 9174 800 18610 856
rect 18834 800 28270 856
rect 28494 800 35492 856
<< metal3 >>
rect 0 39388 800 39628
rect 35200 31908 36000 32148
rect 0 29868 800 30108
rect 35200 21708 36000 21948
rect 0 19668 800 19908
rect 35200 11508 36000 11748
rect 0 9468 800 9708
rect 35200 1988 36000 2228
<< obsm3 >>
rect 800 39708 35266 39745
rect 880 39308 35266 39708
rect 800 32228 35266 39308
rect 800 31828 35120 32228
rect 800 30188 35266 31828
rect 880 29788 35266 30188
rect 800 22028 35266 29788
rect 800 21628 35120 22028
rect 800 19988 35266 21628
rect 880 19588 35266 19988
rect 800 11828 35266 19588
rect 800 11428 35120 11828
rect 800 9788 35266 11428
rect 880 9388 35266 9788
rect 800 2308 35266 9388
rect 800 2075 35120 2308
<< metal4 >>
rect 5164 2128 5484 39760
rect 9384 2128 9704 39760
rect 13605 2128 13925 39760
rect 17825 2128 18145 39760
rect 22046 2128 22366 39760
rect 26266 2128 26586 39760
rect 30487 2128 30807 39760
rect 34707 2128 35027 39760
<< labels >>
rlabel metal3 s 35200 21708 36000 21948 6 clk
port 1 nsew signal input
rlabel metal3 s 0 39388 800 39628 6 enc0_a
port 2 nsew signal input
rlabel metal3 s 35200 31908 36000 32148 6 enc0_b
port 3 nsew signal input
rlabel metal3 s 35200 1988 36000 2228 6 enc1_a
port 4 nsew signal input
rlabel metal2 s 16734 41200 16846 42000 6 enc1_b
port 5 nsew signal input
rlabel metal2 s -10 0 102 800 6 enc2_a
port 6 nsew signal input
rlabel metal2 s 28326 0 28438 800 6 enc2_b
port 7 nsew signal input
rlabel metal2 s 9006 0 9118 800 6 io_oeb[0]
port 8 nsew signal output
rlabel metal2 s 26394 41200 26506 42000 6 io_oeb[1]
port 9 nsew signal output
rlabel metal3 s 0 9468 800 9708 6 io_oeb[2]
port 10 nsew signal output
rlabel metal3 s 0 19668 800 19908 6 io_oeb[3]
port 11 nsew signal output
rlabel metal2 s 35410 41200 35522 42000 6 pwm0_out
port 12 nsew signal output
rlabel metal2 s 18666 0 18778 800 6 pwm1_out
port 13 nsew signal output
rlabel metal3 s 0 29868 800 30108 6 pwm2_out
port 14 nsew signal output
rlabel metal2 s 7074 41200 7186 42000 6 reset
port 15 nsew signal input
rlabel metal3 s 35200 11508 36000 11748 6 sync
port 16 nsew signal output
rlabel metal4 s 5164 2128 5484 39760 6 vccd1
port 17 nsew power bidirectional
rlabel metal4 s 13605 2128 13925 39760 6 vccd1
port 17 nsew power bidirectional
rlabel metal4 s 22046 2128 22366 39760 6 vccd1
port 17 nsew power bidirectional
rlabel metal4 s 30487 2128 30807 39760 6 vccd1
port 17 nsew power bidirectional
rlabel metal4 s 9384 2128 9704 39760 6 vssd1
port 18 nsew ground bidirectional
rlabel metal4 s 17825 2128 18145 39760 6 vssd1
port 18 nsew ground bidirectional
rlabel metal4 s 26266 2128 26586 39760 6 vssd1
port 18 nsew ground bidirectional
rlabel metal4 s 34707 2128 35027 39760 6 vssd1
port 18 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 36000 42000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 1885278
string GDS_FILE /home/zerotoasic/asic_tools/caravel_user_project/openlane/rgb_mixer/runs/23_10_04_17_00/results/signoff/rgb_mixer.magic.gds
string GDS_START 275110
<< end >>

