magic
tech sky130A
magscale 1 2
timestamp 1696431770
<< viali >>
rect 26525 39593 26559 39627
rect 34437 39593 34471 39627
rect 1409 39389 1443 39423
rect 7205 39389 7239 39423
rect 16865 39389 16899 39423
rect 34161 39321 34195 39355
rect 1593 39253 1627 39287
rect 7389 39253 7423 39287
rect 17049 39253 17083 39287
rect 26341 33949 26375 33983
rect 26525 33949 26559 33983
rect 26433 33813 26467 33847
rect 27169 33541 27203 33575
rect 23121 33473 23155 33507
rect 23949 33473 23983 33507
rect 25881 33473 25915 33507
rect 26341 33473 26375 33507
rect 26801 33473 26835 33507
rect 26985 33473 27019 33507
rect 28632 33473 28666 33507
rect 29837 33473 29871 33507
rect 30113 33473 30147 33507
rect 30573 33473 30607 33507
rect 31033 33473 31067 33507
rect 22937 33405 22971 33439
rect 25973 33405 26007 33439
rect 26433 33405 26467 33439
rect 28365 33405 28399 33439
rect 30021 33405 30055 33439
rect 30389 33405 30423 33439
rect 26249 33337 26283 33371
rect 26525 33337 26559 33371
rect 29745 33337 29779 33371
rect 30757 33337 30791 33371
rect 23305 33269 23339 33303
rect 24133 33269 24167 33303
rect 26663 33269 26697 33303
rect 27353 33269 27387 33303
rect 29929 33269 29963 33303
rect 30297 33269 30331 33303
rect 30849 33269 30883 33303
rect 24225 33065 24259 33099
rect 29561 33065 29595 33099
rect 28641 32997 28675 33031
rect 24409 32929 24443 32963
rect 26341 32929 26375 32963
rect 26709 32929 26743 32963
rect 27261 32929 27295 32963
rect 28733 32929 28767 32963
rect 23581 32861 23615 32895
rect 23949 32861 23983 32895
rect 24041 32861 24075 32895
rect 24665 32861 24699 32895
rect 26065 32861 26099 32895
rect 26249 32861 26283 32895
rect 26617 32861 26651 32895
rect 28917 32861 28951 32895
rect 29101 32861 29135 32895
rect 29377 32861 29411 32895
rect 29745 32861 29779 32895
rect 31217 32861 31251 32895
rect 31493 32861 31527 32895
rect 27506 32793 27540 32827
rect 30972 32793 31006 32827
rect 23765 32725 23799 32759
rect 25789 32725 25823 32759
rect 25881 32725 25915 32759
rect 26433 32725 26467 32759
rect 27077 32725 27111 32759
rect 29193 32725 29227 32759
rect 29837 32725 29871 32759
rect 31309 32725 31343 32759
rect 26985 32521 27019 32555
rect 27537 32521 27571 32555
rect 29929 32521 29963 32555
rect 30113 32521 30147 32555
rect 29745 32453 29779 32487
rect 30748 32453 30782 32487
rect 17601 32385 17635 32419
rect 18696 32385 18730 32419
rect 20269 32385 20303 32419
rect 21005 32385 21039 32419
rect 22946 32385 22980 32419
rect 23213 32385 23247 32419
rect 25441 32385 25475 32419
rect 25697 32385 25731 32419
rect 25789 32385 25823 32419
rect 25973 32385 26007 32419
rect 26065 32385 26099 32419
rect 26341 32385 26375 32419
rect 26801 32385 26835 32419
rect 27166 32383 27200 32417
rect 27445 32385 27479 32419
rect 27629 32385 27663 32419
rect 29121 32385 29155 32419
rect 29377 32385 29411 32419
rect 30021 32385 30055 32419
rect 34529 32385 34563 32419
rect 17877 32317 17911 32351
rect 18429 32317 18463 32351
rect 20085 32317 20119 32351
rect 20729 32317 20763 32351
rect 26157 32317 26191 32351
rect 27353 32317 27387 32351
rect 30481 32317 30515 32351
rect 19809 32249 19843 32283
rect 20453 32249 20487 32283
rect 26525 32249 26559 32283
rect 17417 32181 17451 32215
rect 17785 32181 17819 32215
rect 20821 32181 20855 32215
rect 21189 32181 21223 32215
rect 21833 32181 21867 32215
rect 24317 32181 24351 32215
rect 26709 32181 26743 32215
rect 27997 32181 28031 32215
rect 30297 32181 30331 32215
rect 31861 32181 31895 32215
rect 34345 32181 34379 32215
rect 18429 31977 18463 32011
rect 18981 31977 19015 32011
rect 20729 31977 20763 32011
rect 21741 31977 21775 32011
rect 26157 31977 26191 32011
rect 26249 31977 26283 32011
rect 29101 31977 29135 32011
rect 31125 31977 31159 32011
rect 20591 31909 20625 31943
rect 20821 31909 20855 31943
rect 25973 31909 26007 31943
rect 19901 31841 19935 31875
rect 26157 31841 26191 31875
rect 28733 31841 28767 31875
rect 30757 31841 30791 31875
rect 32229 31841 32263 31875
rect 17049 31773 17083 31807
rect 17316 31773 17350 31807
rect 18797 31773 18831 31807
rect 18981 31773 19015 31807
rect 19625 31773 19659 31807
rect 19993 31773 20027 31807
rect 20453 31773 20487 31807
rect 20913 31773 20947 31807
rect 21005 31773 21039 31807
rect 21189 31773 21223 31807
rect 21281 31773 21315 31807
rect 21419 31773 21453 31807
rect 21557 31773 21591 31807
rect 21833 31773 21867 31807
rect 22017 31773 22051 31807
rect 26341 31773 26375 31807
rect 28917 31773 28951 31807
rect 30481 31773 30515 31807
rect 30665 31773 30699 31807
rect 30941 31773 30975 31807
rect 31401 31773 31435 31807
rect 31585 31773 31619 31807
rect 31861 31773 31895 31807
rect 32059 31773 32093 31807
rect 19533 31637 19567 31671
rect 19717 31637 19751 31671
rect 20361 31637 20395 31671
rect 21925 31637 21959 31671
rect 30297 31637 30331 31671
rect 31769 31637 31803 31671
rect 18245 31433 18279 31467
rect 19257 31433 19291 31467
rect 20269 31433 20303 31467
rect 21005 31433 21039 31467
rect 23121 31433 23155 31467
rect 31309 31433 31343 31467
rect 32137 31433 32171 31467
rect 21097 31365 21131 31399
rect 21281 31365 21315 31399
rect 16937 31297 16971 31331
rect 18153 31297 18187 31331
rect 18429 31297 18463 31331
rect 19441 31297 19475 31331
rect 19533 31297 19567 31331
rect 19809 31297 19843 31331
rect 20085 31297 20119 31331
rect 20177 31297 20211 31331
rect 20361 31297 20395 31331
rect 20637 31297 20671 31331
rect 23305 31297 23339 31331
rect 23397 31297 23431 31331
rect 23664 31297 23698 31331
rect 24869 31297 24903 31331
rect 25053 31297 25087 31331
rect 25237 31297 25271 31331
rect 25421 31297 25455 31331
rect 27905 31297 27939 31331
rect 28089 31297 28123 31331
rect 29929 31297 29963 31331
rect 30389 31297 30423 31331
rect 30665 31297 30699 31331
rect 30849 31297 30883 31331
rect 31217 31297 31251 31331
rect 31585 31297 31619 31331
rect 31861 31297 31895 31331
rect 33250 31297 33284 31331
rect 33517 31297 33551 31331
rect 16681 31229 16715 31263
rect 20729 31229 20763 31263
rect 25329 31229 25363 31263
rect 31125 31229 31159 31263
rect 31493 31229 31527 31263
rect 18429 31161 18463 31195
rect 19717 31161 19751 31195
rect 30481 31161 30515 31195
rect 30573 31161 30607 31195
rect 18061 31093 18095 31127
rect 19993 31093 20027 31127
rect 21465 31093 21499 31127
rect 24777 31093 24811 31127
rect 25513 31093 25547 31127
rect 28089 31093 28123 31127
rect 29745 31093 29779 31127
rect 30113 31093 30147 31127
rect 30941 31093 30975 31127
rect 31769 31093 31803 31127
rect 16773 30889 16807 30923
rect 17601 30889 17635 30923
rect 17785 30889 17819 30923
rect 24685 30889 24719 30923
rect 27261 30889 27295 30923
rect 32413 30889 32447 30923
rect 32689 30889 32723 30923
rect 17877 30821 17911 30855
rect 25421 30821 25455 30855
rect 26985 30821 27019 30855
rect 27537 30821 27571 30855
rect 27905 30821 27939 30855
rect 18245 30753 18279 30787
rect 25881 30753 25915 30787
rect 26709 30753 26743 30787
rect 28181 30753 28215 30787
rect 31033 30753 31067 30787
rect 16957 30685 16991 30719
rect 17141 30685 17175 30719
rect 17233 30685 17267 30719
rect 17877 30685 17911 30719
rect 18061 30685 18095 30719
rect 18521 30685 18555 30719
rect 18797 30685 18831 30719
rect 18981 30685 19015 30719
rect 19257 30685 19291 30719
rect 19441 30685 19475 30719
rect 19533 30685 19567 30719
rect 19625 30685 19659 30719
rect 19809 30685 19843 30719
rect 22017 30685 22051 30719
rect 23673 30685 23707 30719
rect 23765 30685 23799 30719
rect 23949 30685 23983 30719
rect 24133 30685 24167 30719
rect 24409 30685 24443 30719
rect 24501 30685 24535 30719
rect 24869 30685 24903 30719
rect 25237 30685 25271 30719
rect 25513 30685 25547 30719
rect 25697 30685 25731 30719
rect 25789 30685 25823 30719
rect 26065 30685 26099 30719
rect 26617 30685 26651 30719
rect 27445 30685 27479 30719
rect 27629 30685 27663 30719
rect 27721 30685 27755 30719
rect 28273 30685 28307 30719
rect 28733 30685 28767 30719
rect 28825 30685 28859 30719
rect 29561 30685 29595 30719
rect 29828 30685 29862 30719
rect 32505 30685 32539 30719
rect 17417 30617 17451 30651
rect 22284 30617 22318 30651
rect 24685 30617 24719 30651
rect 25053 30617 25087 30651
rect 25145 30617 25179 30651
rect 31300 30617 31334 30651
rect 17617 30549 17651 30583
rect 18337 30549 18371 30583
rect 19993 30549 20027 30583
rect 23397 30549 23431 30583
rect 23489 30549 23523 30583
rect 24041 30549 24075 30583
rect 26249 30549 26283 30583
rect 28549 30549 28583 30583
rect 30941 30549 30975 30583
rect 18061 30345 18095 30379
rect 18981 30345 19015 30379
rect 25881 30345 25915 30379
rect 31401 30345 31435 30379
rect 1777 30277 1811 30311
rect 18613 30277 18647 30311
rect 18705 30277 18739 30311
rect 24869 30277 24903 30311
rect 28733 30277 28767 30311
rect 16313 30209 16347 30243
rect 16497 30209 16531 30243
rect 16937 30209 16971 30243
rect 18337 30209 18371 30243
rect 18457 30209 18491 30243
rect 18843 30209 18877 30243
rect 19257 30209 19291 30243
rect 20269 30209 20303 30243
rect 20453 30209 20487 30243
rect 20729 30209 20763 30243
rect 20913 30209 20947 30243
rect 21097 30209 21131 30243
rect 21281 30209 21315 30243
rect 21465 30209 21499 30243
rect 22946 30209 22980 30243
rect 23213 30209 23247 30243
rect 23305 30209 23339 30243
rect 23561 30209 23595 30243
rect 24777 30209 24811 30243
rect 25145 30209 25179 30243
rect 25329 30209 25363 30243
rect 25421 30209 25455 30243
rect 25697 30209 25731 30243
rect 25973 30209 26007 30243
rect 26157 30209 26191 30243
rect 26341 30209 26375 30243
rect 26525 30209 26559 30243
rect 27261 30209 27295 30243
rect 27629 30209 27663 30243
rect 27721 30209 27755 30243
rect 27813 30209 27847 30243
rect 27997 30209 28031 30243
rect 28549 30209 28583 30243
rect 28641 30209 28675 30243
rect 28825 30209 28859 30243
rect 30113 30209 30147 30243
rect 30205 30209 30239 30243
rect 30297 30209 30331 30243
rect 30481 30209 30515 30243
rect 30665 30209 30699 30243
rect 30757 30209 30791 30243
rect 30941 30209 30975 30243
rect 31217 30209 31251 30243
rect 31861 30209 31895 30243
rect 16681 30141 16715 30175
rect 21005 30141 21039 30175
rect 25513 30141 25547 30175
rect 26249 30141 26283 30175
rect 27169 30141 27203 30175
rect 28273 30141 28307 30175
rect 28457 30141 28491 30175
rect 20637 30073 20671 30107
rect 21833 30073 21867 30107
rect 26985 30073 27019 30107
rect 28365 30073 28399 30107
rect 1501 30005 1535 30039
rect 16497 30005 16531 30039
rect 19165 30005 19199 30039
rect 24685 30005 24719 30039
rect 26709 30005 26743 30039
rect 28181 30005 28215 30039
rect 29837 30005 29871 30039
rect 31677 30005 31711 30039
rect 16681 29801 16715 29835
rect 17233 29801 17267 29835
rect 18153 29801 18187 29835
rect 21189 29801 21223 29835
rect 22661 29801 22695 29835
rect 23305 29801 23339 29835
rect 23673 29801 23707 29835
rect 24041 29801 24075 29835
rect 24225 29801 24259 29835
rect 24961 29801 24995 29835
rect 25145 29801 25179 29835
rect 25973 29801 26007 29835
rect 27629 29801 27663 29835
rect 19809 29733 19843 29767
rect 20453 29733 20487 29767
rect 17141 29665 17175 29699
rect 17601 29665 17635 29699
rect 19533 29665 19567 29699
rect 20361 29665 20395 29699
rect 20729 29665 20763 29699
rect 21281 29665 21315 29699
rect 23121 29665 23155 29699
rect 27721 29665 27755 29699
rect 29561 29665 29595 29699
rect 16865 29597 16899 29631
rect 17049 29597 17083 29631
rect 17417 29597 17451 29631
rect 18337 29597 18371 29631
rect 18521 29597 18555 29631
rect 18613 29597 18647 29631
rect 18705 29597 18739 29631
rect 18889 29597 18923 29631
rect 19441 29597 19475 29631
rect 20269 29597 20303 29631
rect 20545 29597 20579 29631
rect 20821 29597 20855 29631
rect 21005 29597 21039 29631
rect 21465 29597 21499 29631
rect 21557 29597 21591 29631
rect 22845 29597 22879 29631
rect 23029 29597 23063 29631
rect 23489 29597 23523 29631
rect 23765 29597 23799 29631
rect 24869 29597 24903 29631
rect 25324 29597 25358 29631
rect 25421 29597 25455 29631
rect 25696 29597 25730 29631
rect 25789 29597 25823 29631
rect 27086 29597 27120 29631
rect 27353 29597 27387 29631
rect 27445 29597 27479 29631
rect 27537 29597 27571 29631
rect 29377 29597 29411 29631
rect 29828 29597 29862 29631
rect 31309 29597 31343 29631
rect 31576 29597 31610 29631
rect 20085 29529 20119 29563
rect 21281 29529 21315 29563
rect 23857 29529 23891 29563
rect 25513 29529 25547 29563
rect 29110 29529 29144 29563
rect 24057 29461 24091 29495
rect 27997 29461 28031 29495
rect 30941 29461 30975 29495
rect 32689 29461 32723 29495
rect 19073 29257 19107 29291
rect 19717 29257 19751 29291
rect 20821 29257 20855 29291
rect 23029 29257 23063 29291
rect 28917 29257 28951 29291
rect 17049 29121 17083 29155
rect 17233 29121 17267 29155
rect 19165 29121 19199 29155
rect 19625 29121 19659 29155
rect 19809 29121 19843 29155
rect 20071 29121 20105 29155
rect 20361 29121 20395 29155
rect 20637 29121 20671 29155
rect 20821 29121 20855 29155
rect 21097 29121 21131 29155
rect 21281 29121 21315 29155
rect 21373 29121 21407 29155
rect 21833 29121 21867 29155
rect 22017 29121 22051 29155
rect 22937 29121 22971 29155
rect 23121 29121 23155 29155
rect 25053 29121 25087 29155
rect 28273 29121 28307 29155
rect 28436 29124 28470 29158
rect 28549 29121 28583 29155
rect 28641 29121 28675 29155
rect 31585 29121 31619 29155
rect 32137 29121 32171 29155
rect 32321 29121 32355 29155
rect 19901 29053 19935 29087
rect 20913 29053 20947 29087
rect 21649 29053 21683 29087
rect 32505 29053 32539 29087
rect 20269 28985 20303 29019
rect 20499 28985 20533 29019
rect 21465 28985 21499 29019
rect 21833 28985 21867 29019
rect 17049 28917 17083 28951
rect 21557 28917 21591 28951
rect 25145 28917 25179 28951
rect 31769 28917 31803 28951
rect 17785 28713 17819 28747
rect 17969 28713 18003 28747
rect 18797 28713 18831 28747
rect 21281 28713 21315 28747
rect 23673 28713 23707 28747
rect 23857 28713 23891 28747
rect 24777 28713 24811 28747
rect 25881 28713 25915 28747
rect 17693 28645 17727 28679
rect 16313 28577 16347 28611
rect 25513 28577 25547 28611
rect 27537 28577 27571 28611
rect 28089 28577 28123 28611
rect 18245 28509 18279 28543
rect 18613 28509 18647 28543
rect 20545 28509 20579 28543
rect 20729 28509 20763 28543
rect 20821 28509 20855 28543
rect 20913 28509 20947 28543
rect 22661 28509 22695 28543
rect 23029 28509 23063 28543
rect 23213 28509 23247 28543
rect 24685 28509 24719 28543
rect 25145 28509 25179 28543
rect 25329 28509 25363 28543
rect 25421 28509 25455 28543
rect 25697 28509 25731 28543
rect 27261 28509 27295 28543
rect 27353 28509 27387 28543
rect 27813 28509 27847 28543
rect 27905 28509 27939 28543
rect 30021 28509 30055 28543
rect 31585 28509 31619 28543
rect 31852 28509 31886 28543
rect 16580 28441 16614 28475
rect 18153 28441 18187 28475
rect 18429 28441 18463 28475
rect 18521 28441 18555 28475
rect 21189 28441 21223 28475
rect 22394 28441 22428 28475
rect 24041 28441 24075 28475
rect 30288 28441 30322 28475
rect 17943 28373 17977 28407
rect 23121 28373 23155 28407
rect 23831 28373 23865 28407
rect 27537 28373 27571 28407
rect 28089 28373 28123 28407
rect 31401 28373 31435 28407
rect 32965 28373 32999 28407
rect 16865 28169 16899 28203
rect 18613 28169 18647 28203
rect 23673 28169 23707 28203
rect 25145 28169 25179 28203
rect 26801 28169 26835 28203
rect 28181 28169 28215 28203
rect 29009 28169 29043 28203
rect 30389 28169 30423 28203
rect 32321 28169 32355 28203
rect 17417 28101 17451 28135
rect 31493 28101 31527 28135
rect 32505 28101 32539 28135
rect 17049 28033 17083 28067
rect 17233 28033 17267 28067
rect 17601 28033 17635 28067
rect 17877 28033 17911 28067
rect 18061 28033 18095 28067
rect 18245 28033 18279 28067
rect 18429 28033 18463 28067
rect 19349 28033 19383 28067
rect 22293 28033 22327 28067
rect 22560 28033 22594 28067
rect 23765 28033 23799 28067
rect 24032 28033 24066 28067
rect 25688 28033 25722 28067
rect 27169 28033 27203 28067
rect 27721 28033 27755 28067
rect 27997 28033 28031 28067
rect 28457 28033 28491 28067
rect 28917 28033 28951 28067
rect 29101 28033 29135 28067
rect 29193 28033 29227 28067
rect 29377 28033 29411 28067
rect 30573 28033 30607 28067
rect 30665 28033 30699 28067
rect 30849 28033 30883 28067
rect 31033 28033 31067 28067
rect 31125 28033 31159 28067
rect 31769 28033 31803 28067
rect 32137 28033 32171 28067
rect 32413 28033 32447 28067
rect 17325 27965 17359 27999
rect 17785 27965 17819 27999
rect 19441 27965 19475 27999
rect 25421 27965 25455 27999
rect 27261 27965 27295 27999
rect 27905 27965 27939 27999
rect 28549 27965 28583 27999
rect 29285 27965 29319 27999
rect 31677 27965 31711 27999
rect 19717 27897 19751 27931
rect 27537 27897 27571 27931
rect 27813 27897 27847 27931
rect 28825 27897 28859 27931
rect 18061 27829 18095 27863
rect 31309 27829 31343 27863
rect 31677 27829 31711 27863
rect 31953 27829 31987 27863
rect 32689 27829 32723 27863
rect 17969 27625 18003 27659
rect 18245 27625 18279 27659
rect 22937 27625 22971 27659
rect 24225 27625 24259 27659
rect 25237 27625 25271 27659
rect 25973 27625 26007 27659
rect 27813 27625 27847 27659
rect 32413 27625 32447 27659
rect 24593 27557 24627 27591
rect 29561 27557 29595 27591
rect 18337 27489 18371 27523
rect 21005 27489 21039 27523
rect 23305 27489 23339 27523
rect 23581 27489 23615 27523
rect 24409 27489 24443 27523
rect 25145 27489 25179 27523
rect 27633 27489 27667 27523
rect 16589 27421 16623 27455
rect 16856 27421 16890 27455
rect 18061 27421 18095 27455
rect 18153 27421 18187 27455
rect 19073 27421 19107 27455
rect 19717 27421 19751 27455
rect 19809 27421 19843 27455
rect 19901 27421 19935 27455
rect 20085 27421 20119 27455
rect 20361 27421 20395 27455
rect 20621 27421 20655 27455
rect 20729 27421 20763 27455
rect 20821 27421 20855 27455
rect 23121 27421 23155 27455
rect 23397 27421 23431 27455
rect 23765 27421 23799 27455
rect 23949 27421 23983 27455
rect 24041 27421 24075 27455
rect 24225 27421 24259 27455
rect 24685 27421 24719 27455
rect 25421 27421 25455 27455
rect 25513 27421 25547 27455
rect 25605 27421 25639 27455
rect 25789 27421 25823 27455
rect 26249 27421 26283 27455
rect 26341 27421 26375 27455
rect 26433 27421 26467 27455
rect 26617 27421 26651 27455
rect 27261 27421 27295 27455
rect 27445 27421 27479 27455
rect 27537 27421 27571 27455
rect 27905 27421 27939 27455
rect 28733 27421 28767 27455
rect 28917 27421 28951 27455
rect 29009 27421 29043 27455
rect 29101 27421 29135 27455
rect 30941 27421 30975 27455
rect 31033 27421 31067 27455
rect 31300 27421 31334 27455
rect 20177 27353 20211 27387
rect 24409 27353 24443 27387
rect 24777 27353 24811 27387
rect 24961 27353 24995 27387
rect 27077 27353 27111 27387
rect 27629 27353 27663 27387
rect 28365 27353 28399 27387
rect 29377 27353 29411 27387
rect 30674 27353 30708 27387
rect 18981 27285 19015 27319
rect 19441 27285 19475 27319
rect 20545 27285 20579 27319
rect 21005 27285 21039 27319
rect 28089 27285 28123 27319
rect 17141 27081 17175 27115
rect 18245 27081 18279 27115
rect 18337 27081 18371 27115
rect 20729 27081 20763 27115
rect 21097 27081 21131 27115
rect 23397 27081 23431 27115
rect 23673 27081 23707 27115
rect 24961 27081 24995 27115
rect 25881 27081 25915 27115
rect 29101 27081 29135 27115
rect 31217 27081 31251 27115
rect 17969 27013 18003 27047
rect 19450 27013 19484 27047
rect 20085 27013 20119 27047
rect 29285 27013 29319 27047
rect 17141 26945 17175 26979
rect 17601 26945 17635 26979
rect 17694 26945 17728 26979
rect 17877 26945 17911 26979
rect 18107 26945 18141 26979
rect 19809 26945 19843 26979
rect 20269 26945 20303 26979
rect 20545 26945 20579 26979
rect 20821 26945 20855 26979
rect 21189 26945 21223 26979
rect 21373 26945 21407 26979
rect 22946 26945 22980 26979
rect 23213 26945 23247 26979
rect 23581 26945 23615 26979
rect 23857 26945 23891 26979
rect 24869 26945 24903 26979
rect 25329 26945 25363 26979
rect 25513 26945 25547 26979
rect 25605 26945 25639 26979
rect 25697 26945 25731 26979
rect 28733 26945 28767 26979
rect 28917 26945 28951 26979
rect 29193 26945 29227 26979
rect 29377 26945 29411 26979
rect 30941 26945 30975 26979
rect 31033 26945 31067 26979
rect 31677 26945 31711 26979
rect 31769 26945 31803 26979
rect 31953 26945 31987 26979
rect 32505 26945 32539 26979
rect 16865 26877 16899 26911
rect 19717 26877 19751 26911
rect 20085 26877 20119 26911
rect 20361 26877 20395 26911
rect 20453 26877 20487 26911
rect 21097 26877 21131 26911
rect 21281 26877 21315 26911
rect 17049 26809 17083 26843
rect 19901 26741 19935 26775
rect 20913 26741 20947 26775
rect 21833 26741 21867 26775
rect 32321 26741 32355 26775
rect 17693 26537 17727 26571
rect 20177 26537 20211 26571
rect 20913 26537 20947 26571
rect 21189 26537 21223 26571
rect 22017 26537 22051 26571
rect 24409 26537 24443 26571
rect 24593 26537 24627 26571
rect 25237 26537 25271 26571
rect 25881 26537 25915 26571
rect 29009 26537 29043 26571
rect 22661 26469 22695 26503
rect 22753 26469 22787 26503
rect 29837 26469 29871 26503
rect 33333 26469 33367 26503
rect 20729 26401 20763 26435
rect 22201 26401 22235 26435
rect 16313 26333 16347 26367
rect 16580 26333 16614 26367
rect 19349 26333 19383 26367
rect 19441 26333 19475 26367
rect 20637 26333 20671 26367
rect 21089 26335 21123 26369
rect 21281 26333 21315 26367
rect 21373 26333 21407 26367
rect 21557 26333 21591 26367
rect 21649 26333 21683 26367
rect 21741 26333 21775 26367
rect 22109 26333 22143 26367
rect 22293 26333 22327 26367
rect 22753 26333 22787 26367
rect 22845 26333 22879 26367
rect 23101 26333 23135 26367
rect 24869 26333 24903 26367
rect 25421 26333 25455 26367
rect 25605 26333 25639 26367
rect 25789 26333 25823 26367
rect 26249 26333 26283 26367
rect 26341 26333 26375 26367
rect 27169 26333 27203 26367
rect 27353 26333 27387 26367
rect 27445 26333 27479 26367
rect 27537 26333 27571 26367
rect 28089 26333 28123 26367
rect 28825 26333 28859 26367
rect 29561 26333 29595 26367
rect 31953 26333 31987 26367
rect 32220 26333 32254 26367
rect 20269 26265 20303 26299
rect 22477 26265 22511 26299
rect 24777 26265 24811 26299
rect 25513 26265 25547 26299
rect 26065 26265 26099 26299
rect 27905 26265 27939 26299
rect 28273 26265 28307 26299
rect 24225 26197 24259 26231
rect 24577 26197 24611 26231
rect 24961 26197 24995 26231
rect 26433 26197 26467 26231
rect 27813 26197 27847 26231
rect 30021 26197 30055 26231
rect 17509 25993 17543 26027
rect 17677 25993 17711 26027
rect 21097 25993 21131 26027
rect 23765 25993 23799 26027
rect 24133 25993 24167 26027
rect 26709 25993 26743 26027
rect 27261 25993 27295 26027
rect 27629 25993 27663 26027
rect 28349 25993 28383 26027
rect 28641 25993 28675 26027
rect 29377 25993 29411 26027
rect 32597 25993 32631 26027
rect 17877 25925 17911 25959
rect 21281 25925 21315 25959
rect 23949 25925 23983 25959
rect 25881 25925 25915 25959
rect 25973 25925 26007 25959
rect 26157 25925 26191 25959
rect 28549 25925 28583 25959
rect 17141 25857 17175 25891
rect 17233 25857 17267 25891
rect 17417 25857 17451 25891
rect 18061 25857 18095 25891
rect 18337 25857 18371 25891
rect 18429 25857 18463 25891
rect 18889 25857 18923 25891
rect 19073 25857 19107 25891
rect 19165 25857 19199 25891
rect 21465 25857 21499 25891
rect 22201 25857 22235 25891
rect 22468 25857 22502 25891
rect 23673 25857 23707 25891
rect 25246 25857 25280 25891
rect 25513 25857 25547 25891
rect 25605 25857 25639 25891
rect 25697 25857 25731 25891
rect 26249 25857 26283 25891
rect 26525 25857 26559 25891
rect 26801 25857 26835 25891
rect 26985 25857 27019 25891
rect 27353 25857 27387 25891
rect 27905 25857 27939 25891
rect 28641 25857 28675 25891
rect 28825 25857 28859 25891
rect 29561 25857 29595 25891
rect 29653 25857 29687 25891
rect 29929 25857 29963 25891
rect 30205 25857 30239 25891
rect 30297 25857 30331 25891
rect 30573 25857 30607 25891
rect 30941 25857 30975 25891
rect 31033 25857 31067 25891
rect 31217 25857 31251 25891
rect 31401 25857 31435 25891
rect 31493 25857 31527 25891
rect 32413 25857 32447 25891
rect 18153 25789 18187 25823
rect 27261 25789 27295 25823
rect 27997 25789 28031 25823
rect 29837 25789 29871 25823
rect 32321 25789 32355 25823
rect 32689 25789 32723 25823
rect 32781 25789 32815 25823
rect 17417 25721 17451 25755
rect 23949 25721 23983 25755
rect 26525 25721 26559 25755
rect 27077 25721 27111 25755
rect 30481 25721 30515 25755
rect 17693 25653 17727 25687
rect 18613 25653 18647 25687
rect 18705 25653 18739 25687
rect 23581 25653 23615 25687
rect 25881 25653 25915 25687
rect 25973 25653 26007 25687
rect 28181 25653 28215 25687
rect 28365 25653 28399 25687
rect 30021 25653 30055 25687
rect 30757 25653 30791 25687
rect 31677 25653 31711 25687
rect 32137 25653 32171 25687
rect 18061 25449 18095 25483
rect 18429 25449 18463 25483
rect 19809 25449 19843 25483
rect 22845 25449 22879 25483
rect 24685 25449 24719 25483
rect 27077 25449 27111 25483
rect 28549 25449 28583 25483
rect 29377 25449 29411 25483
rect 30021 25449 30055 25483
rect 33057 25449 33091 25483
rect 17509 25381 17543 25415
rect 19349 25381 19383 25415
rect 20637 25381 20671 25415
rect 25053 25381 25087 25415
rect 29837 25381 29871 25415
rect 23029 25313 23063 25347
rect 25145 25313 25179 25347
rect 16865 25245 16899 25279
rect 17049 25245 17083 25279
rect 17233 25245 17267 25279
rect 18245 25245 18279 25279
rect 18521 25245 18555 25279
rect 18981 25245 19015 25279
rect 19073 25245 19107 25279
rect 19533 25245 19567 25279
rect 19625 25245 19659 25279
rect 19901 25245 19935 25279
rect 19993 25245 20027 25279
rect 20177 25245 20211 25279
rect 20361 25245 20395 25279
rect 20637 25245 20671 25279
rect 22661 25245 22695 25279
rect 22845 25245 22879 25279
rect 23213 25245 23247 25279
rect 24869 25245 24903 25279
rect 25697 25245 25731 25279
rect 27169 25245 27203 25279
rect 27436 25245 27470 25279
rect 29193 25245 29227 25279
rect 29389 25245 29423 25279
rect 30205 25245 30239 25279
rect 30472 25245 30506 25279
rect 31677 25245 31711 25279
rect 17509 25177 17543 25211
rect 19349 25177 19383 25211
rect 20913 25177 20947 25211
rect 21097 25177 21131 25211
rect 25964 25177 25998 25211
rect 29561 25177 29595 25211
rect 31922 25177 31956 25211
rect 16957 25109 16991 25143
rect 17325 25109 17359 25143
rect 20085 25109 20119 25143
rect 20453 25109 20487 25143
rect 20729 25109 20763 25143
rect 23397 25109 23431 25143
rect 31585 25109 31619 25143
rect 18061 24905 18095 24939
rect 18153 24905 18187 24939
rect 19901 24905 19935 24939
rect 20545 24905 20579 24939
rect 22017 24905 22051 24939
rect 25053 24905 25087 24939
rect 25881 24905 25915 24939
rect 30021 24905 30055 24939
rect 30481 24905 30515 24939
rect 31769 24905 31803 24939
rect 16948 24837 16982 24871
rect 21465 24837 21499 24871
rect 32137 24837 32171 24871
rect 21235 24803 21269 24837
rect 16681 24769 16715 24803
rect 18337 24769 18371 24803
rect 18429 24769 18463 24803
rect 18788 24769 18822 24803
rect 20821 24769 20855 24803
rect 21833 24769 21867 24803
rect 22845 24769 22879 24803
rect 24133 24769 24167 24803
rect 24961 24769 24995 24803
rect 26065 24769 26099 24803
rect 26341 24769 26375 24803
rect 28365 24769 28399 24803
rect 28641 24769 28675 24803
rect 28908 24769 28942 24803
rect 30113 24769 30147 24803
rect 30297 24769 30331 24803
rect 30757 24769 30791 24803
rect 30849 24769 30883 24803
rect 31125 24769 31159 24803
rect 31309 24769 31343 24803
rect 31401 24769 31435 24803
rect 31493 24769 31527 24803
rect 32413 24769 32447 24803
rect 32505 24769 32539 24803
rect 32597 24769 32631 24803
rect 32873 24769 32907 24803
rect 33149 24769 33183 24803
rect 18153 24701 18187 24735
rect 18521 24701 18555 24735
rect 20269 24701 20303 24735
rect 20913 24701 20947 24735
rect 23029 24701 23063 24735
rect 26249 24701 26283 24735
rect 28181 24701 28215 24735
rect 32965 24633 32999 24667
rect 21097 24565 21131 24599
rect 21281 24565 21315 24599
rect 22661 24565 22695 24599
rect 24317 24565 24351 24599
rect 28549 24565 28583 24599
rect 31033 24565 31067 24599
rect 32689 24565 32723 24599
rect 18429 24361 18463 24395
rect 19257 24361 19291 24395
rect 21005 24361 21039 24395
rect 22385 24361 22419 24395
rect 23029 24361 23063 24395
rect 23489 24361 23523 24395
rect 29101 24361 29135 24395
rect 30021 24361 30055 24395
rect 33333 24361 33367 24395
rect 19625 24293 19659 24327
rect 22845 24293 22879 24327
rect 17049 24225 17083 24259
rect 19717 24225 19751 24259
rect 21189 24225 21223 24259
rect 31953 24225 31987 24259
rect 17316 24157 17350 24191
rect 19441 24157 19475 24191
rect 20453 24157 20487 24191
rect 20545 24157 20579 24191
rect 20637 24157 20671 24191
rect 20821 24157 20855 24191
rect 20913 24157 20947 24191
rect 22017 24157 22051 24191
rect 22201 24157 22235 24191
rect 22569 24157 22603 24191
rect 22661 24157 22695 24191
rect 22937 24157 22971 24191
rect 23213 24157 23247 24191
rect 23305 24157 23339 24191
rect 23581 24157 23615 24191
rect 23857 24157 23891 24191
rect 23949 24157 23983 24191
rect 24685 24157 24719 24191
rect 24941 24157 24975 24191
rect 29285 24157 29319 24191
rect 31217 24157 31251 24191
rect 31493 24157 31527 24191
rect 21189 24089 21223 24123
rect 22109 24089 22143 24123
rect 29929 24089 29963 24123
rect 32220 24089 32254 24123
rect 20177 24021 20211 24055
rect 24133 24021 24167 24055
rect 26065 24021 26099 24055
rect 31033 24021 31067 24055
rect 31309 24021 31343 24055
rect 21465 23817 21499 23851
rect 23213 23817 23247 23851
rect 25145 23817 25179 23851
rect 25881 23817 25915 23851
rect 26801 23817 26835 23851
rect 32597 23817 32631 23851
rect 20330 23749 20364 23783
rect 25329 23749 25363 23783
rect 26157 23749 26191 23783
rect 27230 23749 27264 23783
rect 30840 23749 30874 23783
rect 20085 23681 20119 23715
rect 21833 23681 21867 23715
rect 22100 23681 22134 23715
rect 23489 23681 23523 23715
rect 24032 23681 24066 23715
rect 25697 23681 25731 23715
rect 26525 23681 26559 23715
rect 26617 23681 26651 23715
rect 26985 23681 27019 23715
rect 29561 23681 29595 23715
rect 29653 23681 29687 23715
rect 29837 23681 29871 23715
rect 30113 23681 30147 23715
rect 30573 23681 30607 23715
rect 32321 23681 32355 23715
rect 32505 23681 32539 23715
rect 32781 23681 32815 23715
rect 23673 23613 23707 23647
rect 23765 23613 23799 23647
rect 32137 23613 32171 23647
rect 31953 23545 31987 23579
rect 23305 23477 23339 23511
rect 26341 23477 26375 23511
rect 28365 23477 28399 23511
rect 29929 23477 29963 23511
rect 22293 23273 22327 23307
rect 23029 23273 23063 23307
rect 23581 23273 23615 23307
rect 24409 23273 24443 23307
rect 25513 23273 25547 23307
rect 27537 23273 27571 23307
rect 30941 23273 30975 23307
rect 23213 23205 23247 23239
rect 23765 23205 23799 23239
rect 29285 23137 29319 23171
rect 17325 23069 17359 23103
rect 17509 23069 17543 23103
rect 20637 23069 20671 23103
rect 21741 23069 21775 23103
rect 22477 23069 22511 23103
rect 23489 23069 23523 23103
rect 24593 23069 24627 23103
rect 25421 23069 25455 23103
rect 25881 23069 25915 23103
rect 27537 23069 27571 23103
rect 27629 23069 27663 23103
rect 27813 23069 27847 23103
rect 29561 23069 29595 23103
rect 31217 23069 31251 23103
rect 20370 23001 20404 23035
rect 24041 23001 24075 23035
rect 26148 23001 26182 23035
rect 29018 23001 29052 23035
rect 29828 23001 29862 23035
rect 17417 22933 17451 22967
rect 19257 22933 19291 22967
rect 21833 22933 21867 22967
rect 27261 22933 27295 22967
rect 27353 22933 27387 22967
rect 27905 22933 27939 22967
rect 31033 22933 31067 22967
rect 18337 22729 18371 22763
rect 19158 22729 19192 22763
rect 23397 22729 23431 22763
rect 25789 22729 25823 22763
rect 26525 22729 26559 22763
rect 27537 22729 27571 22763
rect 29009 22729 29043 22763
rect 32505 22729 32539 22763
rect 17224 22661 17258 22695
rect 18889 22661 18923 22695
rect 19257 22661 19291 22695
rect 21649 22661 21683 22695
rect 24593 22661 24627 22695
rect 25513 22661 25547 22695
rect 25881 22661 25915 22695
rect 27445 22661 27479 22695
rect 29561 22661 29595 22695
rect 30748 22661 30782 22695
rect 32873 22661 32907 22695
rect 18613 22593 18647 22627
rect 18705 22593 18739 22627
rect 18981 22593 19015 22627
rect 19073 22593 19107 22627
rect 21373 22593 21407 22627
rect 22109 22593 22143 22627
rect 22201 22593 22235 22627
rect 22293 22593 22327 22627
rect 22477 22593 22511 22627
rect 23213 22593 23247 22627
rect 23765 22593 23799 22627
rect 23857 22593 23891 22627
rect 24501 22593 24535 22627
rect 24961 22593 24995 22627
rect 26157 22593 26191 22627
rect 26341 22593 26375 22627
rect 27629 22593 27663 22627
rect 27905 22593 27939 22627
rect 28089 22593 28123 22627
rect 28549 22593 28583 22627
rect 28641 22593 28675 22627
rect 28825 22593 28859 22627
rect 32413 22593 32447 22627
rect 16957 22525 16991 22559
rect 18889 22525 18923 22559
rect 21649 22525 21683 22559
rect 24777 22525 24811 22559
rect 25329 22525 25363 22559
rect 28273 22525 28307 22559
rect 30481 22525 30515 22559
rect 27261 22457 27295 22491
rect 32689 22457 32723 22491
rect 21465 22389 21499 22423
rect 21833 22389 21867 22423
rect 24041 22389 24075 22423
rect 25145 22389 25179 22423
rect 27813 22389 27847 22423
rect 28365 22389 28399 22423
rect 29837 22389 29871 22423
rect 31861 22389 31895 22423
rect 21373 22185 21407 22219
rect 26341 22185 26375 22219
rect 26709 22185 26743 22219
rect 30665 22185 30699 22219
rect 34345 22185 34379 22219
rect 19717 22049 19751 22083
rect 21741 22049 21775 22083
rect 26065 22049 26099 22083
rect 26985 22049 27019 22083
rect 27353 22049 27387 22083
rect 31677 22049 31711 22083
rect 17049 21981 17083 22015
rect 18616 21981 18650 22015
rect 18889 21981 18923 22015
rect 21649 21981 21683 22015
rect 21997 21981 22031 22015
rect 24593 21981 24627 22015
rect 26157 21981 26191 22015
rect 26617 21981 26651 22015
rect 27169 21981 27203 22015
rect 28181 21981 28215 22015
rect 29929 21981 29963 22015
rect 30389 21981 30423 22015
rect 30481 21981 30515 22015
rect 31033 21981 31067 22015
rect 31125 21981 31159 22015
rect 31217 21981 31251 22015
rect 31401 21981 31435 22015
rect 31861 21981 31895 22015
rect 32137 21981 32171 22015
rect 33793 21981 33827 22015
rect 34529 21981 34563 22015
rect 17316 21913 17350 21947
rect 18705 21913 18739 21947
rect 19984 21913 20018 21947
rect 21373 21913 21407 21947
rect 24041 21913 24075 21947
rect 25798 21913 25832 21947
rect 32045 21913 32079 21947
rect 32404 21913 32438 21947
rect 18429 21845 18463 21879
rect 19073 21845 19107 21879
rect 21097 21845 21131 21879
rect 21557 21845 21591 21879
rect 23121 21845 23155 21879
rect 23949 21845 23983 21879
rect 24409 21845 24443 21879
rect 24685 21845 24719 21879
rect 28365 21845 28399 21879
rect 30113 21845 30147 21879
rect 30757 21845 30791 21879
rect 33517 21845 33551 21879
rect 33609 21845 33643 21879
rect 17693 21641 17727 21675
rect 18321 21641 18355 21675
rect 20361 21641 20395 21675
rect 21649 21641 21683 21675
rect 22385 21641 22419 21675
rect 24593 21641 24627 21675
rect 25881 21641 25915 21675
rect 32137 21641 32171 21675
rect 33425 21641 33459 21675
rect 17417 21573 17451 21607
rect 18521 21573 18555 21607
rect 18613 21573 18647 21607
rect 19165 21573 19199 21607
rect 21281 21573 21315 21607
rect 21497 21573 21531 21607
rect 23388 21573 23422 21607
rect 25053 21573 25087 21607
rect 29570 21573 29604 21607
rect 30196 21573 30230 21607
rect 17693 21505 17727 21539
rect 18797 21505 18831 21539
rect 18889 21505 18923 21539
rect 19349 21505 19383 21539
rect 19441 21505 19475 21539
rect 19717 21505 19751 21539
rect 19901 21505 19935 21539
rect 20085 21505 20119 21539
rect 20545 21505 20579 21539
rect 20913 21505 20947 21539
rect 21097 21505 21131 21539
rect 21189 21505 21223 21539
rect 22385 21505 22419 21539
rect 22845 21505 22879 21539
rect 23029 21505 23063 21539
rect 25697 21505 25731 21539
rect 25973 21505 26007 21539
rect 26157 21505 26191 21539
rect 28098 21505 28132 21539
rect 29837 21505 29871 21539
rect 29929 21505 29963 21539
rect 32413 21505 32447 21539
rect 32873 21505 32907 21539
rect 33149 21505 33183 21539
rect 19809 21437 19843 21471
rect 20821 21437 20855 21471
rect 21833 21437 21867 21471
rect 22477 21437 22511 21471
rect 22661 21437 22695 21471
rect 23121 21437 23155 21471
rect 25605 21437 25639 21471
rect 26065 21437 26099 21471
rect 28365 21437 28399 21471
rect 32965 21437 32999 21471
rect 33241 21437 33275 21471
rect 33517 21437 33551 21471
rect 33609 21437 33643 21471
rect 17601 21369 17635 21403
rect 18613 21369 18647 21403
rect 20913 21369 20947 21403
rect 24777 21369 24811 21403
rect 25237 21369 25271 21403
rect 31309 21369 31343 21403
rect 32597 21369 32631 21403
rect 18153 21301 18187 21335
rect 18337 21301 18371 21335
rect 19625 21301 19659 21335
rect 20269 21301 20303 21335
rect 20729 21301 20763 21335
rect 21465 21301 21499 21335
rect 24501 21301 24535 21335
rect 25145 21301 25179 21335
rect 26985 21301 27019 21335
rect 28457 21301 28491 21335
rect 32505 21301 32539 21335
rect 32689 21301 32723 21335
rect 20177 21097 20211 21131
rect 20453 21097 20487 21131
rect 21925 21097 21959 21131
rect 23673 21097 23707 21131
rect 24961 21097 24995 21131
rect 27077 21097 27111 21131
rect 27537 21097 27571 21131
rect 30021 21097 30055 21131
rect 31953 21097 31987 21131
rect 33885 21097 33919 21131
rect 27721 21029 27755 21063
rect 27997 21029 28031 21063
rect 18153 20961 18187 20995
rect 24133 20961 24167 20995
rect 25053 20961 25087 20995
rect 27169 20961 27203 20995
rect 30389 20961 30423 20995
rect 17877 20893 17911 20927
rect 17969 20893 18003 20927
rect 20269 20893 20303 20927
rect 20545 20893 20579 20927
rect 21833 20893 21867 20927
rect 22017 20893 22051 20927
rect 23857 20893 23891 20927
rect 23949 20893 23983 20927
rect 24225 20893 24259 20927
rect 24685 20893 24719 20927
rect 24777 20893 24811 20927
rect 25329 20893 25363 20927
rect 25421 20893 25455 20927
rect 26433 20893 26467 20927
rect 26617 20893 26651 20927
rect 26709 20893 26743 20927
rect 26801 20893 26835 20927
rect 27445 20893 27479 20927
rect 27629 20893 27663 20927
rect 27905 20893 27939 20927
rect 29377 20893 29411 20927
rect 30205 20893 30239 20927
rect 30573 20893 30607 20927
rect 30840 20893 30874 20927
rect 32505 20893 32539 20927
rect 25145 20825 25179 20859
rect 29110 20825 29144 20859
rect 32772 20825 32806 20859
rect 18153 20757 18187 20791
rect 24501 20757 24535 20791
rect 20269 20553 20303 20587
rect 27261 20553 27295 20587
rect 27721 20553 27755 20587
rect 27813 20553 27847 20587
rect 28733 20553 28767 20587
rect 32597 20553 32631 20587
rect 33333 20553 33367 20587
rect 19809 20485 19843 20519
rect 22385 20485 22419 20519
rect 32873 20485 32907 20519
rect 17233 20417 17267 20451
rect 17417 20417 17451 20451
rect 17693 20417 17727 20451
rect 18225 20417 18259 20451
rect 19579 20417 19613 20451
rect 19717 20417 19751 20451
rect 19992 20417 20026 20451
rect 20085 20417 20119 20451
rect 20361 20417 20395 20451
rect 22569 20417 22603 20451
rect 23397 20417 23431 20451
rect 23489 20417 23523 20451
rect 23581 20417 23615 20451
rect 23765 20417 23799 20451
rect 23857 20417 23891 20451
rect 24041 20417 24075 20451
rect 26157 20417 26191 20451
rect 26341 20417 26375 20451
rect 26617 20417 26651 20451
rect 27169 20417 27203 20451
rect 27445 20417 27479 20451
rect 27905 20417 27939 20451
rect 27997 20417 28031 20451
rect 28181 20417 28215 20451
rect 28365 20417 28399 20451
rect 28549 20417 28583 20451
rect 31033 20417 31067 20451
rect 31125 20417 31159 20451
rect 31309 20417 31343 20451
rect 31585 20417 31619 20451
rect 32137 20417 32171 20451
rect 32413 20417 32447 20451
rect 33241 20417 33275 20451
rect 33517 20417 33551 20451
rect 17325 20349 17359 20383
rect 17877 20349 17911 20383
rect 17969 20349 18003 20383
rect 23949 20349 23983 20383
rect 25973 20349 26007 20383
rect 27537 20349 27571 20383
rect 32229 20349 32263 20383
rect 32689 20281 32723 20315
rect 17509 20213 17543 20247
rect 19349 20213 19383 20247
rect 19441 20213 19475 20247
rect 22753 20213 22787 20247
rect 23121 20213 23155 20247
rect 26433 20213 26467 20247
rect 26985 20213 27019 20247
rect 31401 20213 31435 20247
rect 32413 20213 32447 20247
rect 33057 20213 33091 20247
rect 18153 20009 18187 20043
rect 18521 20009 18555 20043
rect 19993 20009 20027 20043
rect 22385 20009 22419 20043
rect 24225 20009 24259 20043
rect 26801 20009 26835 20043
rect 28273 20009 28307 20043
rect 29561 20009 29595 20043
rect 33517 20009 33551 20043
rect 32413 19941 32447 19975
rect 18245 19873 18279 19907
rect 21557 19873 21591 19907
rect 21741 19873 21775 19907
rect 22201 19873 22235 19907
rect 22661 19873 22695 19907
rect 22845 19873 22879 19907
rect 30941 19873 30975 19907
rect 31033 19873 31067 19907
rect 32505 19873 32539 19907
rect 1409 19805 1443 19839
rect 17693 19805 17727 19839
rect 17969 19805 18003 19839
rect 19441 19805 19475 19839
rect 20085 19805 20119 19839
rect 21189 19805 21223 19839
rect 21465 19805 21499 19839
rect 21833 19805 21867 19839
rect 22109 19805 22143 19839
rect 22569 19805 22603 19839
rect 22753 19805 22787 19839
rect 23112 19805 23146 19839
rect 25421 19805 25455 19839
rect 25688 19805 25722 19839
rect 26893 19805 26927 19839
rect 27149 19805 27183 19839
rect 32781 19805 32815 19839
rect 33149 19805 33183 19839
rect 33333 19805 33367 19839
rect 17448 19737 17482 19771
rect 17785 19737 17819 19771
rect 18505 19737 18539 19771
rect 18705 19737 18739 19771
rect 19625 19737 19659 19771
rect 30674 19737 30708 19771
rect 31300 19737 31334 19771
rect 33057 19737 33091 19771
rect 16313 19669 16347 19703
rect 18337 19669 18371 19703
rect 19257 19669 19291 19703
rect 21005 19669 21039 19703
rect 21373 19669 21407 19703
rect 21557 19669 21591 19703
rect 32689 19669 32723 19703
rect 32873 19669 32907 19703
rect 21005 19465 21039 19499
rect 21649 19465 21683 19499
rect 23213 19465 23247 19499
rect 26341 19465 26375 19499
rect 27353 19465 27387 19499
rect 29377 19465 29411 19499
rect 30481 19465 30515 19499
rect 31953 19465 31987 19499
rect 33701 19465 33735 19499
rect 19073 19397 19107 19431
rect 22845 19397 22879 19431
rect 30818 19397 30852 19431
rect 32588 19397 32622 19431
rect 17233 19329 17267 19363
rect 17417 19329 17451 19363
rect 18889 19329 18923 19363
rect 18981 19329 19015 19363
rect 19257 19329 19291 19363
rect 19625 19329 19659 19363
rect 19892 19329 19926 19363
rect 21281 19329 21315 19363
rect 21925 19329 21959 19363
rect 22017 19329 22051 19363
rect 22201 19329 22235 19363
rect 23397 19329 23431 19363
rect 24602 19329 24636 19363
rect 24869 19329 24903 19363
rect 24961 19329 24995 19363
rect 25228 19329 25262 19363
rect 26985 19329 27019 19363
rect 27169 19329 27203 19363
rect 28273 19329 28307 19363
rect 28733 19329 28767 19363
rect 28917 19329 28951 19363
rect 29009 19329 29043 19363
rect 29101 19329 29135 19363
rect 30297 19329 30331 19363
rect 17325 19261 17359 19295
rect 21373 19261 21407 19295
rect 30573 19261 30607 19295
rect 32321 19261 32355 19295
rect 22109 19193 22143 19227
rect 18705 19125 18739 19159
rect 22385 19125 22419 19159
rect 22569 19125 22603 19159
rect 23489 19125 23523 19159
rect 28457 19125 28491 19159
rect 17969 18921 18003 18955
rect 18981 18921 19015 18955
rect 20177 18921 20211 18955
rect 21373 18921 21407 18955
rect 21741 18921 21775 18955
rect 22937 18921 22971 18955
rect 23857 18921 23891 18955
rect 28825 18921 28859 18955
rect 29561 18921 29595 18955
rect 30021 18921 30055 18955
rect 31217 18921 31251 18955
rect 32597 18921 32631 18955
rect 28733 18853 28767 18887
rect 19533 18785 19567 18819
rect 21281 18785 21315 18819
rect 21465 18785 21499 18819
rect 21557 18785 21591 18819
rect 29193 18785 29227 18819
rect 30757 18785 30791 18819
rect 31585 18785 31619 18819
rect 16129 18717 16163 18751
rect 17785 18717 17819 18751
rect 18061 18717 18095 18751
rect 19073 18717 19107 18751
rect 19257 18717 19291 18751
rect 19441 18717 19475 18751
rect 19625 18717 19659 18751
rect 19809 18717 19843 18751
rect 20453 18717 20487 18751
rect 20545 18717 20579 18751
rect 20637 18717 20671 18751
rect 20821 18717 20855 18751
rect 21189 18717 21223 18751
rect 21833 18717 21867 18751
rect 22845 18717 22879 18751
rect 23029 18717 23063 18751
rect 23213 18717 23247 18751
rect 23397 18717 23431 18751
rect 23489 18717 23523 18751
rect 23581 18717 23615 18751
rect 27261 18717 27295 18751
rect 27353 18717 27387 18751
rect 29009 18717 29043 18751
rect 29837 18717 29871 18751
rect 29929 18717 29963 18751
rect 30113 18717 30147 18751
rect 30297 18717 30331 18751
rect 30573 18717 30607 18751
rect 31401 18717 31435 18751
rect 32229 18717 32263 18751
rect 32413 18717 32447 18751
rect 16396 18649 16430 18683
rect 17601 18649 17635 18683
rect 27620 18649 27654 18683
rect 17509 18581 17543 18615
rect 19993 18581 20027 18615
rect 21557 18581 21591 18615
rect 27077 18581 27111 18615
rect 30389 18581 30423 18615
rect 17141 18377 17175 18411
rect 17995 18377 18029 18411
rect 25513 18377 25547 18411
rect 27537 18377 27571 18411
rect 29653 18377 29687 18411
rect 29745 18377 29779 18411
rect 17785 18309 17819 18343
rect 18889 18309 18923 18343
rect 17049 18241 17083 18275
rect 17233 18241 17267 18275
rect 17509 18241 17543 18275
rect 18659 18241 18693 18275
rect 18797 18241 18831 18275
rect 19072 18241 19106 18275
rect 19165 18241 19199 18275
rect 20913 18241 20947 18275
rect 22569 18241 22603 18275
rect 22753 18241 22787 18275
rect 24961 18241 24995 18275
rect 25789 18241 25823 18275
rect 25881 18241 25915 18275
rect 25973 18241 26007 18275
rect 26157 18241 26191 18275
rect 26433 18241 26467 18275
rect 26985 18241 27019 18275
rect 27721 18241 27755 18275
rect 27813 18241 27847 18275
rect 27997 18241 28031 18275
rect 28181 18241 28215 18275
rect 28540 18241 28574 18275
rect 30858 18241 30892 18275
rect 17693 18173 17727 18207
rect 26617 18173 26651 18207
rect 28273 18173 28307 18207
rect 31125 18173 31159 18207
rect 21097 18105 21131 18139
rect 17325 18037 17359 18071
rect 17969 18037 18003 18071
rect 18153 18037 18187 18071
rect 18521 18037 18555 18071
rect 22753 18037 22787 18071
rect 24777 18037 24811 18071
rect 26249 18037 26283 18071
rect 27169 18037 27203 18071
rect 17509 17833 17543 17867
rect 18061 17833 18095 17867
rect 19349 17833 19383 17867
rect 23121 17833 23155 17867
rect 23857 17833 23891 17867
rect 23949 17833 23983 17867
rect 25789 17833 25823 17867
rect 29837 17833 29871 17867
rect 20591 17765 20625 17799
rect 21189 17765 21223 17799
rect 21833 17765 21867 17799
rect 30113 17765 30147 17799
rect 15209 17697 15243 17731
rect 18337 17697 18371 17731
rect 20453 17697 20487 17731
rect 24041 17697 24075 17731
rect 15577 17629 15611 17663
rect 17325 17629 17359 17663
rect 17601 17629 17635 17663
rect 18245 17629 18279 17663
rect 18429 17629 18463 17663
rect 19441 17629 19475 17663
rect 20177 17629 20211 17663
rect 20269 17629 20303 17663
rect 20729 17629 20763 17663
rect 20821 17629 20855 17663
rect 21005 17629 21039 17663
rect 21281 17629 21315 17663
rect 21373 17629 21407 17663
rect 21557 17629 21591 17663
rect 21649 17629 21683 17663
rect 21833 17629 21867 17663
rect 22017 17629 22051 17663
rect 22201 17629 22235 17663
rect 22937 17629 22971 17663
rect 23213 17629 23247 17663
rect 23305 17629 23339 17663
rect 23489 17629 23523 17663
rect 23673 17629 23707 17663
rect 23765 17629 23799 17663
rect 24409 17629 24443 17663
rect 24676 17629 24710 17663
rect 25881 17629 25915 17663
rect 28466 17629 28500 17663
rect 28733 17629 28767 17663
rect 29653 17629 29687 17663
rect 31493 17629 31527 17663
rect 17003 17561 17037 17595
rect 17785 17561 17819 17595
rect 22109 17561 22143 17595
rect 22477 17561 22511 17595
rect 22661 17561 22695 17595
rect 26126 17561 26160 17595
rect 31226 17561 31260 17595
rect 17141 17493 17175 17527
rect 20085 17493 20119 17527
rect 20361 17493 20395 17527
rect 21465 17493 21499 17527
rect 22293 17493 22327 17527
rect 22753 17493 22787 17527
rect 27261 17493 27295 17527
rect 27353 17493 27387 17527
rect 16221 17289 16255 17323
rect 18061 17289 18095 17323
rect 20177 17289 20211 17323
rect 25053 17289 25087 17323
rect 25789 17289 25823 17323
rect 25881 17289 25915 17323
rect 26985 17289 27019 17323
rect 29285 17289 29319 17323
rect 29745 17289 29779 17323
rect 30849 17289 30883 17323
rect 16948 17221 16982 17255
rect 29837 17221 29871 17255
rect 15577 17153 15611 17187
rect 16129 17153 16163 17187
rect 16681 17153 16715 17187
rect 18153 17153 18187 17187
rect 18337 17153 18371 17187
rect 18425 17153 18459 17187
rect 18613 17153 18647 17187
rect 18797 17153 18831 17187
rect 18889 17153 18923 17187
rect 19165 17153 19199 17187
rect 19717 17153 19751 17187
rect 19809 17153 19843 17187
rect 20085 17153 20119 17187
rect 20361 17153 20395 17187
rect 20545 17153 20579 17187
rect 20637 17153 20671 17187
rect 20729 17153 20763 17187
rect 20913 17153 20947 17187
rect 21189 17153 21223 17187
rect 22017 17153 22051 17187
rect 22201 17153 22235 17187
rect 22293 17153 22327 17187
rect 22477 17153 22511 17187
rect 22753 17153 22787 17187
rect 22937 17153 22971 17187
rect 23029 17153 23063 17187
rect 23305 17153 23339 17187
rect 23489 17153 23523 17187
rect 24694 17153 24728 17187
rect 24961 17153 24995 17187
rect 25237 17153 25271 17187
rect 25605 17153 25639 17187
rect 26157 17153 26191 17187
rect 26617 17153 26651 17187
rect 27169 17153 27203 17187
rect 27261 17153 27295 17187
rect 29469 17153 29503 17187
rect 30665 17153 30699 17187
rect 18981 17085 19015 17119
rect 19993 17085 20027 17119
rect 21281 17085 21315 17119
rect 21649 17085 21683 17119
rect 23121 17085 23155 17119
rect 25421 17085 25455 17119
rect 26341 17085 26375 17119
rect 29561 17085 29595 17119
rect 29929 17085 29963 17119
rect 21005 17017 21039 17051
rect 22385 17017 22419 17051
rect 23581 17017 23615 17051
rect 26249 17017 26283 17051
rect 18153 16949 18187 16983
rect 19349 16949 19383 16983
rect 19533 16949 19567 16983
rect 26433 16949 26467 16983
rect 18889 16745 18923 16779
rect 19533 16745 19567 16779
rect 20729 16745 20763 16779
rect 21741 16745 21775 16779
rect 22293 16745 22327 16779
rect 22569 16745 22603 16779
rect 22937 16745 22971 16779
rect 23397 16745 23431 16779
rect 25881 16745 25915 16779
rect 29377 16745 29411 16779
rect 30113 16745 30147 16779
rect 20913 16677 20947 16711
rect 22661 16677 22695 16711
rect 30573 16677 30607 16711
rect 17509 16609 17543 16643
rect 19625 16609 19659 16643
rect 20545 16609 20579 16643
rect 22109 16609 22143 16643
rect 22477 16609 22511 16643
rect 23765 16609 23799 16643
rect 26065 16609 26099 16643
rect 26157 16609 26191 16643
rect 26433 16609 26467 16643
rect 29561 16609 29595 16643
rect 19257 16541 19291 16575
rect 19809 16541 19843 16575
rect 19993 16541 20027 16575
rect 20453 16541 20487 16575
rect 21097 16541 21131 16575
rect 21189 16541 21223 16575
rect 21373 16541 21407 16575
rect 21557 16541 21591 16575
rect 22017 16541 22051 16575
rect 22753 16541 22787 16575
rect 22845 16541 22879 16575
rect 23029 16541 23063 16575
rect 23167 16541 23201 16575
rect 23305 16541 23339 16575
rect 23581 16541 23615 16575
rect 26525 16541 26559 16575
rect 26617 16541 26651 16575
rect 28273 16541 28307 16575
rect 29101 16541 29135 16575
rect 29193 16541 29227 16575
rect 29745 16541 29779 16575
rect 29837 16541 29871 16575
rect 30205 16541 30239 16575
rect 30389 16541 30423 16575
rect 30757 16541 30791 16575
rect 17776 16473 17810 16507
rect 19717 16473 19751 16507
rect 29377 16473 29411 16507
rect 31024 16473 31058 16507
rect 19349 16405 19383 16439
rect 19901 16405 19935 16439
rect 26249 16405 26283 16439
rect 26801 16405 26835 16439
rect 28457 16405 28491 16439
rect 28917 16405 28951 16439
rect 29929 16405 29963 16439
rect 32137 16405 32171 16439
rect 20361 16201 20395 16235
rect 25881 16201 25915 16235
rect 26157 16201 26191 16235
rect 26985 16201 27019 16235
rect 29837 16201 29871 16235
rect 31309 16201 31343 16235
rect 17877 16133 17911 16167
rect 19064 16133 19098 16167
rect 28098 16133 28132 16167
rect 28702 16133 28736 16167
rect 18061 16065 18095 16099
rect 18337 16065 18371 16099
rect 20453 16065 20487 16099
rect 24685 16065 24719 16099
rect 25145 16065 25179 16099
rect 25789 16065 25823 16099
rect 25973 16065 26007 16099
rect 26617 16065 26651 16099
rect 26801 16065 26835 16099
rect 28365 16065 28399 16099
rect 28457 16065 28491 16099
rect 30185 16065 30219 16099
rect 31585 16065 31619 16099
rect 31677 16065 31711 16099
rect 18797 15997 18831 16031
rect 24869 15997 24903 16031
rect 25329 15997 25363 16031
rect 26433 15997 26467 16031
rect 29929 15997 29963 16031
rect 18245 15929 18279 15963
rect 20177 15929 20211 15963
rect 25605 15929 25639 15963
rect 24501 15861 24535 15895
rect 24961 15861 24995 15895
rect 31401 15861 31435 15895
rect 25881 15657 25915 15691
rect 28365 15657 28399 15691
rect 29745 15657 29779 15691
rect 30021 15657 30055 15691
rect 31493 15657 31527 15691
rect 28825 15521 28859 15555
rect 24041 15453 24075 15487
rect 24409 15453 24443 15487
rect 27261 15453 27295 15487
rect 28181 15453 28215 15487
rect 28549 15453 28583 15487
rect 28733 15453 28767 15487
rect 29009 15453 29043 15487
rect 29193 15453 29227 15487
rect 29561 15453 29595 15487
rect 31401 15453 31435 15487
rect 31677 15453 31711 15487
rect 24676 15385 24710 15419
rect 26994 15385 27028 15419
rect 31134 15385 31168 15419
rect 24225 15317 24259 15351
rect 25789 15317 25823 15351
rect 27997 15317 28031 15351
rect 21189 15113 21223 15147
rect 25881 15113 25915 15147
rect 26433 15113 26467 15147
rect 26709 15113 26743 15147
rect 29009 15113 29043 15147
rect 30021 15113 30055 15147
rect 31677 15113 31711 15147
rect 24746 15045 24780 15079
rect 25973 15045 26007 15079
rect 27896 15045 27930 15079
rect 19809 14977 19843 15011
rect 20076 14977 20110 15011
rect 23029 14977 23063 15011
rect 23296 14977 23330 15011
rect 26157 14977 26191 15011
rect 26249 14977 26283 15011
rect 26525 14977 26559 15011
rect 27629 14977 27663 15011
rect 29837 14977 29871 15011
rect 31493 14977 31527 15011
rect 24501 14909 24535 14943
rect 31309 14909 31343 14943
rect 24409 14773 24443 14807
rect 25973 14773 26007 14807
rect 23397 14569 23431 14603
rect 24593 14569 24627 14603
rect 26157 14569 26191 14603
rect 28273 14569 28307 14603
rect 22477 14433 22511 14467
rect 25789 14433 25823 14467
rect 22661 14365 22695 14399
rect 22845 14365 22879 14399
rect 23213 14365 23247 14399
rect 24409 14365 24443 14399
rect 25973 14365 26007 14399
rect 27905 14365 27939 14399
rect 28089 14365 28123 14399
rect 33977 12189 34011 12223
rect 34161 12053 34195 12087
rect 34161 11713 34195 11747
rect 34437 11577 34471 11611
rect 1409 10013 1443 10047
rect 28457 2601 28491 2635
rect 34345 2601 34379 2635
rect 1685 2465 1719 2499
rect 1409 2397 1443 2431
rect 9137 2397 9171 2431
rect 19625 2397 19659 2431
rect 28641 2397 28675 2431
rect 34529 2397 34563 2431
rect 19349 2261 19383 2295
<< metal1 >>
rect 1104 39738 34868 39760
rect 1104 39686 5170 39738
rect 5222 39686 5234 39738
rect 5286 39686 5298 39738
rect 5350 39686 5362 39738
rect 5414 39686 5426 39738
rect 5478 39686 13611 39738
rect 13663 39686 13675 39738
rect 13727 39686 13739 39738
rect 13791 39686 13803 39738
rect 13855 39686 13867 39738
rect 13919 39686 22052 39738
rect 22104 39686 22116 39738
rect 22168 39686 22180 39738
rect 22232 39686 22244 39738
rect 22296 39686 22308 39738
rect 22360 39686 30493 39738
rect 30545 39686 30557 39738
rect 30609 39686 30621 39738
rect 30673 39686 30685 39738
rect 30737 39686 30749 39738
rect 30801 39686 34868 39738
rect 1104 39664 34868 39686
rect 26418 39584 26424 39636
rect 26476 39624 26482 39636
rect 26513 39627 26571 39633
rect 26513 39624 26525 39627
rect 26476 39596 26525 39624
rect 26476 39584 26482 39596
rect 26513 39593 26525 39596
rect 26559 39593 26571 39627
rect 26513 39587 26571 39593
rect 34425 39627 34483 39633
rect 34425 39593 34437 39627
rect 34471 39624 34483 39627
rect 35434 39624 35440 39636
rect 34471 39596 35440 39624
rect 34471 39593 34483 39596
rect 34425 39587 34483 39593
rect 35434 39584 35440 39596
rect 35492 39584 35498 39636
rect 934 39380 940 39432
rect 992 39420 998 39432
rect 1397 39423 1455 39429
rect 1397 39420 1409 39423
rect 992 39392 1409 39420
rect 992 39380 998 39392
rect 1397 39389 1409 39392
rect 1443 39389 1455 39423
rect 1397 39383 1455 39389
rect 7098 39380 7104 39432
rect 7156 39420 7162 39432
rect 7193 39423 7251 39429
rect 7193 39420 7205 39423
rect 7156 39392 7205 39420
rect 7156 39380 7162 39392
rect 7193 39389 7205 39392
rect 7239 39389 7251 39423
rect 7193 39383 7251 39389
rect 16758 39380 16764 39432
rect 16816 39420 16822 39432
rect 16853 39423 16911 39429
rect 16853 39420 16865 39423
rect 16816 39392 16865 39420
rect 16816 39380 16822 39392
rect 16853 39389 16865 39392
rect 16899 39389 16911 39423
rect 16853 39383 16911 39389
rect 34146 39312 34152 39364
rect 34204 39312 34210 39364
rect 1578 39244 1584 39296
rect 1636 39244 1642 39296
rect 7377 39287 7435 39293
rect 7377 39253 7389 39287
rect 7423 39284 7435 39287
rect 16114 39284 16120 39296
rect 7423 39256 16120 39284
rect 7423 39253 7435 39256
rect 7377 39247 7435 39253
rect 16114 39244 16120 39256
rect 16172 39244 16178 39296
rect 17037 39287 17095 39293
rect 17037 39253 17049 39287
rect 17083 39284 17095 39287
rect 17586 39284 17592 39296
rect 17083 39256 17592 39284
rect 17083 39253 17095 39256
rect 17037 39247 17095 39253
rect 17586 39244 17592 39256
rect 17644 39244 17650 39296
rect 1104 39194 35027 39216
rect 1104 39142 9390 39194
rect 9442 39142 9454 39194
rect 9506 39142 9518 39194
rect 9570 39142 9582 39194
rect 9634 39142 9646 39194
rect 9698 39142 17831 39194
rect 17883 39142 17895 39194
rect 17947 39142 17959 39194
rect 18011 39142 18023 39194
rect 18075 39142 18087 39194
rect 18139 39142 26272 39194
rect 26324 39142 26336 39194
rect 26388 39142 26400 39194
rect 26452 39142 26464 39194
rect 26516 39142 26528 39194
rect 26580 39142 34713 39194
rect 34765 39142 34777 39194
rect 34829 39142 34841 39194
rect 34893 39142 34905 39194
rect 34957 39142 34969 39194
rect 35021 39142 35027 39194
rect 1104 39120 35027 39142
rect 1104 38650 34868 38672
rect 1104 38598 5170 38650
rect 5222 38598 5234 38650
rect 5286 38598 5298 38650
rect 5350 38598 5362 38650
rect 5414 38598 5426 38650
rect 5478 38598 13611 38650
rect 13663 38598 13675 38650
rect 13727 38598 13739 38650
rect 13791 38598 13803 38650
rect 13855 38598 13867 38650
rect 13919 38598 22052 38650
rect 22104 38598 22116 38650
rect 22168 38598 22180 38650
rect 22232 38598 22244 38650
rect 22296 38598 22308 38650
rect 22360 38598 30493 38650
rect 30545 38598 30557 38650
rect 30609 38598 30621 38650
rect 30673 38598 30685 38650
rect 30737 38598 30749 38650
rect 30801 38598 34868 38650
rect 1104 38576 34868 38598
rect 1104 38106 35027 38128
rect 1104 38054 9390 38106
rect 9442 38054 9454 38106
rect 9506 38054 9518 38106
rect 9570 38054 9582 38106
rect 9634 38054 9646 38106
rect 9698 38054 17831 38106
rect 17883 38054 17895 38106
rect 17947 38054 17959 38106
rect 18011 38054 18023 38106
rect 18075 38054 18087 38106
rect 18139 38054 26272 38106
rect 26324 38054 26336 38106
rect 26388 38054 26400 38106
rect 26452 38054 26464 38106
rect 26516 38054 26528 38106
rect 26580 38054 34713 38106
rect 34765 38054 34777 38106
rect 34829 38054 34841 38106
rect 34893 38054 34905 38106
rect 34957 38054 34969 38106
rect 35021 38054 35027 38106
rect 1104 38032 35027 38054
rect 1104 37562 34868 37584
rect 1104 37510 5170 37562
rect 5222 37510 5234 37562
rect 5286 37510 5298 37562
rect 5350 37510 5362 37562
rect 5414 37510 5426 37562
rect 5478 37510 13611 37562
rect 13663 37510 13675 37562
rect 13727 37510 13739 37562
rect 13791 37510 13803 37562
rect 13855 37510 13867 37562
rect 13919 37510 22052 37562
rect 22104 37510 22116 37562
rect 22168 37510 22180 37562
rect 22232 37510 22244 37562
rect 22296 37510 22308 37562
rect 22360 37510 30493 37562
rect 30545 37510 30557 37562
rect 30609 37510 30621 37562
rect 30673 37510 30685 37562
rect 30737 37510 30749 37562
rect 30801 37510 34868 37562
rect 1104 37488 34868 37510
rect 1104 37018 35027 37040
rect 1104 36966 9390 37018
rect 9442 36966 9454 37018
rect 9506 36966 9518 37018
rect 9570 36966 9582 37018
rect 9634 36966 9646 37018
rect 9698 36966 17831 37018
rect 17883 36966 17895 37018
rect 17947 36966 17959 37018
rect 18011 36966 18023 37018
rect 18075 36966 18087 37018
rect 18139 36966 26272 37018
rect 26324 36966 26336 37018
rect 26388 36966 26400 37018
rect 26452 36966 26464 37018
rect 26516 36966 26528 37018
rect 26580 36966 34713 37018
rect 34765 36966 34777 37018
rect 34829 36966 34841 37018
rect 34893 36966 34905 37018
rect 34957 36966 34969 37018
rect 35021 36966 35027 37018
rect 1104 36944 35027 36966
rect 1104 36474 34868 36496
rect 1104 36422 5170 36474
rect 5222 36422 5234 36474
rect 5286 36422 5298 36474
rect 5350 36422 5362 36474
rect 5414 36422 5426 36474
rect 5478 36422 13611 36474
rect 13663 36422 13675 36474
rect 13727 36422 13739 36474
rect 13791 36422 13803 36474
rect 13855 36422 13867 36474
rect 13919 36422 22052 36474
rect 22104 36422 22116 36474
rect 22168 36422 22180 36474
rect 22232 36422 22244 36474
rect 22296 36422 22308 36474
rect 22360 36422 30493 36474
rect 30545 36422 30557 36474
rect 30609 36422 30621 36474
rect 30673 36422 30685 36474
rect 30737 36422 30749 36474
rect 30801 36422 34868 36474
rect 1104 36400 34868 36422
rect 1104 35930 35027 35952
rect 1104 35878 9390 35930
rect 9442 35878 9454 35930
rect 9506 35878 9518 35930
rect 9570 35878 9582 35930
rect 9634 35878 9646 35930
rect 9698 35878 17831 35930
rect 17883 35878 17895 35930
rect 17947 35878 17959 35930
rect 18011 35878 18023 35930
rect 18075 35878 18087 35930
rect 18139 35878 26272 35930
rect 26324 35878 26336 35930
rect 26388 35878 26400 35930
rect 26452 35878 26464 35930
rect 26516 35878 26528 35930
rect 26580 35878 34713 35930
rect 34765 35878 34777 35930
rect 34829 35878 34841 35930
rect 34893 35878 34905 35930
rect 34957 35878 34969 35930
rect 35021 35878 35027 35930
rect 1104 35856 35027 35878
rect 1104 35386 34868 35408
rect 1104 35334 5170 35386
rect 5222 35334 5234 35386
rect 5286 35334 5298 35386
rect 5350 35334 5362 35386
rect 5414 35334 5426 35386
rect 5478 35334 13611 35386
rect 13663 35334 13675 35386
rect 13727 35334 13739 35386
rect 13791 35334 13803 35386
rect 13855 35334 13867 35386
rect 13919 35334 22052 35386
rect 22104 35334 22116 35386
rect 22168 35334 22180 35386
rect 22232 35334 22244 35386
rect 22296 35334 22308 35386
rect 22360 35334 30493 35386
rect 30545 35334 30557 35386
rect 30609 35334 30621 35386
rect 30673 35334 30685 35386
rect 30737 35334 30749 35386
rect 30801 35334 34868 35386
rect 1104 35312 34868 35334
rect 1104 34842 35027 34864
rect 1104 34790 9390 34842
rect 9442 34790 9454 34842
rect 9506 34790 9518 34842
rect 9570 34790 9582 34842
rect 9634 34790 9646 34842
rect 9698 34790 17831 34842
rect 17883 34790 17895 34842
rect 17947 34790 17959 34842
rect 18011 34790 18023 34842
rect 18075 34790 18087 34842
rect 18139 34790 26272 34842
rect 26324 34790 26336 34842
rect 26388 34790 26400 34842
rect 26452 34790 26464 34842
rect 26516 34790 26528 34842
rect 26580 34790 34713 34842
rect 34765 34790 34777 34842
rect 34829 34790 34841 34842
rect 34893 34790 34905 34842
rect 34957 34790 34969 34842
rect 35021 34790 35027 34842
rect 1104 34768 35027 34790
rect 1104 34298 34868 34320
rect 1104 34246 5170 34298
rect 5222 34246 5234 34298
rect 5286 34246 5298 34298
rect 5350 34246 5362 34298
rect 5414 34246 5426 34298
rect 5478 34246 13611 34298
rect 13663 34246 13675 34298
rect 13727 34246 13739 34298
rect 13791 34246 13803 34298
rect 13855 34246 13867 34298
rect 13919 34246 22052 34298
rect 22104 34246 22116 34298
rect 22168 34246 22180 34298
rect 22232 34246 22244 34298
rect 22296 34246 22308 34298
rect 22360 34246 30493 34298
rect 30545 34246 30557 34298
rect 30609 34246 30621 34298
rect 30673 34246 30685 34298
rect 30737 34246 30749 34298
rect 30801 34246 34868 34298
rect 1104 34224 34868 34246
rect 25958 33940 25964 33992
rect 26016 33980 26022 33992
rect 26329 33983 26387 33989
rect 26329 33980 26341 33983
rect 26016 33952 26341 33980
rect 26016 33940 26022 33952
rect 26329 33949 26341 33952
rect 26375 33949 26387 33983
rect 26329 33943 26387 33949
rect 26513 33983 26571 33989
rect 26513 33949 26525 33983
rect 26559 33949 26571 33983
rect 26513 33943 26571 33949
rect 26528 33912 26556 33943
rect 26878 33912 26884 33924
rect 26160 33884 26884 33912
rect 26160 33856 26188 33884
rect 26878 33872 26884 33884
rect 26936 33872 26942 33924
rect 26142 33804 26148 33856
rect 26200 33804 26206 33856
rect 26421 33847 26479 33853
rect 26421 33813 26433 33847
rect 26467 33844 26479 33847
rect 26786 33844 26792 33856
rect 26467 33816 26792 33844
rect 26467 33813 26479 33816
rect 26421 33807 26479 33813
rect 26786 33804 26792 33816
rect 26844 33804 26850 33856
rect 1104 33754 35027 33776
rect 1104 33702 9390 33754
rect 9442 33702 9454 33754
rect 9506 33702 9518 33754
rect 9570 33702 9582 33754
rect 9634 33702 9646 33754
rect 9698 33702 17831 33754
rect 17883 33702 17895 33754
rect 17947 33702 17959 33754
rect 18011 33702 18023 33754
rect 18075 33702 18087 33754
rect 18139 33702 26272 33754
rect 26324 33702 26336 33754
rect 26388 33702 26400 33754
rect 26452 33702 26464 33754
rect 26516 33702 26528 33754
rect 26580 33702 34713 33754
rect 34765 33702 34777 33754
rect 34829 33702 34841 33754
rect 34893 33702 34905 33754
rect 34957 33702 34969 33754
rect 35021 33702 35027 33754
rect 1104 33680 35027 33702
rect 26786 33600 26792 33652
rect 26844 33600 26850 33652
rect 26804 33572 26832 33600
rect 27157 33575 27215 33581
rect 27157 33572 27169 33575
rect 26804 33544 27169 33572
rect 27157 33541 27169 33544
rect 27203 33541 27215 33575
rect 27157 33535 27215 33541
rect 30576 33544 32260 33572
rect 1578 33464 1584 33516
rect 1636 33504 1642 33516
rect 23109 33507 23167 33513
rect 23109 33504 23121 33507
rect 1636 33476 23121 33504
rect 1636 33464 1642 33476
rect 23109 33473 23121 33476
rect 23155 33473 23167 33507
rect 23109 33467 23167 33473
rect 23934 33464 23940 33516
rect 23992 33464 23998 33516
rect 25498 33464 25504 33516
rect 25556 33504 25562 33516
rect 25869 33507 25927 33513
rect 25869 33504 25881 33507
rect 25556 33476 25881 33504
rect 25556 33464 25562 33476
rect 25869 33473 25881 33476
rect 25915 33473 25927 33507
rect 25869 33467 25927 33473
rect 26329 33507 26387 33513
rect 26329 33473 26341 33507
rect 26375 33504 26387 33507
rect 26789 33507 26847 33513
rect 26375 33476 26740 33504
rect 26375 33473 26387 33476
rect 26329 33467 26387 33473
rect 22925 33439 22983 33445
rect 22925 33405 22937 33439
rect 22971 33436 22983 33439
rect 23842 33436 23848 33448
rect 22971 33408 23848 33436
rect 22971 33405 22983 33408
rect 22925 33399 22983 33405
rect 23842 33396 23848 33408
rect 23900 33396 23906 33448
rect 25961 33439 26019 33445
rect 25961 33405 25973 33439
rect 26007 33436 26019 33439
rect 26142 33436 26148 33448
rect 26007 33408 26148 33436
rect 26007 33405 26019 33408
rect 25961 33399 26019 33405
rect 26142 33396 26148 33408
rect 26200 33396 26206 33448
rect 26421 33439 26479 33445
rect 26421 33405 26433 33439
rect 26467 33436 26479 33439
rect 26602 33436 26608 33448
rect 26467 33408 26608 33436
rect 26467 33405 26479 33408
rect 26421 33399 26479 33405
rect 26602 33396 26608 33408
rect 26660 33396 26666 33448
rect 26712 33436 26740 33476
rect 26789 33473 26801 33507
rect 26835 33504 26847 33507
rect 26970 33504 26976 33516
rect 26835 33476 26976 33504
rect 26835 33473 26847 33476
rect 26789 33467 26847 33473
rect 26970 33464 26976 33476
rect 27028 33464 27034 33516
rect 28620 33507 28678 33513
rect 28620 33473 28632 33507
rect 28666 33504 28678 33507
rect 29546 33504 29552 33516
rect 28666 33476 29552 33504
rect 28666 33473 28678 33476
rect 28620 33467 28678 33473
rect 29546 33464 29552 33476
rect 29604 33464 29610 33516
rect 29825 33507 29883 33513
rect 29825 33473 29837 33507
rect 29871 33473 29883 33507
rect 29825 33467 29883 33473
rect 30101 33507 30159 33513
rect 30101 33473 30113 33507
rect 30147 33504 30159 33507
rect 30190 33504 30196 33516
rect 30147 33476 30196 33504
rect 30147 33473 30159 33476
rect 30101 33467 30159 33473
rect 27062 33436 27068 33448
rect 26712 33408 27068 33436
rect 27062 33396 27068 33408
rect 27120 33396 27126 33448
rect 27246 33396 27252 33448
rect 27304 33436 27310 33448
rect 28350 33436 28356 33448
rect 27304 33408 28356 33436
rect 27304 33396 27310 33408
rect 28350 33396 28356 33408
rect 28408 33396 28414 33448
rect 26234 33328 26240 33380
rect 26292 33368 26298 33380
rect 26513 33371 26571 33377
rect 26513 33368 26525 33371
rect 26292 33340 26525 33368
rect 26292 33328 26298 33340
rect 26513 33337 26525 33340
rect 26559 33337 26571 33371
rect 27430 33368 27436 33380
rect 26513 33331 26571 33337
rect 27080 33340 27436 33368
rect 23293 33303 23351 33309
rect 23293 33269 23305 33303
rect 23339 33300 23351 33303
rect 23474 33300 23480 33312
rect 23339 33272 23480 33300
rect 23339 33269 23351 33272
rect 23293 33263 23351 33269
rect 23474 33260 23480 33272
rect 23532 33260 23538 33312
rect 24121 33303 24179 33309
rect 24121 33269 24133 33303
rect 24167 33300 24179 33303
rect 24486 33300 24492 33312
rect 24167 33272 24492 33300
rect 24167 33269 24179 33272
rect 24121 33263 24179 33269
rect 24486 33260 24492 33272
rect 24544 33260 24550 33312
rect 26326 33260 26332 33312
rect 26384 33300 26390 33312
rect 26651 33303 26709 33309
rect 26651 33300 26663 33303
rect 26384 33272 26663 33300
rect 26384 33260 26390 33272
rect 26651 33269 26663 33272
rect 26697 33300 26709 33303
rect 27080 33300 27108 33340
rect 27430 33328 27436 33340
rect 27488 33328 27494 33380
rect 29733 33371 29791 33377
rect 29733 33337 29745 33371
rect 29779 33368 29791 33371
rect 29840 33368 29868 33467
rect 30190 33464 30196 33476
rect 30248 33464 30254 33516
rect 30282 33464 30288 33516
rect 30340 33504 30346 33516
rect 30576 33513 30604 33544
rect 32232 33516 32260 33544
rect 30561 33507 30619 33513
rect 30561 33504 30573 33507
rect 30340 33476 30573 33504
rect 30340 33464 30346 33476
rect 30561 33473 30573 33476
rect 30607 33473 30619 33507
rect 30561 33467 30619 33473
rect 31018 33464 31024 33516
rect 31076 33464 31082 33516
rect 32214 33464 32220 33516
rect 32272 33464 32278 33516
rect 30006 33396 30012 33448
rect 30064 33396 30070 33448
rect 30377 33439 30435 33445
rect 30377 33436 30389 33439
rect 30116 33408 30389 33436
rect 30116 33368 30144 33408
rect 30377 33405 30389 33408
rect 30423 33405 30435 33439
rect 30377 33399 30435 33405
rect 29779 33340 30144 33368
rect 29779 33337 29791 33340
rect 29733 33331 29791 33337
rect 30116 33312 30144 33340
rect 30745 33371 30803 33377
rect 30745 33337 30757 33371
rect 30791 33368 30803 33371
rect 31294 33368 31300 33380
rect 30791 33340 31300 33368
rect 30791 33337 30803 33340
rect 30745 33331 30803 33337
rect 31294 33328 31300 33340
rect 31352 33328 31358 33380
rect 26697 33272 27108 33300
rect 26697 33269 26709 33272
rect 26651 33263 26709 33269
rect 27154 33260 27160 33312
rect 27212 33300 27218 33312
rect 27341 33303 27399 33309
rect 27341 33300 27353 33303
rect 27212 33272 27353 33300
rect 27212 33260 27218 33272
rect 27341 33269 27353 33272
rect 27387 33269 27399 33303
rect 27341 33263 27399 33269
rect 29914 33260 29920 33312
rect 29972 33260 29978 33312
rect 30098 33260 30104 33312
rect 30156 33260 30162 33312
rect 30285 33303 30343 33309
rect 30285 33269 30297 33303
rect 30331 33300 30343 33303
rect 30374 33300 30380 33312
rect 30331 33272 30380 33300
rect 30331 33269 30343 33272
rect 30285 33263 30343 33269
rect 30374 33260 30380 33272
rect 30432 33260 30438 33312
rect 30834 33260 30840 33312
rect 30892 33260 30898 33312
rect 1104 33210 34868 33232
rect 1104 33158 5170 33210
rect 5222 33158 5234 33210
rect 5286 33158 5298 33210
rect 5350 33158 5362 33210
rect 5414 33158 5426 33210
rect 5478 33158 13611 33210
rect 13663 33158 13675 33210
rect 13727 33158 13739 33210
rect 13791 33158 13803 33210
rect 13855 33158 13867 33210
rect 13919 33158 22052 33210
rect 22104 33158 22116 33210
rect 22168 33158 22180 33210
rect 22232 33158 22244 33210
rect 22296 33158 22308 33210
rect 22360 33158 30493 33210
rect 30545 33158 30557 33210
rect 30609 33158 30621 33210
rect 30673 33158 30685 33210
rect 30737 33158 30749 33210
rect 30801 33158 34868 33210
rect 1104 33136 34868 33158
rect 23934 33056 23940 33108
rect 23992 33096 23998 33108
rect 24213 33099 24271 33105
rect 24213 33096 24225 33099
rect 23992 33068 24225 33096
rect 23992 33056 23998 33068
rect 24213 33065 24225 33068
rect 24259 33065 24271 33099
rect 24213 33059 24271 33065
rect 25590 33056 25596 33108
rect 25648 33096 25654 33108
rect 27246 33096 27252 33108
rect 25648 33068 27252 33096
rect 25648 33056 25654 33068
rect 27246 33056 27252 33068
rect 27304 33056 27310 33108
rect 29546 33056 29552 33108
rect 29604 33056 29610 33108
rect 26142 32988 26148 33040
rect 26200 32988 26206 33040
rect 26970 33028 26976 33040
rect 26344 33000 26976 33028
rect 23382 32920 23388 32972
rect 23440 32960 23446 32972
rect 24397 32963 24455 32969
rect 24397 32960 24409 32963
rect 23440 32932 24409 32960
rect 23440 32920 23446 32932
rect 24397 32929 24409 32932
rect 24443 32929 24455 32963
rect 24397 32923 24455 32929
rect 23474 32852 23480 32904
rect 23532 32892 23538 32904
rect 23569 32895 23627 32901
rect 23569 32892 23581 32895
rect 23532 32864 23581 32892
rect 23532 32852 23538 32864
rect 23569 32861 23581 32864
rect 23615 32861 23627 32895
rect 23569 32855 23627 32861
rect 23934 32852 23940 32904
rect 23992 32852 23998 32904
rect 24029 32895 24087 32901
rect 24029 32861 24041 32895
rect 24075 32892 24087 32895
rect 24302 32892 24308 32904
rect 24075 32864 24308 32892
rect 24075 32861 24087 32864
rect 24029 32855 24087 32861
rect 24302 32852 24308 32864
rect 24360 32852 24366 32904
rect 24486 32852 24492 32904
rect 24544 32892 24550 32904
rect 24653 32895 24711 32901
rect 24653 32892 24665 32895
rect 24544 32864 24665 32892
rect 24544 32852 24550 32864
rect 24653 32861 24665 32864
rect 24699 32861 24711 32895
rect 24653 32855 24711 32861
rect 26053 32895 26111 32901
rect 26053 32861 26065 32895
rect 26099 32892 26111 32895
rect 26160 32892 26188 32988
rect 26344 32969 26372 33000
rect 26970 32988 26976 33000
rect 27028 32988 27034 33040
rect 26329 32963 26387 32969
rect 26329 32929 26341 32963
rect 26375 32929 26387 32963
rect 26329 32923 26387 32929
rect 26697 32963 26755 32969
rect 26697 32929 26709 32963
rect 26743 32960 26755 32963
rect 27154 32960 27160 32972
rect 26743 32932 27160 32960
rect 26743 32929 26755 32932
rect 26697 32923 26755 32929
rect 27154 32920 27160 32932
rect 27212 32920 27218 32972
rect 27264 32969 27292 33056
rect 28629 33031 28687 33037
rect 28629 32997 28641 33031
rect 28675 33028 28687 33031
rect 28675 33000 28764 33028
rect 28675 32997 28687 33000
rect 28629 32991 28687 32997
rect 28736 32969 28764 33000
rect 27249 32963 27307 32969
rect 27249 32929 27261 32963
rect 27295 32929 27307 32963
rect 27249 32923 27307 32929
rect 28721 32963 28779 32969
rect 28721 32929 28733 32963
rect 28767 32960 28779 32963
rect 28767 32932 29960 32960
rect 28767 32929 28779 32932
rect 28721 32923 28779 32929
rect 29932 32904 29960 32932
rect 26099 32864 26188 32892
rect 26099 32861 26111 32864
rect 26053 32855 26111 32861
rect 26234 32852 26240 32904
rect 26292 32852 26298 32904
rect 26605 32895 26663 32901
rect 26605 32861 26617 32895
rect 26651 32892 26663 32895
rect 27338 32892 27344 32904
rect 26651 32864 27344 32892
rect 26651 32861 26663 32864
rect 26605 32855 26663 32861
rect 27338 32852 27344 32864
rect 27396 32852 27402 32904
rect 28905 32895 28963 32901
rect 28905 32861 28917 32895
rect 28951 32861 28963 32895
rect 28905 32855 28963 32861
rect 29089 32895 29147 32901
rect 29089 32861 29101 32895
rect 29135 32892 29147 32895
rect 29365 32895 29423 32901
rect 29365 32892 29377 32895
rect 29135 32864 29377 32892
rect 29135 32861 29147 32864
rect 29089 32855 29147 32861
rect 29365 32861 29377 32864
rect 29411 32861 29423 32895
rect 29365 32855 29423 32861
rect 27494 32827 27552 32833
rect 27494 32824 27506 32827
rect 23768 32796 27506 32824
rect 23768 32765 23796 32796
rect 27494 32793 27506 32796
rect 27540 32793 27552 32827
rect 27494 32787 27552 32793
rect 28920 32824 28948 32855
rect 29730 32852 29736 32904
rect 29788 32852 29794 32904
rect 29914 32852 29920 32904
rect 29972 32852 29978 32904
rect 31202 32852 31208 32904
rect 31260 32852 31266 32904
rect 31294 32852 31300 32904
rect 31352 32892 31358 32904
rect 31481 32895 31539 32901
rect 31481 32892 31493 32895
rect 31352 32864 31493 32892
rect 31352 32852 31358 32864
rect 31481 32861 31493 32864
rect 31527 32861 31539 32895
rect 31481 32855 31539 32861
rect 30282 32824 30288 32836
rect 28920 32796 30288 32824
rect 28920 32768 28948 32796
rect 30282 32784 30288 32796
rect 30340 32784 30346 32836
rect 30960 32827 31018 32833
rect 30960 32793 30972 32827
rect 31006 32824 31018 32827
rect 31006 32796 31340 32824
rect 31006 32793 31018 32796
rect 30960 32787 31018 32793
rect 23753 32759 23811 32765
rect 23753 32725 23765 32759
rect 23799 32725 23811 32759
rect 23753 32719 23811 32725
rect 25682 32716 25688 32768
rect 25740 32756 25746 32768
rect 25777 32759 25835 32765
rect 25777 32756 25789 32759
rect 25740 32728 25789 32756
rect 25740 32716 25746 32728
rect 25777 32725 25789 32728
rect 25823 32725 25835 32759
rect 25777 32719 25835 32725
rect 25866 32716 25872 32768
rect 25924 32716 25930 32768
rect 26142 32716 26148 32768
rect 26200 32756 26206 32768
rect 26421 32759 26479 32765
rect 26421 32756 26433 32759
rect 26200 32728 26433 32756
rect 26200 32716 26206 32728
rect 26421 32725 26433 32728
rect 26467 32725 26479 32759
rect 26421 32719 26479 32725
rect 27062 32716 27068 32768
rect 27120 32716 27126 32768
rect 28902 32716 28908 32768
rect 28960 32716 28966 32768
rect 29086 32716 29092 32768
rect 29144 32756 29150 32768
rect 29181 32759 29239 32765
rect 29181 32756 29193 32759
rect 29144 32728 29193 32756
rect 29144 32716 29150 32728
rect 29181 32725 29193 32728
rect 29227 32725 29239 32759
rect 29181 32719 29239 32725
rect 29825 32759 29883 32765
rect 29825 32725 29837 32759
rect 29871 32756 29883 32759
rect 30006 32756 30012 32768
rect 29871 32728 30012 32756
rect 29871 32725 29883 32728
rect 29825 32719 29883 32725
rect 30006 32716 30012 32728
rect 30064 32716 30070 32768
rect 31312 32765 31340 32796
rect 31297 32759 31355 32765
rect 31297 32725 31309 32759
rect 31343 32725 31355 32759
rect 31297 32719 31355 32725
rect 1104 32666 35027 32688
rect 1104 32614 9390 32666
rect 9442 32614 9454 32666
rect 9506 32614 9518 32666
rect 9570 32614 9582 32666
rect 9634 32614 9646 32666
rect 9698 32614 17831 32666
rect 17883 32614 17895 32666
rect 17947 32614 17959 32666
rect 18011 32614 18023 32666
rect 18075 32614 18087 32666
rect 18139 32614 26272 32666
rect 26324 32614 26336 32666
rect 26388 32614 26400 32666
rect 26452 32614 26464 32666
rect 26516 32614 26528 32666
rect 26580 32614 34713 32666
rect 34765 32614 34777 32666
rect 34829 32614 34841 32666
rect 34893 32614 34905 32666
rect 34957 32614 34969 32666
rect 35021 32614 35027 32666
rect 1104 32592 35027 32614
rect 25774 32552 25780 32564
rect 25444 32524 25780 32552
rect 17589 32419 17647 32425
rect 17589 32385 17601 32419
rect 17635 32416 17647 32419
rect 18322 32416 18328 32428
rect 17635 32388 18328 32416
rect 17635 32385 17647 32388
rect 17589 32379 17647 32385
rect 18322 32376 18328 32388
rect 18380 32376 18386 32428
rect 18690 32425 18696 32428
rect 18684 32379 18696 32425
rect 18690 32376 18696 32379
rect 18748 32376 18754 32428
rect 20257 32419 20315 32425
rect 20257 32385 20269 32419
rect 20303 32416 20315 32419
rect 20530 32416 20536 32428
rect 20303 32388 20536 32416
rect 20303 32385 20315 32388
rect 20257 32379 20315 32385
rect 20530 32376 20536 32388
rect 20588 32376 20594 32428
rect 20640 32388 20944 32416
rect 17865 32351 17923 32357
rect 17865 32317 17877 32351
rect 17911 32348 17923 32351
rect 18138 32348 18144 32360
rect 17911 32320 18144 32348
rect 17911 32317 17923 32320
rect 17865 32311 17923 32317
rect 18138 32308 18144 32320
rect 18196 32308 18202 32360
rect 18417 32351 18475 32357
rect 18417 32317 18429 32351
rect 18463 32317 18475 32351
rect 18417 32311 18475 32317
rect 20073 32351 20131 32357
rect 20073 32317 20085 32351
rect 20119 32348 20131 32351
rect 20640 32348 20668 32388
rect 20119 32320 20668 32348
rect 20119 32317 20131 32320
rect 20073 32311 20131 32317
rect 17126 32240 17132 32292
rect 17184 32280 17190 32292
rect 18432 32280 18460 32311
rect 17184 32252 18460 32280
rect 17184 32240 17190 32252
rect 19794 32240 19800 32292
rect 19852 32280 19858 32292
rect 20088 32280 20116 32311
rect 20714 32308 20720 32360
rect 20772 32348 20778 32360
rect 20916 32348 20944 32388
rect 20990 32376 20996 32428
rect 21048 32376 21054 32428
rect 21726 32376 21732 32428
rect 21784 32416 21790 32428
rect 22934 32419 22992 32425
rect 22934 32416 22946 32419
rect 21784 32388 22946 32416
rect 21784 32376 21790 32388
rect 22934 32385 22946 32388
rect 22980 32385 22992 32419
rect 22934 32379 22992 32385
rect 23201 32419 23259 32425
rect 23201 32385 23213 32419
rect 23247 32416 23259 32419
rect 23382 32416 23388 32428
rect 23247 32388 23388 32416
rect 23247 32385 23259 32388
rect 23201 32379 23259 32385
rect 23382 32376 23388 32388
rect 23440 32376 23446 32428
rect 25444 32425 25472 32524
rect 25774 32512 25780 32524
rect 25832 32512 25838 32564
rect 25866 32512 25872 32564
rect 25924 32512 25930 32564
rect 25958 32512 25964 32564
rect 26016 32552 26022 32564
rect 26016 32524 26832 32552
rect 26016 32512 26022 32524
rect 25590 32444 25596 32496
rect 25648 32484 25654 32496
rect 25884 32484 25912 32512
rect 26602 32484 26608 32496
rect 25648 32456 25721 32484
rect 25884 32456 26004 32484
rect 25648 32444 25654 32456
rect 25693 32425 25721 32456
rect 25976 32425 26004 32456
rect 26068 32456 26608 32484
rect 26068 32425 26096 32456
rect 26602 32444 26608 32456
rect 26660 32444 26666 32496
rect 26804 32425 26832 32524
rect 26970 32512 26976 32564
rect 27028 32512 27034 32564
rect 27154 32512 27160 32564
rect 27212 32552 27218 32564
rect 27212 32524 27384 32552
rect 27212 32512 27218 32524
rect 26878 32444 26884 32496
rect 26936 32444 26942 32496
rect 27356 32484 27384 32524
rect 27430 32512 27436 32564
rect 27488 32552 27494 32564
rect 27525 32555 27583 32561
rect 27525 32552 27537 32555
rect 27488 32524 27537 32552
rect 27488 32512 27494 32524
rect 27525 32521 27537 32524
rect 27571 32521 27583 32555
rect 27525 32515 27583 32521
rect 28350 32512 28356 32564
rect 28408 32552 28414 32564
rect 28408 32524 29316 32552
rect 28408 32512 28414 32524
rect 27356 32456 27660 32484
rect 25429 32419 25487 32425
rect 25429 32385 25441 32419
rect 25475 32385 25487 32419
rect 25429 32379 25487 32385
rect 25685 32419 25743 32425
rect 25685 32385 25697 32419
rect 25731 32385 25743 32419
rect 25685 32379 25743 32385
rect 25777 32419 25835 32425
rect 25777 32385 25789 32419
rect 25823 32416 25835 32419
rect 25961 32419 26019 32425
rect 25823 32388 25912 32416
rect 25823 32385 25835 32388
rect 25777 32379 25835 32385
rect 25884 32360 25912 32388
rect 25961 32385 25973 32419
rect 26007 32385 26019 32419
rect 25961 32379 26019 32385
rect 26053 32419 26111 32425
rect 26053 32385 26065 32419
rect 26099 32385 26111 32419
rect 26053 32379 26111 32385
rect 26329 32419 26387 32425
rect 26329 32385 26341 32419
rect 26375 32416 26387 32419
rect 26789 32419 26847 32425
rect 26375 32388 26740 32416
rect 26375 32385 26387 32388
rect 26329 32379 26387 32385
rect 20772 32320 20852 32348
rect 20916 32320 21956 32348
rect 20772 32308 20778 32320
rect 19852 32252 20116 32280
rect 19852 32240 19858 32252
rect 20438 32240 20444 32292
rect 20496 32280 20502 32292
rect 20824 32280 20852 32320
rect 20496 32252 20852 32280
rect 20496 32240 20502 32252
rect 21928 32224 21956 32320
rect 25866 32308 25872 32360
rect 25924 32308 25930 32360
rect 26145 32351 26203 32357
rect 26145 32317 26157 32351
rect 26191 32348 26203 32351
rect 26234 32348 26240 32360
rect 26191 32320 26240 32348
rect 26191 32317 26203 32320
rect 26145 32311 26203 32317
rect 26234 32308 26240 32320
rect 26292 32308 26298 32360
rect 25774 32240 25780 32292
rect 25832 32280 25838 32292
rect 26513 32283 26571 32289
rect 26513 32280 26525 32283
rect 25832 32252 26525 32280
rect 25832 32240 25838 32252
rect 26513 32249 26525 32252
rect 26559 32249 26571 32283
rect 26712 32280 26740 32388
rect 26789 32385 26801 32419
rect 26835 32385 26847 32419
rect 26896 32416 26924 32444
rect 27154 32417 27212 32423
rect 26896 32414 27117 32416
rect 27154 32414 27166 32417
rect 26896 32388 27166 32414
rect 27089 32386 27166 32388
rect 26789 32379 26847 32385
rect 27154 32383 27166 32386
rect 27200 32383 27212 32417
rect 26804 32348 26832 32379
rect 27154 32377 27212 32383
rect 27430 32376 27436 32428
rect 27488 32376 27494 32428
rect 27632 32425 27660 32456
rect 27617 32419 27675 32425
rect 27617 32385 27629 32419
rect 27663 32385 27675 32419
rect 27617 32379 27675 32385
rect 29086 32376 29092 32428
rect 29144 32425 29150 32428
rect 29144 32419 29167 32425
rect 29155 32385 29167 32419
rect 29288 32416 29316 32524
rect 29914 32512 29920 32564
rect 29972 32512 29978 32564
rect 30098 32512 30104 32564
rect 30156 32512 30162 32564
rect 29454 32444 29460 32496
rect 29512 32484 29518 32496
rect 29733 32487 29791 32493
rect 29733 32484 29745 32487
rect 29512 32456 29745 32484
rect 29512 32444 29518 32456
rect 29733 32453 29745 32456
rect 29779 32484 29791 32487
rect 30190 32484 30196 32496
rect 29779 32456 30196 32484
rect 29779 32453 29791 32456
rect 29733 32447 29791 32453
rect 30190 32444 30196 32456
rect 30248 32444 30254 32496
rect 30736 32487 30794 32493
rect 30736 32453 30748 32487
rect 30782 32484 30794 32487
rect 30834 32484 30840 32496
rect 30782 32456 30840 32484
rect 30782 32453 30794 32456
rect 30736 32447 30794 32453
rect 30834 32444 30840 32456
rect 30892 32444 30898 32496
rect 29365 32419 29423 32425
rect 29365 32416 29377 32419
rect 29288 32388 29377 32416
rect 29144 32379 29167 32385
rect 29365 32385 29377 32388
rect 29411 32385 29423 32419
rect 29365 32379 29423 32385
rect 29144 32376 29150 32379
rect 27341 32351 27399 32357
rect 27341 32348 27353 32351
rect 26804 32320 27353 32348
rect 27341 32317 27353 32320
rect 27387 32317 27399 32351
rect 29380 32348 29408 32379
rect 30006 32376 30012 32428
rect 30064 32376 30070 32428
rect 31202 32416 31208 32428
rect 30484 32388 31208 32416
rect 30484 32357 30512 32388
rect 31202 32376 31208 32388
rect 31260 32376 31266 32428
rect 34517 32419 34575 32425
rect 34517 32385 34529 32419
rect 34563 32416 34575 32419
rect 34882 32416 34888 32428
rect 34563 32388 34888 32416
rect 34563 32385 34575 32388
rect 34517 32379 34575 32385
rect 34882 32376 34888 32388
rect 34940 32376 34946 32428
rect 30469 32351 30527 32357
rect 30469 32348 30481 32351
rect 29380 32320 30481 32348
rect 27341 32311 27399 32317
rect 30469 32317 30481 32320
rect 30515 32317 30527 32351
rect 30469 32311 30527 32317
rect 26513 32243 26571 32249
rect 26620 32252 26740 32280
rect 17310 32172 17316 32224
rect 17368 32212 17374 32224
rect 17405 32215 17463 32221
rect 17405 32212 17417 32215
rect 17368 32184 17417 32212
rect 17368 32172 17374 32184
rect 17405 32181 17417 32184
rect 17451 32181 17463 32215
rect 17405 32175 17463 32181
rect 17770 32172 17776 32224
rect 17828 32172 17834 32224
rect 20622 32172 20628 32224
rect 20680 32212 20686 32224
rect 20809 32215 20867 32221
rect 20809 32212 20821 32215
rect 20680 32184 20821 32212
rect 20680 32172 20686 32184
rect 20809 32181 20821 32184
rect 20855 32181 20867 32215
rect 20809 32175 20867 32181
rect 21174 32172 21180 32224
rect 21232 32172 21238 32224
rect 21818 32172 21824 32224
rect 21876 32172 21882 32224
rect 21910 32172 21916 32224
rect 21968 32172 21974 32224
rect 24305 32215 24363 32221
rect 24305 32181 24317 32215
rect 24351 32212 24363 32215
rect 25498 32212 25504 32224
rect 24351 32184 25504 32212
rect 24351 32181 24363 32184
rect 24305 32175 24363 32181
rect 25498 32172 25504 32184
rect 25556 32212 25562 32224
rect 26620 32212 26648 32252
rect 29454 32240 29460 32292
rect 29512 32240 29518 32292
rect 25556 32184 26648 32212
rect 25556 32172 25562 32184
rect 26694 32172 26700 32224
rect 26752 32172 26758 32224
rect 27985 32215 28043 32221
rect 27985 32181 27997 32215
rect 28031 32212 28043 32215
rect 29472 32212 29500 32240
rect 28031 32184 29500 32212
rect 30285 32215 30343 32221
rect 28031 32181 28043 32184
rect 27985 32175 28043 32181
rect 30285 32181 30297 32215
rect 30331 32212 30343 32215
rect 31110 32212 31116 32224
rect 30331 32184 31116 32212
rect 30331 32181 30343 32184
rect 30285 32175 30343 32181
rect 31110 32172 31116 32184
rect 31168 32172 31174 32224
rect 31386 32172 31392 32224
rect 31444 32212 31450 32224
rect 31849 32215 31907 32221
rect 31849 32212 31861 32215
rect 31444 32184 31861 32212
rect 31444 32172 31450 32184
rect 31849 32181 31861 32184
rect 31895 32181 31907 32215
rect 31849 32175 31907 32181
rect 32030 32172 32036 32224
rect 32088 32212 32094 32224
rect 34333 32215 34391 32221
rect 34333 32212 34345 32215
rect 32088 32184 34345 32212
rect 32088 32172 32094 32184
rect 34333 32181 34345 32184
rect 34379 32181 34391 32215
rect 34333 32175 34391 32181
rect 1104 32122 34868 32144
rect 1104 32070 5170 32122
rect 5222 32070 5234 32122
rect 5286 32070 5298 32122
rect 5350 32070 5362 32122
rect 5414 32070 5426 32122
rect 5478 32070 13611 32122
rect 13663 32070 13675 32122
rect 13727 32070 13739 32122
rect 13791 32070 13803 32122
rect 13855 32070 13867 32122
rect 13919 32070 22052 32122
rect 22104 32070 22116 32122
rect 22168 32070 22180 32122
rect 22232 32070 22244 32122
rect 22296 32070 22308 32122
rect 22360 32070 30493 32122
rect 30545 32070 30557 32122
rect 30609 32070 30621 32122
rect 30673 32070 30685 32122
rect 30737 32070 30749 32122
rect 30801 32070 34868 32122
rect 1104 32048 34868 32070
rect 18138 31968 18144 32020
rect 18196 32008 18202 32020
rect 18417 32011 18475 32017
rect 18417 32008 18429 32011
rect 18196 31980 18429 32008
rect 18196 31968 18202 31980
rect 18417 31977 18429 31980
rect 18463 31977 18475 32011
rect 18417 31971 18475 31977
rect 18690 31968 18696 32020
rect 18748 32008 18754 32020
rect 18969 32011 19027 32017
rect 18969 32008 18981 32011
rect 18748 31980 18981 32008
rect 18748 31968 18754 31980
rect 18969 31977 18981 31980
rect 19015 31977 19027 32011
rect 18969 31971 19027 31977
rect 19794 31968 19800 32020
rect 19852 31968 19858 32020
rect 20438 31968 20444 32020
rect 20496 31968 20502 32020
rect 20717 32011 20775 32017
rect 20717 31977 20729 32011
rect 20763 32008 20775 32011
rect 20990 32008 20996 32020
rect 20763 31980 20996 32008
rect 20763 31977 20775 31980
rect 20717 31971 20775 31977
rect 20990 31968 20996 31980
rect 21048 31968 21054 32020
rect 21174 31968 21180 32020
rect 21232 31968 21238 32020
rect 21726 31968 21732 32020
rect 21784 31968 21790 32020
rect 24302 31968 24308 32020
rect 24360 32008 24366 32020
rect 26145 32011 26203 32017
rect 26145 32008 26157 32011
rect 24360 31980 26157 32008
rect 24360 31968 24366 31980
rect 26145 31977 26157 31980
rect 26191 31977 26203 32011
rect 26145 31971 26203 31977
rect 26237 32011 26295 32017
rect 26237 31977 26249 32011
rect 26283 32008 26295 32011
rect 27062 32008 27068 32020
rect 26283 31980 27068 32008
rect 26283 31977 26295 31980
rect 26237 31971 26295 31977
rect 27062 31968 27068 31980
rect 27120 32008 27126 32020
rect 29089 32011 29147 32017
rect 27120 31980 27660 32008
rect 27120 31968 27126 31980
rect 16666 31764 16672 31816
rect 16724 31804 16730 31816
rect 17037 31807 17095 31813
rect 17037 31804 17049 31807
rect 16724 31776 17049 31804
rect 16724 31764 16730 31776
rect 17037 31773 17049 31776
rect 17083 31804 17095 31807
rect 17126 31804 17132 31816
rect 17083 31776 17132 31804
rect 17083 31773 17095 31776
rect 17037 31767 17095 31773
rect 17126 31764 17132 31776
rect 17184 31764 17190 31816
rect 17310 31813 17316 31816
rect 17304 31804 17316 31813
rect 17271 31776 17316 31804
rect 17304 31767 17316 31776
rect 17310 31764 17316 31767
rect 17368 31764 17374 31816
rect 18506 31764 18512 31816
rect 18564 31804 18570 31816
rect 18785 31807 18843 31813
rect 18785 31804 18797 31807
rect 18564 31776 18797 31804
rect 18564 31764 18570 31776
rect 18785 31773 18797 31776
rect 18831 31773 18843 31807
rect 18785 31767 18843 31773
rect 18966 31764 18972 31816
rect 19024 31764 19030 31816
rect 19613 31807 19671 31813
rect 19613 31773 19625 31807
rect 19659 31804 19671 31807
rect 19812 31804 19840 31968
rect 19889 31875 19947 31881
rect 19889 31841 19901 31875
rect 19935 31872 19947 31875
rect 19935 31844 20208 31872
rect 19935 31841 19947 31844
rect 19889 31835 19947 31841
rect 20180 31816 20208 31844
rect 19659 31776 19840 31804
rect 19981 31807 20039 31813
rect 19659 31773 19671 31776
rect 19613 31767 19671 31773
rect 19981 31773 19993 31807
rect 20027 31773 20039 31807
rect 19981 31767 20039 31773
rect 19794 31736 19800 31748
rect 16684 31708 19800 31736
rect 16684 31680 16712 31708
rect 19794 31696 19800 31708
rect 19852 31696 19858 31748
rect 16666 31628 16672 31680
rect 16724 31628 16730 31680
rect 19518 31628 19524 31680
rect 19576 31628 19582 31680
rect 19702 31628 19708 31680
rect 19760 31628 19766 31680
rect 19996 31668 20024 31767
rect 20162 31764 20168 31816
rect 20220 31764 20226 31816
rect 20456 31813 20484 31968
rect 20622 31949 20628 31952
rect 20579 31943 20628 31949
rect 20579 31909 20591 31943
rect 20625 31909 20628 31943
rect 20579 31903 20628 31909
rect 20622 31900 20628 31903
rect 20680 31900 20686 31952
rect 20809 31943 20867 31949
rect 20809 31909 20821 31943
rect 20855 31940 20867 31943
rect 20855 31912 21128 31940
rect 20855 31909 20867 31912
rect 20809 31903 20867 31909
rect 20732 31844 20944 31872
rect 20441 31807 20499 31813
rect 20441 31773 20453 31807
rect 20487 31773 20499 31807
rect 20441 31767 20499 31773
rect 20732 31736 20760 31844
rect 20916 31816 20944 31844
rect 20898 31764 20904 31816
rect 20956 31764 20962 31816
rect 20993 31807 21051 31813
rect 20993 31773 21005 31807
rect 21039 31773 21051 31807
rect 20993 31767 21051 31773
rect 20364 31708 20760 31736
rect 20364 31680 20392 31708
rect 20254 31668 20260 31680
rect 19996 31640 20260 31668
rect 20254 31628 20260 31640
rect 20312 31628 20318 31680
rect 20346 31628 20352 31680
rect 20404 31628 20410 31680
rect 20806 31628 20812 31680
rect 20864 31668 20870 31680
rect 21008 31668 21036 31767
rect 21100 31736 21128 31912
rect 21192 31813 21220 31968
rect 21818 31900 21824 31952
rect 21876 31900 21882 31952
rect 25961 31943 26019 31949
rect 25961 31909 25973 31943
rect 26007 31940 26019 31943
rect 26050 31940 26056 31952
rect 26007 31912 26056 31940
rect 26007 31909 26019 31912
rect 25961 31903 26019 31909
rect 26050 31900 26056 31912
rect 26108 31900 26114 31952
rect 21836 31872 21864 31900
rect 27632 31884 27660 31980
rect 29089 31977 29101 32011
rect 29135 32008 29147 32011
rect 29730 32008 29736 32020
rect 29135 31980 29736 32008
rect 29135 31977 29147 31980
rect 29089 31971 29147 31977
rect 29730 31968 29736 31980
rect 29788 31968 29794 32020
rect 31018 31968 31024 32020
rect 31076 32008 31082 32020
rect 31113 32011 31171 32017
rect 31113 32008 31125 32011
rect 31076 31980 31125 32008
rect 31076 31968 31082 31980
rect 31113 31977 31125 31980
rect 31159 31977 31171 32011
rect 31386 32008 31392 32020
rect 31113 31971 31171 31977
rect 31312 31980 31392 32008
rect 25866 31872 25872 31884
rect 21560 31844 21864 31872
rect 22112 31844 25872 31872
rect 21560 31816 21588 31844
rect 21450 31813 21456 31816
rect 21177 31807 21235 31813
rect 21177 31773 21189 31807
rect 21223 31773 21235 31807
rect 21177 31767 21235 31773
rect 21269 31807 21327 31813
rect 21269 31773 21281 31807
rect 21315 31804 21327 31807
rect 21407 31807 21456 31813
rect 21315 31776 21349 31804
rect 21315 31773 21327 31776
rect 21269 31767 21327 31773
rect 21407 31773 21419 31807
rect 21453 31773 21456 31807
rect 21407 31767 21456 31773
rect 21284 31736 21312 31767
rect 21450 31764 21456 31767
rect 21508 31764 21514 31816
rect 21542 31764 21548 31816
rect 21600 31764 21606 31816
rect 21818 31764 21824 31816
rect 21876 31764 21882 31816
rect 21910 31764 21916 31816
rect 21968 31804 21974 31816
rect 22005 31807 22063 31813
rect 22005 31804 22017 31807
rect 21968 31776 22017 31804
rect 21968 31764 21974 31776
rect 22005 31773 22017 31776
rect 22051 31773 22063 31807
rect 22005 31767 22063 31773
rect 22112 31736 22140 31844
rect 25866 31832 25872 31844
rect 25924 31832 25930 31884
rect 26142 31832 26148 31884
rect 26200 31832 26206 31884
rect 26694 31832 26700 31884
rect 26752 31832 26758 31884
rect 27614 31832 27620 31884
rect 27672 31832 27678 31884
rect 28721 31875 28779 31881
rect 28721 31841 28733 31875
rect 28767 31872 28779 31875
rect 29454 31872 29460 31884
rect 28767 31844 29460 31872
rect 28767 31841 28779 31844
rect 28721 31835 28779 31841
rect 29454 31832 29460 31844
rect 29512 31832 29518 31884
rect 30006 31832 30012 31884
rect 30064 31872 30070 31884
rect 30745 31875 30803 31881
rect 30745 31872 30757 31875
rect 30064 31844 30757 31872
rect 30064 31832 30070 31844
rect 30745 31841 30757 31844
rect 30791 31841 30803 31875
rect 31312 31872 31340 31980
rect 31386 31968 31392 31980
rect 31444 31968 31450 32020
rect 31662 31872 31668 31884
rect 30745 31835 30803 31841
rect 30852 31844 31340 31872
rect 31404 31844 31668 31872
rect 23934 31764 23940 31816
rect 23992 31804 23998 31816
rect 26329 31807 26387 31813
rect 23992 31776 26280 31804
rect 23992 31764 23998 31776
rect 21100 31708 21312 31736
rect 21376 31708 22140 31736
rect 26252 31736 26280 31776
rect 26329 31773 26341 31807
rect 26375 31804 26387 31807
rect 26712 31804 26740 31832
rect 28902 31804 28908 31816
rect 26375 31776 26740 31804
rect 26804 31776 28908 31804
rect 26375 31773 26387 31776
rect 26329 31767 26387 31773
rect 26804 31736 26832 31776
rect 28902 31764 28908 31776
rect 28960 31764 28966 31816
rect 30469 31807 30527 31813
rect 30469 31773 30481 31807
rect 30515 31804 30527 31807
rect 30653 31807 30711 31813
rect 30515 31776 30604 31804
rect 30515 31773 30527 31776
rect 30469 31767 30527 31773
rect 26252 31708 26832 31736
rect 30576 31736 30604 31776
rect 30653 31773 30665 31807
rect 30699 31804 30711 31807
rect 30852 31804 30880 31844
rect 30699 31776 30880 31804
rect 30929 31807 30987 31813
rect 30699 31773 30711 31776
rect 30653 31767 30711 31773
rect 30929 31773 30941 31807
rect 30975 31804 30987 31807
rect 31202 31804 31208 31816
rect 30975 31776 31208 31804
rect 30975 31773 30987 31776
rect 30929 31767 30987 31773
rect 30944 31736 30972 31767
rect 31202 31764 31208 31776
rect 31260 31804 31266 31816
rect 31404 31813 31432 31844
rect 31662 31832 31668 31844
rect 31720 31832 31726 31884
rect 32214 31832 32220 31884
rect 32272 31832 32278 31884
rect 31389 31807 31447 31813
rect 31260 31776 31340 31804
rect 31260 31764 31266 31776
rect 30576 31708 30972 31736
rect 31312 31736 31340 31776
rect 31389 31773 31401 31807
rect 31435 31773 31447 31807
rect 31573 31807 31631 31813
rect 31573 31804 31585 31807
rect 31389 31767 31447 31773
rect 31496 31776 31585 31804
rect 31496 31736 31524 31776
rect 31573 31773 31585 31776
rect 31619 31773 31631 31807
rect 31573 31767 31631 31773
rect 31846 31764 31852 31816
rect 31904 31764 31910 31816
rect 32030 31764 32036 31816
rect 32088 31813 32094 31816
rect 32088 31807 32105 31813
rect 32093 31773 32105 31807
rect 32088 31767 32105 31773
rect 32088 31764 32094 31767
rect 31312 31708 31524 31736
rect 21376 31668 21404 31708
rect 20864 31640 21404 31668
rect 20864 31628 20870 31640
rect 21910 31628 21916 31680
rect 21968 31628 21974 31680
rect 30282 31628 30288 31680
rect 30340 31628 30346 31680
rect 31757 31671 31815 31677
rect 31757 31637 31769 31671
rect 31803 31668 31815 31671
rect 32122 31668 32128 31680
rect 31803 31640 32128 31668
rect 31803 31637 31815 31640
rect 31757 31631 31815 31637
rect 32122 31628 32128 31640
rect 32180 31628 32186 31680
rect 1104 31578 35027 31600
rect 1104 31526 9390 31578
rect 9442 31526 9454 31578
rect 9506 31526 9518 31578
rect 9570 31526 9582 31578
rect 9634 31526 9646 31578
rect 9698 31526 17831 31578
rect 17883 31526 17895 31578
rect 17947 31526 17959 31578
rect 18011 31526 18023 31578
rect 18075 31526 18087 31578
rect 18139 31526 26272 31578
rect 26324 31526 26336 31578
rect 26388 31526 26400 31578
rect 26452 31526 26464 31578
rect 26516 31526 26528 31578
rect 26580 31526 34713 31578
rect 34765 31526 34777 31578
rect 34829 31526 34841 31578
rect 34893 31526 34905 31578
rect 34957 31526 34969 31578
rect 35021 31526 35027 31578
rect 1104 31504 35027 31526
rect 18230 31424 18236 31476
rect 18288 31464 18294 31476
rect 18874 31464 18880 31476
rect 18288 31436 18880 31464
rect 18288 31424 18294 31436
rect 18874 31424 18880 31436
rect 18932 31424 18938 31476
rect 18966 31424 18972 31476
rect 19024 31464 19030 31476
rect 19245 31467 19303 31473
rect 19245 31464 19257 31467
rect 19024 31436 19257 31464
rect 19024 31424 19030 31436
rect 19245 31433 19257 31436
rect 19291 31433 19303 31467
rect 19245 31427 19303 31433
rect 20257 31467 20315 31473
rect 20257 31433 20269 31467
rect 20303 31464 20315 31467
rect 20622 31464 20628 31476
rect 20303 31436 20628 31464
rect 20303 31433 20315 31436
rect 20257 31427 20315 31433
rect 17678 31356 17684 31408
rect 17736 31396 17742 31408
rect 20272 31396 20300 31427
rect 20622 31424 20628 31436
rect 20680 31424 20686 31476
rect 20990 31424 20996 31476
rect 21048 31424 21054 31476
rect 23109 31467 23167 31473
rect 23109 31433 23121 31467
rect 23155 31464 23167 31467
rect 23382 31464 23388 31476
rect 23155 31436 23388 31464
rect 23155 31433 23167 31436
rect 23109 31427 23167 31433
rect 23382 31424 23388 31436
rect 23440 31424 23446 31476
rect 30282 31424 30288 31476
rect 30340 31424 30346 31476
rect 31297 31467 31355 31473
rect 31297 31464 31309 31467
rect 30668 31436 31309 31464
rect 20438 31396 20444 31408
rect 17736 31368 18184 31396
rect 17736 31356 17742 31368
rect 16758 31288 16764 31340
rect 16816 31328 16822 31340
rect 18156 31337 18184 31368
rect 19444 31368 20300 31396
rect 20364 31368 20444 31396
rect 16925 31331 16983 31337
rect 16925 31328 16937 31331
rect 16816 31300 16937 31328
rect 16816 31288 16822 31300
rect 16925 31297 16937 31300
rect 16971 31297 16983 31331
rect 16925 31291 16983 31297
rect 18141 31331 18199 31337
rect 18141 31297 18153 31331
rect 18187 31297 18199 31331
rect 18141 31291 18199 31297
rect 18414 31288 18420 31340
rect 18472 31288 18478 31340
rect 19444 31337 19472 31368
rect 19429 31331 19487 31337
rect 19429 31297 19441 31331
rect 19475 31297 19487 31331
rect 19429 31291 19487 31297
rect 19521 31331 19579 31337
rect 19521 31297 19533 31331
rect 19567 31328 19579 31331
rect 19702 31328 19708 31340
rect 19567 31300 19708 31328
rect 19567 31297 19579 31300
rect 19521 31291 19579 31297
rect 19702 31288 19708 31300
rect 19760 31288 19766 31340
rect 19797 31331 19855 31337
rect 19797 31297 19809 31331
rect 19843 31297 19855 31331
rect 19797 31291 19855 31297
rect 20073 31331 20131 31337
rect 20073 31297 20085 31331
rect 20119 31297 20131 31331
rect 20073 31291 20131 31297
rect 16666 31220 16672 31272
rect 16724 31220 16730 31272
rect 18322 31220 18328 31272
rect 18380 31260 18386 31272
rect 19812 31260 19840 31291
rect 18380 31232 18460 31260
rect 18380 31220 18386 31232
rect 18432 31201 18460 31232
rect 19536 31232 19840 31260
rect 20088 31260 20116 31291
rect 20162 31288 20168 31340
rect 20220 31288 20226 31340
rect 20254 31288 20260 31340
rect 20312 31328 20318 31340
rect 20364 31337 20392 31368
rect 20438 31356 20444 31368
rect 20496 31356 20502 31408
rect 20714 31356 20720 31408
rect 20772 31396 20778 31408
rect 21085 31399 21143 31405
rect 21085 31396 21097 31399
rect 20772 31368 21097 31396
rect 20772 31356 20778 31368
rect 21085 31365 21097 31368
rect 21131 31365 21143 31399
rect 21085 31359 21143 31365
rect 21269 31399 21327 31405
rect 21269 31365 21281 31399
rect 21315 31396 21327 31399
rect 21910 31396 21916 31408
rect 21315 31368 21916 31396
rect 21315 31365 21327 31368
rect 21269 31359 21327 31365
rect 21910 31356 21916 31368
rect 21968 31356 21974 31408
rect 24486 31356 24492 31408
rect 24544 31396 24550 31408
rect 24544 31368 25268 31396
rect 24544 31356 24550 31368
rect 20349 31331 20407 31337
rect 20349 31328 20361 31331
rect 20312 31300 20361 31328
rect 20312 31288 20318 31300
rect 20349 31297 20361 31300
rect 20395 31297 20407 31331
rect 20349 31291 20407 31297
rect 20625 31331 20683 31337
rect 20625 31297 20637 31331
rect 20671 31328 20683 31331
rect 21542 31328 21548 31340
rect 20671 31300 21548 31328
rect 20671 31297 20683 31300
rect 20625 31291 20683 31297
rect 20640 31260 20668 31291
rect 21542 31288 21548 31300
rect 21600 31288 21606 31340
rect 23290 31288 23296 31340
rect 23348 31328 23354 31340
rect 25240 31337 25268 31368
rect 27908 31368 28856 31396
rect 23385 31331 23443 31337
rect 23385 31328 23397 31331
rect 23348 31300 23397 31328
rect 23348 31288 23354 31300
rect 23385 31297 23397 31300
rect 23431 31297 23443 31331
rect 23385 31291 23443 31297
rect 23652 31331 23710 31337
rect 23652 31297 23664 31331
rect 23698 31328 23710 31331
rect 24857 31331 24915 31337
rect 24857 31328 24869 31331
rect 23698 31300 24869 31328
rect 23698 31297 23710 31300
rect 23652 31291 23710 31297
rect 24857 31297 24869 31300
rect 24903 31297 24915 31331
rect 24857 31291 24915 31297
rect 25041 31331 25099 31337
rect 25041 31297 25053 31331
rect 25087 31297 25099 31331
rect 25041 31291 25099 31297
rect 25225 31331 25283 31337
rect 25225 31297 25237 31331
rect 25271 31297 25283 31331
rect 25409 31331 25467 31337
rect 25409 31328 25421 31331
rect 25225 31291 25283 31297
rect 25332 31300 25421 31328
rect 20088 31232 20668 31260
rect 18417 31195 18475 31201
rect 18417 31161 18429 31195
rect 18463 31161 18475 31195
rect 18417 31155 18475 31161
rect 19536 31136 19564 31232
rect 20714 31220 20720 31272
rect 20772 31260 20778 31272
rect 21266 31260 21272 31272
rect 20772 31232 21272 31260
rect 20772 31220 20778 31232
rect 21266 31220 21272 31232
rect 21324 31260 21330 31272
rect 21818 31260 21824 31272
rect 21324 31232 21824 31260
rect 21324 31220 21330 31232
rect 21818 31220 21824 31232
rect 21876 31220 21882 31272
rect 25056 31260 25084 31291
rect 25332 31269 25360 31300
rect 25409 31297 25421 31300
rect 25455 31297 25467 31331
rect 25409 31291 25467 31297
rect 27430 31288 27436 31340
rect 27488 31328 27494 31340
rect 27908 31337 27936 31368
rect 28828 31340 28856 31368
rect 27893 31331 27951 31337
rect 27893 31328 27905 31331
rect 27488 31300 27905 31328
rect 27488 31288 27494 31300
rect 27893 31297 27905 31300
rect 27939 31297 27951 31331
rect 28077 31331 28135 31337
rect 28077 31328 28089 31331
rect 27893 31291 27951 31297
rect 28000 31300 28089 31328
rect 24688 31232 25084 31260
rect 25317 31263 25375 31269
rect 19705 31195 19763 31201
rect 19705 31161 19717 31195
rect 19751 31192 19763 31195
rect 20346 31192 20352 31204
rect 19751 31164 20352 31192
rect 19751 31161 19763 31164
rect 19705 31155 19763 31161
rect 20346 31152 20352 31164
rect 20404 31152 20410 31204
rect 24688 31136 24716 31232
rect 25317 31229 25329 31263
rect 25363 31229 25375 31263
rect 25317 31223 25375 31229
rect 25332 31192 25360 31223
rect 24780 31164 25360 31192
rect 24780 31136 24808 31164
rect 28000 31136 28028 31300
rect 28077 31297 28089 31300
rect 28123 31297 28135 31331
rect 28077 31291 28135 31297
rect 28810 31288 28816 31340
rect 28868 31288 28874 31340
rect 29917 31331 29975 31337
rect 29917 31297 29929 31331
rect 29963 31328 29975 31331
rect 30300 31328 30328 31424
rect 30668 31337 30696 31436
rect 31297 31433 31309 31436
rect 31343 31464 31355 31467
rect 32125 31467 32183 31473
rect 32125 31464 32137 31467
rect 31343 31436 32137 31464
rect 31343 31433 31355 31436
rect 31297 31427 31355 31433
rect 32125 31433 32137 31436
rect 32171 31433 32183 31467
rect 32125 31427 32183 31433
rect 31110 31356 31116 31408
rect 31168 31396 31174 31408
rect 31168 31368 31616 31396
rect 31168 31356 31174 31368
rect 29963 31300 30328 31328
rect 30377 31331 30435 31337
rect 29963 31297 29975 31300
rect 29917 31291 29975 31297
rect 30377 31297 30389 31331
rect 30423 31297 30435 31331
rect 30377 31291 30435 31297
rect 30653 31331 30711 31337
rect 30653 31297 30665 31331
rect 30699 31297 30711 31331
rect 30653 31291 30711 31297
rect 30392 31260 30420 31291
rect 30742 31288 30748 31340
rect 30800 31288 30806 31340
rect 30837 31331 30895 31337
rect 30837 31297 30849 31331
rect 30883 31328 30895 31331
rect 31205 31331 31263 31337
rect 31205 31328 31217 31331
rect 30883 31300 31217 31328
rect 30883 31297 30895 31300
rect 30837 31291 30895 31297
rect 31205 31297 31217 31300
rect 31251 31328 31263 31331
rect 31386 31328 31392 31340
rect 31251 31300 31392 31328
rect 31251 31297 31263 31300
rect 31205 31291 31263 31297
rect 31386 31288 31392 31300
rect 31444 31288 31450 31340
rect 31588 31337 31616 31368
rect 31662 31356 31668 31408
rect 31720 31356 31726 31408
rect 31956 31368 33548 31396
rect 31573 31331 31631 31337
rect 31573 31297 31585 31331
rect 31619 31297 31631 31331
rect 31573 31291 31631 31297
rect 30760 31260 30788 31288
rect 31113 31263 31171 31269
rect 31113 31260 31125 31263
rect 30392 31232 31125 31260
rect 31113 31229 31125 31232
rect 31159 31229 31171 31263
rect 31113 31223 31171 31229
rect 31481 31263 31539 31269
rect 31481 31229 31493 31263
rect 31527 31260 31539 31263
rect 31680 31260 31708 31356
rect 31956 31340 31984 31368
rect 31849 31331 31907 31337
rect 31849 31297 31861 31331
rect 31895 31328 31907 31331
rect 31938 31328 31944 31340
rect 31895 31300 31944 31328
rect 31895 31297 31907 31300
rect 31849 31291 31907 31297
rect 31938 31288 31944 31300
rect 31996 31288 32002 31340
rect 32674 31288 32680 31340
rect 32732 31328 32738 31340
rect 33520 31337 33548 31368
rect 33238 31331 33296 31337
rect 33238 31328 33250 31331
rect 32732 31300 33250 31328
rect 32732 31288 32738 31300
rect 33238 31297 33250 31300
rect 33284 31297 33296 31331
rect 33238 31291 33296 31297
rect 33505 31331 33563 31337
rect 33505 31297 33517 31331
rect 33551 31297 33563 31331
rect 33505 31291 33563 31297
rect 31527 31232 31708 31260
rect 31527 31229 31539 31232
rect 31481 31223 31539 31229
rect 30374 31152 30380 31204
rect 30432 31192 30438 31204
rect 30469 31195 30527 31201
rect 30469 31192 30481 31195
rect 30432 31164 30481 31192
rect 30432 31152 30438 31164
rect 30469 31161 30481 31164
rect 30515 31161 30527 31195
rect 30469 31155 30527 31161
rect 30561 31195 30619 31201
rect 30561 31161 30573 31195
rect 30607 31192 30619 31195
rect 31496 31192 31524 31223
rect 30607 31164 31524 31192
rect 30607 31161 30619 31164
rect 30561 31155 30619 31161
rect 17954 31084 17960 31136
rect 18012 31124 18018 31136
rect 18049 31127 18107 31133
rect 18049 31124 18061 31127
rect 18012 31096 18061 31124
rect 18012 31084 18018 31096
rect 18049 31093 18061 31096
rect 18095 31124 18107 31127
rect 19150 31124 19156 31136
rect 18095 31096 19156 31124
rect 18095 31093 18107 31096
rect 18049 31087 18107 31093
rect 19150 31084 19156 31096
rect 19208 31084 19214 31136
rect 19518 31084 19524 31136
rect 19576 31084 19582 31136
rect 19978 31084 19984 31136
rect 20036 31084 20042 31136
rect 20438 31084 20444 31136
rect 20496 31124 20502 31136
rect 21453 31127 21511 31133
rect 21453 31124 21465 31127
rect 20496 31096 21465 31124
rect 20496 31084 20502 31096
rect 21453 31093 21465 31096
rect 21499 31093 21511 31127
rect 21453 31087 21511 31093
rect 24670 31084 24676 31136
rect 24728 31084 24734 31136
rect 24762 31084 24768 31136
rect 24820 31084 24826 31136
rect 25498 31084 25504 31136
rect 25556 31084 25562 31136
rect 27982 31084 27988 31136
rect 28040 31084 28046 31136
rect 28074 31084 28080 31136
rect 28132 31084 28138 31136
rect 29733 31127 29791 31133
rect 29733 31093 29745 31127
rect 29779 31124 29791 31127
rect 29822 31124 29828 31136
rect 29779 31096 29828 31124
rect 29779 31093 29791 31096
rect 29733 31087 29791 31093
rect 29822 31084 29828 31096
rect 29880 31084 29886 31136
rect 30098 31084 30104 31136
rect 30156 31084 30162 31136
rect 30926 31084 30932 31136
rect 30984 31084 30990 31136
rect 31018 31084 31024 31136
rect 31076 31124 31082 31136
rect 31294 31124 31300 31136
rect 31076 31096 31300 31124
rect 31076 31084 31082 31096
rect 31294 31084 31300 31096
rect 31352 31124 31358 31136
rect 31757 31127 31815 31133
rect 31757 31124 31769 31127
rect 31352 31096 31769 31124
rect 31352 31084 31358 31096
rect 31757 31093 31769 31096
rect 31803 31093 31815 31127
rect 31757 31087 31815 31093
rect 1104 31034 34868 31056
rect 1104 30982 5170 31034
rect 5222 30982 5234 31034
rect 5286 30982 5298 31034
rect 5350 30982 5362 31034
rect 5414 30982 5426 31034
rect 5478 30982 13611 31034
rect 13663 30982 13675 31034
rect 13727 30982 13739 31034
rect 13791 30982 13803 31034
rect 13855 30982 13867 31034
rect 13919 30982 22052 31034
rect 22104 30982 22116 31034
rect 22168 30982 22180 31034
rect 22232 30982 22244 31034
rect 22296 30982 22308 31034
rect 22360 30982 30493 31034
rect 30545 30982 30557 31034
rect 30609 30982 30621 31034
rect 30673 30982 30685 31034
rect 30737 30982 30749 31034
rect 30801 30982 34868 31034
rect 1104 30960 34868 30982
rect 16758 30880 16764 30932
rect 16816 30880 16822 30932
rect 17586 30880 17592 30932
rect 17644 30880 17650 30932
rect 17678 30880 17684 30932
rect 17736 30920 17742 30932
rect 17773 30923 17831 30929
rect 17773 30920 17785 30923
rect 17736 30892 17785 30920
rect 17736 30880 17742 30892
rect 17773 30889 17785 30892
rect 17819 30920 17831 30923
rect 18414 30920 18420 30932
rect 17819 30892 18000 30920
rect 17819 30889 17831 30892
rect 17773 30883 17831 30889
rect 17865 30855 17923 30861
rect 17865 30821 17877 30855
rect 17911 30821 17923 30855
rect 17865 30815 17923 30821
rect 17880 30784 17908 30815
rect 16960 30756 17908 30784
rect 16960 30725 16988 30756
rect 16945 30719 17003 30725
rect 16945 30685 16957 30719
rect 16991 30685 17003 30719
rect 16945 30679 17003 30685
rect 17126 30676 17132 30728
rect 17184 30676 17190 30728
rect 17221 30719 17279 30725
rect 17221 30685 17233 30719
rect 17267 30716 17279 30719
rect 17865 30719 17923 30725
rect 17267 30688 17448 30716
rect 17267 30685 17279 30688
rect 17221 30679 17279 30685
rect 17420 30657 17448 30688
rect 17865 30685 17877 30719
rect 17911 30716 17923 30719
rect 17972 30716 18000 30892
rect 18064 30892 18420 30920
rect 18064 30725 18092 30892
rect 18414 30880 18420 30892
rect 18472 30920 18478 30932
rect 23382 30920 23388 30932
rect 18472 30892 20300 30920
rect 18472 30880 18478 30892
rect 18506 30852 18512 30864
rect 18248 30824 18512 30852
rect 18248 30793 18276 30824
rect 18506 30812 18512 30824
rect 18564 30812 18570 30864
rect 18874 30812 18880 30864
rect 18932 30852 18938 30864
rect 18932 30824 19656 30852
rect 18932 30812 18938 30824
rect 18233 30787 18291 30793
rect 18233 30753 18245 30787
rect 18279 30753 18291 30787
rect 18233 30747 18291 30753
rect 19058 30744 19064 30796
rect 19116 30784 19122 30796
rect 19116 30756 19288 30784
rect 19116 30744 19122 30756
rect 17911 30688 18000 30716
rect 18049 30719 18107 30725
rect 17911 30685 17923 30688
rect 17865 30679 17923 30685
rect 18049 30685 18061 30719
rect 18095 30685 18107 30719
rect 18049 30679 18107 30685
rect 18509 30719 18567 30725
rect 18509 30685 18521 30719
rect 18555 30716 18567 30719
rect 18690 30716 18696 30728
rect 18555 30688 18696 30716
rect 18555 30685 18567 30688
rect 18509 30679 18567 30685
rect 18690 30676 18696 30688
rect 18748 30676 18754 30728
rect 18785 30719 18843 30725
rect 18785 30685 18797 30719
rect 18831 30685 18843 30719
rect 18785 30679 18843 30685
rect 17405 30651 17463 30657
rect 17405 30617 17417 30651
rect 17451 30648 17463 30651
rect 17954 30648 17960 30660
rect 17451 30620 17960 30648
rect 17451 30617 17463 30620
rect 17405 30611 17463 30617
rect 17954 30608 17960 30620
rect 18012 30608 18018 30660
rect 18800 30648 18828 30679
rect 18874 30676 18880 30728
rect 18932 30716 18938 30728
rect 19260 30725 19288 30756
rect 18969 30719 19027 30725
rect 18969 30716 18981 30719
rect 18932 30688 18981 30716
rect 18932 30676 18938 30688
rect 18969 30685 18981 30688
rect 19015 30685 19027 30719
rect 18969 30679 19027 30685
rect 19245 30719 19303 30725
rect 19245 30685 19257 30719
rect 19291 30685 19303 30719
rect 19245 30679 19303 30685
rect 19334 30676 19340 30728
rect 19392 30716 19398 30728
rect 19429 30719 19487 30725
rect 19429 30716 19441 30719
rect 19392 30688 19441 30716
rect 19392 30676 19398 30688
rect 19429 30685 19441 30688
rect 19475 30685 19487 30719
rect 19429 30679 19487 30685
rect 19518 30676 19524 30728
rect 19576 30676 19582 30728
rect 19628 30725 19656 30824
rect 19794 30812 19800 30864
rect 19852 30852 19858 30864
rect 19852 30824 20116 30852
rect 19852 30812 19858 30824
rect 19978 30744 19984 30796
rect 20036 30744 20042 30796
rect 19613 30719 19671 30725
rect 19613 30685 19625 30719
rect 19659 30685 19671 30719
rect 19613 30679 19671 30685
rect 19797 30719 19855 30725
rect 19797 30685 19809 30719
rect 19843 30716 19855 30719
rect 19996 30716 20024 30744
rect 19843 30688 20024 30716
rect 20088 30716 20116 30824
rect 20272 30796 20300 30892
rect 21928 30892 23388 30920
rect 20254 30744 20260 30796
rect 20312 30744 20318 30796
rect 21928 30716 21956 30892
rect 23382 30880 23388 30892
rect 23440 30880 23446 30932
rect 24670 30880 24676 30932
rect 24728 30880 24734 30932
rect 25498 30920 25504 30932
rect 25240 30892 25504 30920
rect 24486 30812 24492 30864
rect 24544 30812 24550 30864
rect 24504 30784 24532 30812
rect 23124 30756 24072 30784
rect 22005 30719 22063 30725
rect 22005 30716 22017 30719
rect 20088 30688 22017 30716
rect 19843 30685 19855 30688
rect 19797 30679 19855 30685
rect 22005 30685 22017 30688
rect 22051 30685 22063 30719
rect 22005 30679 22063 30685
rect 19812 30648 19840 30679
rect 18800 30620 19840 30648
rect 22272 30651 22330 30657
rect 22272 30617 22284 30651
rect 22318 30648 22330 30651
rect 22646 30648 22652 30660
rect 22318 30620 22652 30648
rect 22318 30617 22330 30620
rect 22272 30611 22330 30617
rect 22646 30608 22652 30620
rect 22704 30608 22710 30660
rect 23124 30592 23152 30756
rect 23658 30676 23664 30728
rect 23716 30676 23722 30728
rect 23753 30719 23811 30725
rect 23753 30685 23765 30719
rect 23799 30685 23811 30719
rect 23753 30679 23811 30685
rect 23768 30648 23796 30679
rect 23842 30676 23848 30728
rect 23900 30716 23906 30728
rect 23937 30719 23995 30725
rect 23937 30716 23949 30719
rect 23900 30688 23949 30716
rect 23900 30676 23906 30688
rect 23937 30685 23949 30688
rect 23983 30685 23995 30719
rect 23937 30679 23995 30685
rect 23400 30620 23796 30648
rect 24044 30648 24072 30756
rect 24412 30756 24532 30784
rect 24121 30719 24179 30725
rect 24121 30685 24133 30719
rect 24167 30716 24179 30719
rect 24210 30716 24216 30728
rect 24167 30688 24216 30716
rect 24167 30685 24179 30688
rect 24121 30679 24179 30685
rect 24210 30676 24216 30688
rect 24268 30716 24274 30728
rect 24412 30725 24440 30756
rect 24397 30719 24455 30725
rect 24397 30716 24409 30719
rect 24268 30688 24409 30716
rect 24268 30676 24274 30688
rect 24397 30685 24409 30688
rect 24443 30685 24455 30719
rect 24397 30679 24455 30685
rect 24489 30719 24547 30725
rect 24489 30685 24501 30719
rect 24535 30716 24547 30719
rect 24762 30716 24768 30728
rect 24535 30688 24768 30716
rect 24535 30685 24547 30688
rect 24489 30679 24547 30685
rect 24762 30676 24768 30688
rect 24820 30676 24826 30728
rect 25240 30725 25268 30892
rect 25498 30880 25504 30892
rect 25556 30880 25562 30932
rect 27249 30923 27307 30929
rect 27249 30889 27261 30923
rect 27295 30920 27307 30923
rect 27338 30920 27344 30932
rect 27295 30892 27344 30920
rect 27295 30889 27307 30892
rect 27249 30883 27307 30889
rect 27338 30880 27344 30892
rect 27396 30880 27402 30932
rect 31018 30920 31024 30932
rect 29564 30892 31024 30920
rect 25409 30855 25467 30861
rect 25409 30821 25421 30855
rect 25455 30821 25467 30855
rect 25516 30852 25544 30880
rect 26973 30855 27031 30861
rect 25516 30824 25912 30852
rect 25409 30815 25467 30821
rect 25424 30784 25452 30815
rect 25884 30793 25912 30824
rect 26973 30821 26985 30855
rect 27019 30821 27031 30855
rect 26973 30815 27031 30821
rect 27525 30855 27583 30861
rect 27525 30821 27537 30855
rect 27571 30852 27583 30855
rect 27893 30855 27951 30861
rect 27893 30852 27905 30855
rect 27571 30824 27905 30852
rect 27571 30821 27583 30824
rect 27525 30815 27583 30821
rect 27893 30821 27905 30824
rect 27939 30852 27951 30855
rect 27982 30852 27988 30864
rect 27939 30824 27988 30852
rect 27939 30821 27951 30824
rect 27893 30815 27951 30821
rect 25869 30787 25927 30793
rect 25424 30756 25728 30784
rect 24857 30719 24915 30725
rect 24857 30685 24869 30719
rect 24903 30685 24915 30719
rect 24857 30679 24915 30685
rect 25225 30719 25283 30725
rect 25225 30685 25237 30719
rect 25271 30685 25283 30719
rect 25225 30679 25283 30685
rect 24302 30648 24308 30660
rect 24044 30620 24308 30648
rect 17494 30540 17500 30592
rect 17552 30580 17558 30592
rect 17605 30583 17663 30589
rect 17605 30580 17617 30583
rect 17552 30552 17617 30580
rect 17552 30540 17558 30552
rect 17605 30549 17617 30552
rect 17651 30549 17663 30583
rect 17605 30543 17663 30549
rect 18230 30540 18236 30592
rect 18288 30580 18294 30592
rect 18325 30583 18383 30589
rect 18325 30580 18337 30583
rect 18288 30552 18337 30580
rect 18288 30540 18294 30552
rect 18325 30549 18337 30552
rect 18371 30549 18383 30583
rect 18325 30543 18383 30549
rect 19242 30540 19248 30592
rect 19300 30580 19306 30592
rect 19981 30583 20039 30589
rect 19981 30580 19993 30583
rect 19300 30552 19993 30580
rect 19300 30540 19306 30552
rect 19981 30549 19993 30552
rect 20027 30549 20039 30583
rect 19981 30543 20039 30549
rect 23106 30540 23112 30592
rect 23164 30540 23170 30592
rect 23198 30540 23204 30592
rect 23256 30580 23262 30592
rect 23400 30589 23428 30620
rect 24302 30608 24308 30620
rect 24360 30648 24366 30660
rect 24673 30651 24731 30657
rect 24673 30648 24685 30651
rect 24360 30620 24685 30648
rect 24360 30608 24366 30620
rect 24673 30617 24685 30620
rect 24719 30617 24731 30651
rect 24673 30611 24731 30617
rect 23385 30583 23443 30589
rect 23385 30580 23397 30583
rect 23256 30552 23397 30580
rect 23256 30540 23262 30552
rect 23385 30549 23397 30552
rect 23431 30549 23443 30583
rect 23385 30543 23443 30549
rect 23474 30540 23480 30592
rect 23532 30540 23538 30592
rect 23566 30540 23572 30592
rect 23624 30580 23630 30592
rect 24029 30583 24087 30589
rect 24029 30580 24041 30583
rect 23624 30552 24041 30580
rect 23624 30540 23630 30552
rect 24029 30549 24041 30552
rect 24075 30549 24087 30583
rect 24872 30580 24900 30679
rect 25406 30676 25412 30728
rect 25464 30676 25470 30728
rect 25501 30719 25559 30725
rect 25501 30685 25513 30719
rect 25547 30716 25559 30719
rect 25590 30716 25596 30728
rect 25547 30688 25596 30716
rect 25547 30685 25559 30688
rect 25501 30679 25559 30685
rect 25590 30676 25596 30688
rect 25648 30676 25654 30728
rect 25700 30725 25728 30756
rect 25869 30753 25881 30787
rect 25915 30753 25927 30787
rect 25869 30747 25927 30753
rect 26697 30787 26755 30793
rect 26697 30753 26709 30787
rect 26743 30784 26755 30787
rect 26878 30784 26884 30796
rect 26743 30756 26884 30784
rect 26743 30753 26755 30756
rect 26697 30747 26755 30753
rect 26878 30744 26884 30756
rect 26936 30744 26942 30796
rect 26988 30784 27016 30815
rect 27982 30812 27988 30824
rect 28040 30852 28046 30864
rect 28040 30824 28764 30852
rect 28040 30812 28046 30824
rect 26988 30756 27568 30784
rect 27540 30728 27568 30756
rect 28166 30744 28172 30796
rect 28224 30744 28230 30796
rect 25685 30719 25743 30725
rect 25685 30685 25697 30719
rect 25731 30685 25743 30719
rect 25685 30679 25743 30685
rect 25774 30676 25780 30728
rect 25832 30676 25838 30728
rect 26053 30719 26111 30725
rect 26053 30685 26065 30719
rect 26099 30685 26111 30719
rect 26053 30679 26111 30685
rect 24946 30608 24952 30660
rect 25004 30648 25010 30660
rect 25041 30651 25099 30657
rect 25041 30648 25053 30651
rect 25004 30620 25053 30648
rect 25004 30608 25010 30620
rect 25041 30617 25053 30620
rect 25087 30617 25099 30651
rect 25041 30611 25099 30617
rect 25133 30651 25191 30657
rect 25133 30617 25145 30651
rect 25179 30648 25191 30651
rect 25424 30648 25452 30676
rect 26068 30648 26096 30679
rect 26602 30676 26608 30728
rect 26660 30676 26666 30728
rect 27430 30676 27436 30728
rect 27488 30676 27494 30728
rect 27522 30676 27528 30728
rect 27580 30716 27586 30728
rect 27617 30719 27675 30725
rect 27617 30716 27629 30719
rect 27580 30688 27629 30716
rect 27580 30676 27586 30688
rect 27617 30685 27629 30688
rect 27663 30685 27675 30719
rect 27617 30679 27675 30685
rect 27706 30676 27712 30728
rect 27764 30676 27770 30728
rect 27798 30676 27804 30728
rect 27856 30716 27862 30728
rect 28736 30725 28764 30824
rect 29564 30728 29592 30892
rect 31018 30880 31024 30892
rect 31076 30880 31082 30932
rect 31662 30880 31668 30932
rect 31720 30920 31726 30932
rect 32401 30923 32459 30929
rect 32401 30920 32413 30923
rect 31720 30892 32413 30920
rect 31720 30880 31726 30892
rect 32401 30889 32413 30892
rect 32447 30889 32459 30923
rect 32401 30883 32459 30889
rect 32674 30880 32680 30932
rect 32732 30880 32738 30932
rect 31036 30793 31064 30880
rect 32122 30812 32128 30864
rect 32180 30812 32186 30864
rect 31021 30787 31079 30793
rect 31021 30753 31033 30787
rect 31067 30753 31079 30787
rect 31021 30747 31079 30753
rect 28261 30719 28319 30725
rect 28261 30716 28273 30719
rect 27856 30688 28273 30716
rect 27856 30676 27862 30688
rect 28261 30685 28273 30688
rect 28307 30685 28319 30719
rect 28261 30679 28319 30685
rect 28721 30719 28779 30725
rect 28721 30685 28733 30719
rect 28767 30685 28779 30719
rect 28721 30679 28779 30685
rect 28810 30676 28816 30728
rect 28868 30676 28874 30728
rect 29546 30676 29552 30728
rect 29604 30676 29610 30728
rect 29822 30725 29828 30728
rect 29816 30716 29828 30725
rect 29783 30688 29828 30716
rect 29816 30679 29828 30688
rect 29822 30676 29828 30679
rect 29880 30676 29886 30728
rect 32140 30716 32168 30812
rect 32493 30719 32551 30725
rect 32493 30716 32505 30719
rect 32140 30688 32505 30716
rect 32493 30685 32505 30688
rect 32539 30685 32551 30719
rect 32493 30679 32551 30685
rect 31288 30651 31346 30657
rect 25179 30620 26096 30648
rect 26252 30620 31064 30648
rect 25179 30617 25191 30620
rect 25133 30611 25191 30617
rect 25682 30580 25688 30592
rect 24872 30552 25688 30580
rect 24029 30543 24087 30549
rect 25682 30540 25688 30552
rect 25740 30540 25746 30592
rect 26252 30589 26280 30620
rect 26237 30583 26295 30589
rect 26237 30549 26249 30583
rect 26283 30549 26295 30583
rect 26237 30543 26295 30549
rect 26878 30540 26884 30592
rect 26936 30580 26942 30592
rect 27890 30580 27896 30592
rect 26936 30552 27896 30580
rect 26936 30540 26942 30552
rect 27890 30540 27896 30552
rect 27948 30580 27954 30592
rect 28166 30580 28172 30592
rect 27948 30552 28172 30580
rect 27948 30540 27954 30552
rect 28166 30540 28172 30552
rect 28224 30540 28230 30592
rect 28534 30540 28540 30592
rect 28592 30540 28598 30592
rect 30006 30540 30012 30592
rect 30064 30580 30070 30592
rect 30650 30580 30656 30592
rect 30064 30552 30656 30580
rect 30064 30540 30070 30552
rect 30650 30540 30656 30552
rect 30708 30580 30714 30592
rect 30929 30583 30987 30589
rect 30929 30580 30941 30583
rect 30708 30552 30941 30580
rect 30708 30540 30714 30552
rect 30929 30549 30941 30552
rect 30975 30549 30987 30583
rect 31036 30580 31064 30620
rect 31288 30617 31300 30651
rect 31334 30648 31346 30651
rect 31386 30648 31392 30660
rect 31334 30620 31392 30648
rect 31334 30617 31346 30620
rect 31288 30611 31346 30617
rect 31386 30608 31392 30620
rect 31444 30608 31450 30660
rect 34146 30580 34152 30592
rect 31036 30552 34152 30580
rect 30929 30543 30987 30549
rect 34146 30540 34152 30552
rect 34204 30540 34210 30592
rect 1104 30490 35027 30512
rect 1104 30438 9390 30490
rect 9442 30438 9454 30490
rect 9506 30438 9518 30490
rect 9570 30438 9582 30490
rect 9634 30438 9646 30490
rect 9698 30438 17831 30490
rect 17883 30438 17895 30490
rect 17947 30438 17959 30490
rect 18011 30438 18023 30490
rect 18075 30438 18087 30490
rect 18139 30438 26272 30490
rect 26324 30438 26336 30490
rect 26388 30438 26400 30490
rect 26452 30438 26464 30490
rect 26516 30438 26528 30490
rect 26580 30438 34713 30490
rect 34765 30438 34777 30490
rect 34829 30438 34841 30490
rect 34893 30438 34905 30490
rect 34957 30438 34969 30490
rect 35021 30438 35027 30490
rect 1104 30416 35027 30438
rect 17586 30336 17592 30388
rect 17644 30376 17650 30388
rect 18049 30379 18107 30385
rect 18049 30376 18061 30379
rect 17644 30348 18061 30376
rect 17644 30336 17650 30348
rect 18049 30345 18061 30348
rect 18095 30376 18107 30379
rect 18969 30379 19027 30385
rect 18095 30348 18460 30376
rect 18095 30345 18107 30348
rect 18049 30339 18107 30345
rect 1765 30311 1823 30317
rect 1765 30277 1777 30311
rect 1811 30308 1823 30311
rect 18230 30308 18236 30320
rect 1811 30280 18236 30308
rect 1811 30277 1823 30280
rect 1765 30271 1823 30277
rect 18230 30268 18236 30280
rect 18288 30268 18294 30320
rect 18432 30308 18460 30348
rect 18969 30345 18981 30379
rect 19015 30376 19027 30379
rect 19058 30376 19064 30388
rect 19015 30348 19064 30376
rect 19015 30345 19027 30348
rect 18969 30339 19027 30345
rect 19058 30336 19064 30348
rect 19116 30336 19122 30388
rect 20254 30336 20260 30388
rect 20312 30376 20318 30388
rect 23106 30376 23112 30388
rect 20312 30348 23112 30376
rect 20312 30336 20318 30348
rect 23106 30336 23112 30348
rect 23164 30336 23170 30388
rect 23382 30336 23388 30388
rect 23440 30336 23446 30388
rect 25774 30336 25780 30388
rect 25832 30376 25838 30388
rect 25869 30379 25927 30385
rect 25869 30376 25881 30379
rect 25832 30348 25881 30376
rect 25832 30336 25838 30348
rect 25869 30345 25881 30348
rect 25915 30345 25927 30379
rect 26602 30376 26608 30388
rect 25869 30339 25927 30345
rect 26068 30348 26608 30376
rect 18601 30311 18659 30317
rect 18601 30308 18613 30311
rect 18432 30280 18613 30308
rect 18601 30277 18613 30280
rect 18647 30277 18659 30311
rect 18601 30271 18659 30277
rect 18693 30311 18751 30317
rect 18693 30277 18705 30311
rect 18739 30308 18751 30311
rect 19518 30308 19524 30320
rect 18739 30280 19524 30308
rect 18739 30277 18751 30280
rect 18693 30271 18751 30277
rect 19518 30268 19524 30280
rect 19576 30268 19582 30320
rect 23400 30308 23428 30336
rect 20180 30280 21312 30308
rect 16301 30243 16359 30249
rect 16301 30209 16313 30243
rect 16347 30240 16359 30243
rect 16485 30243 16543 30249
rect 16347 30212 16436 30240
rect 16347 30209 16359 30212
rect 16301 30203 16359 30209
rect 16408 30048 16436 30212
rect 16485 30209 16497 30243
rect 16531 30240 16543 30243
rect 16531 30212 16620 30240
rect 16531 30209 16543 30212
rect 16485 30203 16543 30209
rect 934 29996 940 30048
rect 992 30036 998 30048
rect 1489 30039 1547 30045
rect 1489 30036 1501 30039
rect 992 30008 1501 30036
rect 992 29996 998 30008
rect 1489 30005 1501 30008
rect 1535 30005 1547 30039
rect 1489 29999 1547 30005
rect 16390 29996 16396 30048
rect 16448 29996 16454 30048
rect 16482 29996 16488 30048
rect 16540 29996 16546 30048
rect 16592 30036 16620 30212
rect 16758 30200 16764 30252
rect 16816 30240 16822 30252
rect 16925 30243 16983 30249
rect 16925 30240 16937 30243
rect 16816 30212 16937 30240
rect 16816 30200 16822 30212
rect 16925 30209 16937 30212
rect 16971 30209 16983 30243
rect 16925 30203 16983 30209
rect 18322 30200 18328 30252
rect 18380 30200 18386 30252
rect 18445 30243 18503 30249
rect 18445 30209 18457 30243
rect 18491 30240 18503 30243
rect 18831 30243 18889 30249
rect 18491 30212 18727 30240
rect 18491 30209 18503 30212
rect 18445 30203 18503 30209
rect 16666 30132 16672 30184
rect 16724 30132 16730 30184
rect 18699 30172 18727 30212
rect 18831 30209 18843 30243
rect 18877 30240 18889 30243
rect 19150 30240 19156 30252
rect 18877 30212 19156 30240
rect 18877 30209 18889 30212
rect 18831 30203 18889 30209
rect 19150 30200 19156 30212
rect 19208 30200 19214 30252
rect 19242 30200 19248 30252
rect 19300 30240 19306 30252
rect 20180 30240 20208 30280
rect 19300 30212 20208 30240
rect 19300 30200 19306 30212
rect 20254 30200 20260 30252
rect 20312 30200 20318 30252
rect 20438 30200 20444 30252
rect 20496 30200 20502 30252
rect 20717 30243 20775 30249
rect 20717 30209 20729 30243
rect 20763 30240 20775 30243
rect 20806 30240 20812 30252
rect 20763 30212 20812 30240
rect 20763 30209 20775 30212
rect 20717 30203 20775 30209
rect 20806 30200 20812 30212
rect 20864 30200 20870 30252
rect 20898 30200 20904 30252
rect 20956 30200 20962 30252
rect 21085 30243 21143 30249
rect 21085 30209 21097 30243
rect 21131 30240 21143 30243
rect 21174 30240 21180 30252
rect 21131 30212 21180 30240
rect 21131 30209 21143 30212
rect 21085 30203 21143 30209
rect 21174 30200 21180 30212
rect 21232 30200 21238 30252
rect 21284 30249 21312 30280
rect 23308 30280 23428 30308
rect 24857 30311 24915 30317
rect 23308 30249 23336 30280
rect 24857 30277 24869 30311
rect 24903 30308 24915 30311
rect 26068 30308 26096 30348
rect 26602 30336 26608 30348
rect 26660 30336 26666 30388
rect 27522 30336 27528 30388
rect 27580 30376 27586 30388
rect 27580 30348 28856 30376
rect 27580 30336 27586 30348
rect 28721 30311 28779 30317
rect 28721 30308 28733 30311
rect 24903 30280 25360 30308
rect 24903 30277 24915 30280
rect 24857 30271 24915 30277
rect 25332 30252 25360 30280
rect 25424 30280 26096 30308
rect 26160 30280 28733 30308
rect 21269 30243 21327 30249
rect 21269 30209 21281 30243
rect 21315 30209 21327 30243
rect 21269 30203 21327 30209
rect 21453 30243 21511 30249
rect 21453 30209 21465 30243
rect 21499 30240 21511 30243
rect 22934 30243 22992 30249
rect 22934 30240 22946 30243
rect 21499 30212 22946 30240
rect 21499 30209 21511 30212
rect 21453 30203 21511 30209
rect 22934 30209 22946 30212
rect 22980 30209 22992 30243
rect 22934 30203 22992 30209
rect 23201 30243 23259 30249
rect 23201 30209 23213 30243
rect 23247 30240 23259 30243
rect 23293 30243 23351 30249
rect 23293 30240 23305 30243
rect 23247 30212 23305 30240
rect 23247 30209 23259 30212
rect 23201 30203 23259 30209
rect 23293 30209 23305 30212
rect 23339 30209 23351 30243
rect 23293 30203 23351 30209
rect 20272 30172 20300 30200
rect 20530 30172 20536 30184
rect 18699 30144 19196 30172
rect 20272 30144 20536 30172
rect 19168 30048 19196 30144
rect 20530 30132 20536 30144
rect 20588 30132 20594 30184
rect 20990 30132 20996 30184
rect 21048 30132 21054 30184
rect 20346 30064 20352 30116
rect 20404 30104 20410 30116
rect 20622 30104 20628 30116
rect 20404 30076 20628 30104
rect 20404 30064 20410 30076
rect 20622 30064 20628 30076
rect 20680 30064 20686 30116
rect 21284 30104 21312 30203
rect 23382 30200 23388 30252
rect 23440 30240 23446 30252
rect 23549 30243 23607 30249
rect 23549 30240 23561 30243
rect 23440 30212 23561 30240
rect 23440 30200 23446 30212
rect 23549 30209 23561 30212
rect 23595 30209 23607 30243
rect 23549 30203 23607 30209
rect 24026 30200 24032 30252
rect 24084 30240 24090 30252
rect 24765 30243 24823 30249
rect 24765 30240 24777 30243
rect 24084 30212 24777 30240
rect 24084 30200 24090 30212
rect 24765 30209 24777 30212
rect 24811 30209 24823 30243
rect 24765 30203 24823 30209
rect 25130 30200 25136 30252
rect 25188 30200 25194 30252
rect 25314 30200 25320 30252
rect 25372 30200 25378 30252
rect 25424 30249 25452 30280
rect 25409 30243 25467 30249
rect 25409 30209 25421 30243
rect 25455 30209 25467 30243
rect 25409 30203 25467 30209
rect 25590 30200 25596 30252
rect 25648 30200 25654 30252
rect 25682 30200 25688 30252
rect 25740 30200 25746 30252
rect 26160 30249 26188 30280
rect 28721 30277 28733 30280
rect 28767 30277 28779 30311
rect 28721 30271 28779 30277
rect 25961 30243 26019 30249
rect 25961 30209 25973 30243
rect 26007 30209 26019 30243
rect 25961 30203 26019 30209
rect 26145 30243 26203 30249
rect 26145 30209 26157 30243
rect 26191 30209 26203 30243
rect 26145 30203 26203 30209
rect 24946 30132 24952 30184
rect 25004 30132 25010 30184
rect 25501 30175 25559 30181
rect 25501 30141 25513 30175
rect 25547 30141 25559 30175
rect 25608 30172 25636 30200
rect 25976 30172 26004 30203
rect 26326 30200 26332 30252
rect 26384 30200 26390 30252
rect 26513 30243 26571 30249
rect 26513 30209 26525 30243
rect 26559 30240 26571 30243
rect 26602 30240 26608 30252
rect 26559 30212 26608 30240
rect 26559 30209 26571 30212
rect 26513 30203 26571 30209
rect 26602 30200 26608 30212
rect 26660 30240 26666 30252
rect 27249 30243 27307 30249
rect 26660 30212 27108 30240
rect 26660 30200 26666 30212
rect 25608 30144 26004 30172
rect 26237 30175 26295 30181
rect 25501 30135 25559 30141
rect 26237 30141 26249 30175
rect 26283 30141 26295 30175
rect 26344 30172 26372 30200
rect 26878 30172 26884 30184
rect 26344 30144 26884 30172
rect 26237 30135 26295 30141
rect 21542 30104 21548 30116
rect 21284 30076 21548 30104
rect 21542 30064 21548 30076
rect 21600 30104 21606 30116
rect 21821 30107 21879 30113
rect 21821 30104 21833 30107
rect 21600 30076 21833 30104
rect 21600 30064 21606 30076
rect 21821 30073 21833 30076
rect 21867 30073 21879 30107
rect 24964 30104 24992 30132
rect 25516 30104 25544 30135
rect 24964 30076 25544 30104
rect 26252 30104 26280 30135
rect 26878 30132 26884 30144
rect 26936 30132 26942 30184
rect 26973 30107 27031 30113
rect 26973 30104 26985 30107
rect 26252 30076 26985 30104
rect 21821 30067 21879 30073
rect 26973 30073 26985 30076
rect 27019 30073 27031 30107
rect 26973 30067 27031 30073
rect 17034 30036 17040 30048
rect 16592 30008 17040 30036
rect 17034 29996 17040 30008
rect 17092 29996 17098 30048
rect 19150 29996 19156 30048
rect 19208 29996 19214 30048
rect 20070 29996 20076 30048
rect 20128 30036 20134 30048
rect 21266 30036 21272 30048
rect 20128 30008 21272 30036
rect 20128 29996 20134 30008
rect 21266 29996 21272 30008
rect 21324 29996 21330 30048
rect 24670 29996 24676 30048
rect 24728 29996 24734 30048
rect 26694 29996 26700 30048
rect 26752 29996 26758 30048
rect 27080 30036 27108 30212
rect 27249 30209 27261 30243
rect 27295 30240 27307 30243
rect 27522 30240 27528 30252
rect 27295 30212 27528 30240
rect 27295 30209 27307 30212
rect 27249 30203 27307 30209
rect 27522 30200 27528 30212
rect 27580 30200 27586 30252
rect 27614 30200 27620 30252
rect 27672 30200 27678 30252
rect 27709 30243 27767 30249
rect 27709 30209 27721 30243
rect 27755 30209 27767 30243
rect 27709 30203 27767 30209
rect 27157 30175 27215 30181
rect 27157 30141 27169 30175
rect 27203 30141 27215 30175
rect 27724 30172 27752 30203
rect 27798 30200 27804 30252
rect 27856 30200 27862 30252
rect 27890 30200 27896 30252
rect 27948 30200 27954 30252
rect 27985 30243 28043 30249
rect 27985 30209 27997 30243
rect 28031 30240 28043 30243
rect 28074 30240 28080 30252
rect 28031 30212 28080 30240
rect 28031 30209 28043 30212
rect 27985 30203 28043 30209
rect 28074 30200 28080 30212
rect 28132 30240 28138 30252
rect 28132 30212 28396 30240
rect 28132 30200 28138 30212
rect 27908 30172 27936 30200
rect 27724 30144 27936 30172
rect 27157 30135 27215 30141
rect 27172 30104 27200 30135
rect 28258 30132 28264 30184
rect 28316 30132 28322 30184
rect 28368 30172 28396 30212
rect 28534 30200 28540 30252
rect 28592 30200 28598 30252
rect 28828 30249 28856 30348
rect 30098 30336 30104 30388
rect 30156 30336 30162 30388
rect 30926 30336 30932 30388
rect 30984 30336 30990 30388
rect 31386 30336 31392 30388
rect 31444 30336 31450 30388
rect 30116 30308 30144 30336
rect 30944 30308 30972 30336
rect 30116 30280 30236 30308
rect 28629 30243 28687 30249
rect 28629 30209 28641 30243
rect 28675 30209 28687 30243
rect 28629 30203 28687 30209
rect 28813 30243 28871 30249
rect 28813 30209 28825 30243
rect 28859 30209 28871 30243
rect 28813 30203 28871 30209
rect 28445 30175 28503 30181
rect 28445 30172 28457 30175
rect 28368 30144 28457 30172
rect 28445 30141 28457 30144
rect 28491 30141 28503 30175
rect 28445 30135 28503 30141
rect 28644 30116 28672 30203
rect 30006 30200 30012 30252
rect 30064 30240 30070 30252
rect 30208 30249 30236 30280
rect 30300 30280 30972 30308
rect 30300 30249 30328 30280
rect 30101 30243 30159 30249
rect 30101 30240 30113 30243
rect 30064 30212 30113 30240
rect 30064 30200 30070 30212
rect 30101 30209 30113 30212
rect 30147 30209 30159 30243
rect 30101 30203 30159 30209
rect 30193 30243 30251 30249
rect 30193 30209 30205 30243
rect 30239 30209 30251 30243
rect 30193 30203 30251 30209
rect 30285 30243 30343 30249
rect 30285 30209 30297 30243
rect 30331 30209 30343 30243
rect 30469 30243 30527 30249
rect 30469 30240 30481 30243
rect 30285 30203 30343 30209
rect 30392 30212 30481 30240
rect 27982 30104 27988 30116
rect 27172 30076 27988 30104
rect 27982 30064 27988 30076
rect 28040 30064 28046 30116
rect 28353 30107 28411 30113
rect 28353 30073 28365 30107
rect 28399 30104 28411 30107
rect 28534 30104 28540 30116
rect 28399 30076 28540 30104
rect 28399 30073 28411 30076
rect 28353 30067 28411 30073
rect 28534 30064 28540 30076
rect 28592 30064 28598 30116
rect 28626 30064 28632 30116
rect 28684 30064 28690 30116
rect 30392 30104 30420 30212
rect 30469 30209 30481 30212
rect 30515 30209 30527 30243
rect 30469 30203 30527 30209
rect 30650 30200 30656 30252
rect 30708 30200 30714 30252
rect 30745 30243 30803 30249
rect 30745 30209 30757 30243
rect 30791 30209 30803 30243
rect 30745 30203 30803 30209
rect 30929 30243 30987 30249
rect 30929 30209 30941 30243
rect 30975 30240 30987 30243
rect 31205 30243 31263 30249
rect 31205 30240 31217 30243
rect 30975 30212 31217 30240
rect 30975 30209 30987 30212
rect 30929 30203 30987 30209
rect 31205 30209 31217 30212
rect 31251 30209 31263 30243
rect 31205 30203 31263 30209
rect 30760 30172 30788 30203
rect 31846 30200 31852 30252
rect 31904 30200 31910 30252
rect 30760 30144 31248 30172
rect 31220 30116 31248 30144
rect 28966 30076 30420 30104
rect 27430 30036 27436 30048
rect 27080 30008 27436 30036
rect 27430 29996 27436 30008
rect 27488 29996 27494 30048
rect 28166 29996 28172 30048
rect 28224 29996 28230 30048
rect 28442 29996 28448 30048
rect 28500 30036 28506 30048
rect 28966 30036 28994 30076
rect 31202 30064 31208 30116
rect 31260 30064 31266 30116
rect 28500 30008 28994 30036
rect 28500 29996 28506 30008
rect 29822 29996 29828 30048
rect 29880 29996 29886 30048
rect 31570 29996 31576 30048
rect 31628 30036 31634 30048
rect 31665 30039 31723 30045
rect 31665 30036 31677 30039
rect 31628 30008 31677 30036
rect 31628 29996 31634 30008
rect 31665 30005 31677 30008
rect 31711 30005 31723 30039
rect 31665 29999 31723 30005
rect 1104 29946 34868 29968
rect 1104 29894 5170 29946
rect 5222 29894 5234 29946
rect 5286 29894 5298 29946
rect 5350 29894 5362 29946
rect 5414 29894 5426 29946
rect 5478 29894 13611 29946
rect 13663 29894 13675 29946
rect 13727 29894 13739 29946
rect 13791 29894 13803 29946
rect 13855 29894 13867 29946
rect 13919 29894 22052 29946
rect 22104 29894 22116 29946
rect 22168 29894 22180 29946
rect 22232 29894 22244 29946
rect 22296 29894 22308 29946
rect 22360 29894 30493 29946
rect 30545 29894 30557 29946
rect 30609 29894 30621 29946
rect 30673 29894 30685 29946
rect 30737 29894 30749 29946
rect 30801 29894 34868 29946
rect 1104 29872 34868 29894
rect 16482 29792 16488 29844
rect 16540 29792 16546 29844
rect 16669 29835 16727 29841
rect 16669 29801 16681 29835
rect 16715 29832 16727 29835
rect 16758 29832 16764 29844
rect 16715 29804 16764 29832
rect 16715 29801 16727 29804
rect 16669 29795 16727 29801
rect 16758 29792 16764 29804
rect 16816 29792 16822 29844
rect 17126 29792 17132 29844
rect 17184 29832 17190 29844
rect 17221 29835 17279 29841
rect 17221 29832 17233 29835
rect 17184 29804 17233 29832
rect 17184 29792 17190 29804
rect 17221 29801 17233 29804
rect 17267 29801 17279 29835
rect 17221 29795 17279 29801
rect 18141 29835 18199 29841
rect 18141 29801 18153 29835
rect 18187 29832 18199 29835
rect 18322 29832 18328 29844
rect 18187 29804 18328 29832
rect 18187 29801 18199 29804
rect 18141 29795 18199 29801
rect 18322 29792 18328 29804
rect 18380 29792 18386 29844
rect 19150 29792 19156 29844
rect 19208 29792 19214 29844
rect 19242 29792 19248 29844
rect 19300 29792 19306 29844
rect 20456 29804 20852 29832
rect 16500 29628 16528 29792
rect 17129 29699 17187 29705
rect 17129 29665 17141 29699
rect 17175 29696 17187 29699
rect 17586 29696 17592 29708
rect 17175 29668 17592 29696
rect 17175 29665 17187 29668
rect 17129 29659 17187 29665
rect 17586 29656 17592 29668
rect 17644 29656 17650 29708
rect 19168 29696 19196 29792
rect 18340 29668 19196 29696
rect 16853 29631 16911 29637
rect 16853 29628 16865 29631
rect 16500 29600 16865 29628
rect 16853 29597 16865 29600
rect 16899 29597 16911 29631
rect 16853 29591 16911 29597
rect 17037 29631 17095 29637
rect 17037 29597 17049 29631
rect 17083 29597 17095 29631
rect 17037 29591 17095 29597
rect 17405 29631 17463 29637
rect 17405 29597 17417 29631
rect 17451 29597 17463 29631
rect 17405 29591 17463 29597
rect 17052 29560 17080 29591
rect 17420 29560 17448 29591
rect 17052 29532 17448 29560
rect 17604 29560 17632 29656
rect 18340 29637 18368 29668
rect 18325 29631 18383 29637
rect 18325 29597 18337 29631
rect 18371 29597 18383 29631
rect 18325 29591 18383 29597
rect 18509 29631 18567 29637
rect 18509 29597 18521 29631
rect 18555 29597 18567 29631
rect 18509 29591 18567 29597
rect 18524 29560 18552 29591
rect 18598 29588 18604 29640
rect 18656 29588 18662 29640
rect 18690 29588 18696 29640
rect 18748 29588 18754 29640
rect 18874 29588 18880 29640
rect 18932 29588 18938 29640
rect 19260 29628 19288 29792
rect 19797 29767 19855 29773
rect 19797 29733 19809 29767
rect 19843 29764 19855 29767
rect 19886 29764 19892 29776
rect 19843 29736 19892 29764
rect 19843 29733 19855 29736
rect 19797 29727 19855 29733
rect 19886 29724 19892 29736
rect 19944 29764 19950 29776
rect 20456 29773 20484 29804
rect 20441 29767 20499 29773
rect 20441 29764 20453 29767
rect 19944 29736 20453 29764
rect 19944 29724 19950 29736
rect 20441 29733 20453 29736
rect 20487 29733 20499 29767
rect 20441 29727 20499 29733
rect 20530 29724 20536 29776
rect 20588 29724 20594 29776
rect 19521 29699 19579 29705
rect 19521 29665 19533 29699
rect 19567 29696 19579 29699
rect 20070 29696 20076 29708
rect 19567 29668 20076 29696
rect 19567 29665 19579 29668
rect 19521 29659 19579 29665
rect 20070 29656 20076 29668
rect 20128 29656 20134 29708
rect 20346 29656 20352 29708
rect 20404 29656 20410 29708
rect 20548 29696 20576 29724
rect 20717 29699 20775 29705
rect 20717 29696 20729 29699
rect 20548 29668 20729 29696
rect 20717 29665 20729 29668
rect 20763 29665 20775 29699
rect 20824 29696 20852 29804
rect 20898 29792 20904 29844
rect 20956 29832 20962 29844
rect 21177 29835 21235 29841
rect 21177 29832 21189 29835
rect 20956 29804 21189 29832
rect 20956 29792 20962 29804
rect 21177 29801 21189 29804
rect 21223 29801 21235 29835
rect 21177 29795 21235 29801
rect 21266 29792 21272 29844
rect 21324 29792 21330 29844
rect 21542 29792 21548 29844
rect 21600 29792 21606 29844
rect 22646 29792 22652 29844
rect 22704 29792 22710 29844
rect 23293 29835 23351 29841
rect 23293 29801 23305 29835
rect 23339 29832 23351 29835
rect 23382 29832 23388 29844
rect 23339 29804 23388 29832
rect 23339 29801 23351 29804
rect 23293 29795 23351 29801
rect 23382 29792 23388 29804
rect 23440 29792 23446 29844
rect 23474 29792 23480 29844
rect 23532 29832 23538 29844
rect 23661 29835 23719 29841
rect 23661 29832 23673 29835
rect 23532 29804 23673 29832
rect 23532 29792 23538 29804
rect 23661 29801 23673 29804
rect 23707 29801 23719 29835
rect 23661 29795 23719 29801
rect 24026 29792 24032 29844
rect 24084 29792 24090 29844
rect 24210 29792 24216 29844
rect 24268 29792 24274 29844
rect 24670 29792 24676 29844
rect 24728 29792 24734 29844
rect 24946 29792 24952 29844
rect 25004 29792 25010 29844
rect 25130 29792 25136 29844
rect 25188 29792 25194 29844
rect 25314 29792 25320 29844
rect 25372 29792 25378 29844
rect 25961 29835 26019 29841
rect 25961 29801 25973 29835
rect 26007 29832 26019 29835
rect 26602 29832 26608 29844
rect 26007 29804 26608 29832
rect 26007 29801 26019 29804
rect 25961 29795 26019 29801
rect 21284 29705 21312 29792
rect 21269 29699 21327 29705
rect 20824 29668 21128 29696
rect 20717 29659 20775 29665
rect 20548 29637 20668 29638
rect 19429 29631 19487 29637
rect 19429 29628 19441 29631
rect 19260 29600 19441 29628
rect 19429 29597 19441 29600
rect 19475 29597 19487 29631
rect 19429 29591 19487 29597
rect 20257 29631 20315 29637
rect 20257 29597 20269 29631
rect 20303 29597 20315 29631
rect 20257 29591 20315 29597
rect 20533 29631 20668 29637
rect 20533 29597 20545 29631
rect 20579 29628 20668 29631
rect 20579 29610 20764 29628
rect 20579 29597 20591 29610
rect 20640 29600 20764 29610
rect 20533 29591 20591 29597
rect 17604 29532 18552 29560
rect 20073 29563 20131 29569
rect 17420 29504 17448 29532
rect 20073 29529 20085 29563
rect 20119 29560 20131 29563
rect 20162 29560 20168 29572
rect 20119 29532 20168 29560
rect 20119 29529 20131 29532
rect 20073 29523 20131 29529
rect 20162 29520 20168 29532
rect 20220 29520 20226 29572
rect 17402 29452 17408 29504
rect 17460 29452 17466 29504
rect 20272 29492 20300 29591
rect 20736 29560 20764 29600
rect 20806 29588 20812 29640
rect 20864 29588 20870 29640
rect 20993 29631 21051 29637
rect 20993 29597 21005 29631
rect 21039 29630 21051 29631
rect 21100 29630 21128 29668
rect 21269 29665 21281 29699
rect 21315 29665 21327 29699
rect 21269 29659 21327 29665
rect 21039 29602 21128 29630
rect 21039 29597 21051 29602
rect 20993 29591 21051 29597
rect 21450 29588 21456 29640
rect 21508 29588 21514 29640
rect 21560 29637 21588 29792
rect 23198 29764 23204 29776
rect 23124 29736 23204 29764
rect 23124 29705 23152 29736
rect 23198 29724 23204 29736
rect 23256 29764 23262 29776
rect 24044 29764 24072 29792
rect 23256 29736 24072 29764
rect 23256 29724 23262 29736
rect 23109 29699 23167 29705
rect 23109 29665 23121 29699
rect 23155 29665 23167 29699
rect 23658 29696 23664 29708
rect 23109 29659 23167 29665
rect 23400 29668 23664 29696
rect 21545 29631 21603 29637
rect 21545 29597 21557 29631
rect 21591 29597 21603 29631
rect 21545 29591 21603 29597
rect 22830 29588 22836 29640
rect 22888 29588 22894 29640
rect 23017 29631 23075 29637
rect 23017 29597 23029 29631
rect 23063 29628 23075 29631
rect 23400 29628 23428 29668
rect 23658 29656 23664 29668
rect 23716 29656 23722 29708
rect 23063 29600 23428 29628
rect 23477 29631 23535 29637
rect 23063 29597 23075 29600
rect 23017 29591 23075 29597
rect 23477 29597 23489 29631
rect 23523 29628 23535 29631
rect 23566 29628 23572 29640
rect 23523 29600 23572 29628
rect 23523 29597 23535 29600
rect 23477 29591 23535 29597
rect 23566 29588 23572 29600
rect 23624 29588 23630 29640
rect 21269 29563 21327 29569
rect 21269 29560 21281 29563
rect 20736 29532 21281 29560
rect 21269 29529 21281 29532
rect 21315 29529 21327 29563
rect 21269 29523 21327 29529
rect 20346 29492 20352 29504
rect 20272 29464 20352 29492
rect 20346 29452 20352 29464
rect 20404 29452 20410 29504
rect 23676 29492 23704 29656
rect 23753 29631 23811 29637
rect 23753 29597 23765 29631
rect 23799 29628 23811 29631
rect 24688 29628 24716 29792
rect 25332 29637 25360 29792
rect 25976 29696 26004 29795
rect 26602 29792 26608 29804
rect 26660 29792 26666 29844
rect 27617 29835 27675 29841
rect 27617 29801 27629 29835
rect 27663 29832 27675 29835
rect 27706 29832 27712 29844
rect 27663 29804 27712 29832
rect 27663 29801 27675 29804
rect 27617 29795 27675 29801
rect 27706 29792 27712 29804
rect 27764 29792 27770 29844
rect 27890 29792 27896 29844
rect 27948 29792 27954 29844
rect 27982 29792 27988 29844
rect 28040 29832 28046 29844
rect 28166 29832 28172 29844
rect 28040 29804 28172 29832
rect 28040 29792 28046 29804
rect 28166 29792 28172 29804
rect 28224 29832 28230 29844
rect 28626 29832 28632 29844
rect 28224 29804 28632 29832
rect 28224 29792 28230 29804
rect 28626 29792 28632 29804
rect 28684 29792 28690 29844
rect 31938 29832 31944 29844
rect 31312 29804 31944 29832
rect 27709 29699 27767 29705
rect 25424 29668 26004 29696
rect 27356 29668 27660 29696
rect 25424 29637 25452 29668
rect 24857 29631 24915 29637
rect 24857 29628 24869 29631
rect 23799 29600 23888 29628
rect 23799 29597 23811 29600
rect 23753 29591 23811 29597
rect 23860 29569 23888 29600
rect 24688 29600 24869 29628
rect 23845 29563 23903 29569
rect 23845 29529 23857 29563
rect 23891 29560 23903 29563
rect 24688 29560 24716 29600
rect 24857 29597 24869 29600
rect 24903 29597 24915 29631
rect 24857 29591 24915 29597
rect 25312 29631 25370 29637
rect 25312 29597 25324 29631
rect 25358 29597 25370 29631
rect 25312 29591 25370 29597
rect 25409 29631 25467 29637
rect 25409 29597 25421 29631
rect 25455 29597 25467 29631
rect 25682 29628 25688 29640
rect 25643 29600 25688 29628
rect 25409 29591 25467 29597
rect 25682 29588 25688 29600
rect 25740 29588 25746 29640
rect 25774 29588 25780 29640
rect 25832 29588 25838 29640
rect 26694 29588 26700 29640
rect 26752 29628 26758 29640
rect 27356 29637 27384 29668
rect 27074 29631 27132 29637
rect 27074 29628 27086 29631
rect 26752 29600 27086 29628
rect 26752 29588 26758 29600
rect 27074 29597 27086 29600
rect 27120 29597 27132 29631
rect 27074 29591 27132 29597
rect 27341 29631 27399 29637
rect 27341 29597 27353 29631
rect 27387 29597 27399 29631
rect 27341 29591 27399 29597
rect 27430 29588 27436 29640
rect 27488 29588 27494 29640
rect 27525 29631 27583 29637
rect 27525 29597 27537 29631
rect 27571 29597 27583 29631
rect 27632 29628 27660 29668
rect 27709 29665 27721 29699
rect 27755 29696 27767 29699
rect 27908 29696 27936 29792
rect 29546 29696 29552 29708
rect 27755 29668 27936 29696
rect 29288 29668 29552 29696
rect 27755 29665 27767 29668
rect 27709 29659 27767 29665
rect 29288 29628 29316 29668
rect 29546 29656 29552 29668
rect 29604 29656 29610 29708
rect 29822 29637 29828 29640
rect 27632 29600 29316 29628
rect 29365 29631 29423 29637
rect 27525 29591 27583 29597
rect 29365 29597 29377 29631
rect 29411 29597 29423 29631
rect 29816 29628 29828 29637
rect 29783 29600 29828 29628
rect 29365 29591 29423 29597
rect 29816 29591 29828 29600
rect 23891 29532 24716 29560
rect 23891 29529 23903 29532
rect 23845 29523 23903 29529
rect 25498 29520 25504 29572
rect 25556 29520 25562 29572
rect 25700 29560 25728 29588
rect 27540 29560 27568 29591
rect 25700 29532 27568 29560
rect 24045 29495 24103 29501
rect 24045 29492 24057 29495
rect 23676 29464 24057 29492
rect 24045 29461 24057 29464
rect 24091 29461 24103 29495
rect 27540 29492 27568 29532
rect 28902 29520 28908 29572
rect 28960 29560 28966 29572
rect 29098 29563 29156 29569
rect 29098 29560 29110 29563
rect 28960 29532 29110 29560
rect 28960 29520 28966 29532
rect 29098 29529 29110 29532
rect 29144 29529 29156 29563
rect 29380 29560 29408 29591
rect 29822 29588 29828 29591
rect 29880 29588 29886 29640
rect 31312 29637 31340 29804
rect 31938 29792 31944 29804
rect 31996 29792 32002 29844
rect 31570 29637 31576 29640
rect 31297 29631 31355 29637
rect 31297 29597 31309 29631
rect 31343 29597 31355 29631
rect 31564 29628 31576 29637
rect 31531 29600 31576 29628
rect 31297 29591 31355 29597
rect 31564 29591 31576 29600
rect 31312 29560 31340 29591
rect 31570 29588 31576 29591
rect 31628 29588 31634 29640
rect 29380 29532 31616 29560
rect 29098 29523 29156 29529
rect 31588 29504 31616 29532
rect 27798 29492 27804 29504
rect 27540 29464 27804 29492
rect 24045 29455 24103 29461
rect 27798 29452 27804 29464
rect 27856 29492 27862 29504
rect 27985 29495 28043 29501
rect 27985 29492 27997 29495
rect 27856 29464 27997 29492
rect 27856 29452 27862 29464
rect 27985 29461 27997 29464
rect 28031 29492 28043 29495
rect 28626 29492 28632 29504
rect 28031 29464 28632 29492
rect 28031 29461 28043 29464
rect 27985 29455 28043 29461
rect 28626 29452 28632 29464
rect 28684 29452 28690 29504
rect 30834 29452 30840 29504
rect 30892 29492 30898 29504
rect 30929 29495 30987 29501
rect 30929 29492 30941 29495
rect 30892 29464 30941 29492
rect 30892 29452 30898 29464
rect 30929 29461 30941 29464
rect 30975 29461 30987 29495
rect 30929 29455 30987 29461
rect 31570 29452 31576 29504
rect 31628 29452 31634 29504
rect 32398 29452 32404 29504
rect 32456 29492 32462 29504
rect 32677 29495 32735 29501
rect 32677 29492 32689 29495
rect 32456 29464 32689 29492
rect 32456 29452 32462 29464
rect 32677 29461 32689 29464
rect 32723 29461 32735 29495
rect 32677 29455 32735 29461
rect 1104 29402 35027 29424
rect 1104 29350 9390 29402
rect 9442 29350 9454 29402
rect 9506 29350 9518 29402
rect 9570 29350 9582 29402
rect 9634 29350 9646 29402
rect 9698 29350 17831 29402
rect 17883 29350 17895 29402
rect 17947 29350 17959 29402
rect 18011 29350 18023 29402
rect 18075 29350 18087 29402
rect 18139 29350 26272 29402
rect 26324 29350 26336 29402
rect 26388 29350 26400 29402
rect 26452 29350 26464 29402
rect 26516 29350 26528 29402
rect 26580 29350 34713 29402
rect 34765 29350 34777 29402
rect 34829 29350 34841 29402
rect 34893 29350 34905 29402
rect 34957 29350 34969 29402
rect 35021 29350 35027 29402
rect 1104 29328 35027 29350
rect 18598 29248 18604 29300
rect 18656 29288 18662 29300
rect 19061 29291 19119 29297
rect 19061 29288 19073 29291
rect 18656 29260 19073 29288
rect 18656 29248 18662 29260
rect 19061 29257 19073 29260
rect 19107 29257 19119 29291
rect 19061 29251 19119 29257
rect 19705 29291 19763 29297
rect 19705 29257 19717 29291
rect 19751 29288 19763 29291
rect 20438 29288 20444 29300
rect 19751 29260 20444 29288
rect 19751 29257 19763 29260
rect 19705 29251 19763 29257
rect 20438 29248 20444 29260
rect 20496 29248 20502 29300
rect 20622 29248 20628 29300
rect 20680 29248 20686 29300
rect 20809 29291 20867 29297
rect 20809 29257 20821 29291
rect 20855 29288 20867 29291
rect 20990 29288 20996 29300
rect 20855 29260 20996 29288
rect 20855 29257 20867 29260
rect 20809 29251 20867 29257
rect 20990 29248 20996 29260
rect 21048 29248 21054 29300
rect 22830 29248 22836 29300
rect 22888 29288 22894 29300
rect 23017 29291 23075 29297
rect 23017 29288 23029 29291
rect 22888 29260 23029 29288
rect 22888 29248 22894 29260
rect 23017 29257 23029 29260
rect 23063 29257 23075 29291
rect 23017 29251 23075 29257
rect 26878 29248 26884 29300
rect 26936 29288 26942 29300
rect 28258 29288 28264 29300
rect 26936 29260 28264 29288
rect 26936 29248 26942 29260
rect 28258 29248 28264 29260
rect 28316 29248 28322 29300
rect 28902 29248 28908 29300
rect 28960 29248 28966 29300
rect 17402 29220 17408 29232
rect 17052 29192 17408 29220
rect 17052 29161 17080 29192
rect 17402 29180 17408 29192
rect 17460 29220 17466 29232
rect 17460 29192 17816 29220
rect 17460 29180 17466 29192
rect 17788 29164 17816 29192
rect 19886 29180 19892 29232
rect 19944 29220 19950 29232
rect 20640 29220 20668 29248
rect 23842 29220 23848 29232
rect 19944 29192 20576 29220
rect 20640 29192 21864 29220
rect 19944 29180 19950 29192
rect 17037 29155 17095 29161
rect 17037 29121 17049 29155
rect 17083 29121 17095 29155
rect 17037 29115 17095 29121
rect 17221 29155 17279 29161
rect 17221 29121 17233 29155
rect 17267 29121 17279 29155
rect 17221 29115 17279 29121
rect 16390 29044 16396 29096
rect 16448 29084 16454 29096
rect 17236 29084 17264 29115
rect 17770 29112 17776 29164
rect 17828 29112 17834 29164
rect 20070 29161 20076 29164
rect 19153 29155 19211 29161
rect 19153 29121 19165 29155
rect 19199 29152 19211 29155
rect 19613 29155 19671 29161
rect 19613 29152 19625 29155
rect 19199 29124 19625 29152
rect 19199 29121 19211 29124
rect 19153 29115 19211 29121
rect 19613 29121 19625 29124
rect 19659 29121 19671 29155
rect 19613 29115 19671 29121
rect 19797 29155 19855 29161
rect 19797 29121 19809 29155
rect 19843 29152 19855 29155
rect 20059 29155 20076 29161
rect 20059 29152 20071 29155
rect 19843 29124 20071 29152
rect 19843 29121 19855 29124
rect 19797 29115 19855 29121
rect 20059 29121 20071 29124
rect 20059 29115 20076 29121
rect 18414 29084 18420 29096
rect 16448 29056 18420 29084
rect 16448 29044 16454 29056
rect 18414 29044 18420 29056
rect 18472 29044 18478 29096
rect 19628 29084 19656 29115
rect 20070 29112 20076 29115
rect 20128 29112 20134 29164
rect 20254 29112 20260 29164
rect 20312 29152 20318 29164
rect 20349 29155 20407 29161
rect 20349 29152 20361 29155
rect 20312 29124 20361 29152
rect 20312 29112 20318 29124
rect 20349 29121 20361 29124
rect 20395 29121 20407 29155
rect 20548 29152 20576 29192
rect 20625 29155 20683 29161
rect 20625 29152 20637 29155
rect 20548 29124 20637 29152
rect 20349 29115 20407 29121
rect 20625 29121 20637 29124
rect 20671 29121 20683 29155
rect 20625 29115 20683 29121
rect 20809 29155 20867 29161
rect 20809 29121 20821 29155
rect 20855 29152 20867 29155
rect 20990 29152 20996 29164
rect 20855 29124 20996 29152
rect 20855 29121 20867 29124
rect 20809 29115 20867 29121
rect 20990 29112 20996 29124
rect 21048 29112 21054 29164
rect 21100 29161 21128 29192
rect 21836 29161 21864 29192
rect 23032 29192 23848 29220
rect 23032 29164 23060 29192
rect 23842 29180 23848 29192
rect 23900 29180 23906 29232
rect 28276 29220 28304 29248
rect 28276 29192 28580 29220
rect 21085 29155 21143 29161
rect 21085 29121 21097 29155
rect 21131 29121 21143 29155
rect 21085 29115 21143 29121
rect 21269 29155 21327 29161
rect 21269 29121 21281 29155
rect 21315 29152 21327 29155
rect 21361 29155 21419 29161
rect 21361 29152 21373 29155
rect 21315 29124 21373 29152
rect 21315 29121 21327 29124
rect 21269 29115 21327 29121
rect 21361 29121 21373 29124
rect 21407 29121 21419 29155
rect 21821 29155 21879 29161
rect 21361 29115 21419 29121
rect 21468 29124 21772 29152
rect 19889 29087 19947 29093
rect 19889 29084 19901 29087
rect 19628 29056 19901 29084
rect 19889 29053 19901 29056
rect 19935 29084 19947 29087
rect 20714 29084 20720 29096
rect 19935 29056 20720 29084
rect 19935 29053 19947 29056
rect 19889 29047 19947 29053
rect 20714 29044 20720 29056
rect 20772 29044 20778 29096
rect 20898 29044 20904 29096
rect 20956 29084 20962 29096
rect 21468 29084 21496 29124
rect 20956 29056 21496 29084
rect 20956 29044 20962 29056
rect 21542 29044 21548 29096
rect 21600 29084 21606 29096
rect 21637 29087 21695 29093
rect 21637 29084 21649 29087
rect 21600 29056 21649 29084
rect 21600 29044 21606 29056
rect 21637 29053 21649 29056
rect 21683 29053 21695 29087
rect 21744 29084 21772 29124
rect 21821 29121 21833 29155
rect 21867 29121 21879 29155
rect 21821 29115 21879 29121
rect 22005 29155 22063 29161
rect 22005 29121 22017 29155
rect 22051 29121 22063 29155
rect 22005 29115 22063 29121
rect 22925 29155 22983 29161
rect 22925 29121 22937 29155
rect 22971 29152 22983 29155
rect 23014 29152 23020 29164
rect 22971 29124 23020 29152
rect 22971 29121 22983 29124
rect 22925 29115 22983 29121
rect 22020 29084 22048 29115
rect 23014 29112 23020 29124
rect 23072 29112 23078 29164
rect 23109 29155 23167 29161
rect 23109 29121 23121 29155
rect 23155 29152 23167 29155
rect 23474 29152 23480 29164
rect 23155 29124 23480 29152
rect 23155 29121 23167 29124
rect 23109 29115 23167 29121
rect 23474 29112 23480 29124
rect 23532 29112 23538 29164
rect 25038 29112 25044 29164
rect 25096 29112 25102 29164
rect 28258 29112 28264 29164
rect 28316 29112 28322 29164
rect 28424 29158 28482 29164
rect 28552 29161 28580 29192
rect 28424 29155 28436 29158
rect 28368 29127 28436 29155
rect 21744 29056 22048 29084
rect 21637 29047 21695 29053
rect 20254 28976 20260 29028
rect 20312 28976 20318 29028
rect 20487 29019 20545 29025
rect 20487 28985 20499 29019
rect 20533 29016 20545 29019
rect 20806 29016 20812 29028
rect 20533 28988 20812 29016
rect 20533 28985 20545 28988
rect 20487 28979 20545 28985
rect 20806 28976 20812 28988
rect 20864 29016 20870 29028
rect 21453 29019 21511 29025
rect 21453 29016 21465 29019
rect 20864 28988 21465 29016
rect 20864 28976 20870 28988
rect 21453 28985 21465 28988
rect 21499 29016 21511 29019
rect 21821 29019 21879 29025
rect 21821 29016 21833 29019
rect 21499 28988 21833 29016
rect 21499 28985 21511 28988
rect 21453 28979 21511 28985
rect 21821 28985 21833 28988
rect 21867 28985 21879 29019
rect 28368 29016 28396 29127
rect 28424 29124 28436 29127
rect 28470 29124 28482 29158
rect 28424 29118 28482 29124
rect 28537 29155 28595 29161
rect 28537 29121 28549 29155
rect 28583 29121 28595 29155
rect 28537 29115 28595 29121
rect 28626 29112 28632 29164
rect 28684 29112 28690 29164
rect 31573 29155 31631 29161
rect 31573 29121 31585 29155
rect 31619 29152 31631 29155
rect 32125 29155 32183 29161
rect 32125 29152 32137 29155
rect 31619 29124 32137 29152
rect 31619 29121 31631 29124
rect 31573 29115 31631 29121
rect 32125 29121 32137 29124
rect 32171 29121 32183 29155
rect 32125 29115 32183 29121
rect 32309 29155 32367 29161
rect 32309 29121 32321 29155
rect 32355 29121 32367 29155
rect 32309 29115 32367 29121
rect 31202 29044 31208 29096
rect 31260 29084 31266 29096
rect 32324 29084 32352 29115
rect 31260 29056 32352 29084
rect 31260 29044 31266 29056
rect 32398 29044 32404 29096
rect 32456 29084 32462 29096
rect 32493 29087 32551 29093
rect 32493 29084 32505 29087
rect 32456 29056 32505 29084
rect 32456 29044 32462 29056
rect 32493 29053 32505 29056
rect 32539 29053 32551 29087
rect 32493 29047 32551 29053
rect 28534 29016 28540 29028
rect 28368 28988 28540 29016
rect 21821 28979 21879 28985
rect 28534 28976 28540 28988
rect 28592 28976 28598 29028
rect 17034 28908 17040 28960
rect 17092 28908 17098 28960
rect 21542 28908 21548 28960
rect 21600 28908 21606 28960
rect 25130 28908 25136 28960
rect 25188 28908 25194 28960
rect 31757 28951 31815 28957
rect 31757 28917 31769 28951
rect 31803 28948 31815 28951
rect 31846 28948 31852 28960
rect 31803 28920 31852 28948
rect 31803 28917 31815 28920
rect 31757 28911 31815 28917
rect 31846 28908 31852 28920
rect 31904 28908 31910 28960
rect 1104 28858 34868 28880
rect 1104 28806 5170 28858
rect 5222 28806 5234 28858
rect 5286 28806 5298 28858
rect 5350 28806 5362 28858
rect 5414 28806 5426 28858
rect 5478 28806 13611 28858
rect 13663 28806 13675 28858
rect 13727 28806 13739 28858
rect 13791 28806 13803 28858
rect 13855 28806 13867 28858
rect 13919 28806 22052 28858
rect 22104 28806 22116 28858
rect 22168 28806 22180 28858
rect 22232 28806 22244 28858
rect 22296 28806 22308 28858
rect 22360 28806 30493 28858
rect 30545 28806 30557 28858
rect 30609 28806 30621 28858
rect 30673 28806 30685 28858
rect 30737 28806 30749 28858
rect 30801 28806 34868 28858
rect 1104 28784 34868 28806
rect 16666 28744 16672 28756
rect 16316 28716 16672 28744
rect 16316 28617 16344 28716
rect 16666 28704 16672 28716
rect 16724 28704 16730 28756
rect 17770 28704 17776 28756
rect 17828 28704 17834 28756
rect 17957 28747 18015 28753
rect 17957 28713 17969 28747
rect 18003 28744 18015 28747
rect 18322 28744 18328 28756
rect 18003 28716 18328 28744
rect 18003 28713 18015 28716
rect 17957 28707 18015 28713
rect 18322 28704 18328 28716
rect 18380 28704 18386 28756
rect 18785 28747 18843 28753
rect 18785 28713 18797 28747
rect 18831 28744 18843 28747
rect 18874 28744 18880 28756
rect 18831 28716 18880 28744
rect 18831 28713 18843 28716
rect 18785 28707 18843 28713
rect 18874 28704 18880 28716
rect 18932 28704 18938 28756
rect 20714 28704 20720 28756
rect 20772 28744 20778 28756
rect 21269 28747 21327 28753
rect 21269 28744 21281 28747
rect 20772 28716 21281 28744
rect 20772 28704 20778 28716
rect 21269 28713 21281 28716
rect 21315 28744 21327 28747
rect 21450 28744 21456 28756
rect 21315 28716 21456 28744
rect 21315 28713 21327 28716
rect 21269 28707 21327 28713
rect 21450 28704 21456 28716
rect 21508 28704 21514 28756
rect 23658 28704 23664 28756
rect 23716 28704 23722 28756
rect 23845 28747 23903 28753
rect 23845 28713 23857 28747
rect 23891 28713 23903 28747
rect 23845 28707 23903 28713
rect 24765 28747 24823 28753
rect 24765 28713 24777 28747
rect 24811 28744 24823 28747
rect 24811 28716 25544 28744
rect 24811 28713 24823 28716
rect 24765 28707 24823 28713
rect 17681 28679 17739 28685
rect 17681 28645 17693 28679
rect 17727 28676 17739 28679
rect 17727 28648 18368 28676
rect 17727 28645 17739 28648
rect 17681 28639 17739 28645
rect 16301 28611 16359 28617
rect 16301 28577 16313 28611
rect 16347 28577 16359 28611
rect 16301 28571 16359 28577
rect 18230 28500 18236 28552
rect 18288 28500 18294 28552
rect 18340 28540 18368 28648
rect 20732 28580 21588 28608
rect 18601 28543 18659 28549
rect 18601 28540 18613 28543
rect 18340 28512 18613 28540
rect 16568 28475 16626 28481
rect 16568 28441 16580 28475
rect 16614 28472 16626 28475
rect 16850 28472 16856 28484
rect 16614 28444 16856 28472
rect 16614 28441 16626 28444
rect 16568 28435 16626 28441
rect 16850 28432 16856 28444
rect 16908 28432 16914 28484
rect 18141 28475 18199 28481
rect 18141 28441 18153 28475
rect 18187 28472 18199 28475
rect 18340 28472 18368 28512
rect 18601 28509 18613 28512
rect 18647 28540 18659 28543
rect 18690 28540 18696 28552
rect 18647 28512 18696 28540
rect 18647 28509 18659 28512
rect 18601 28503 18659 28509
rect 18690 28500 18696 28512
rect 18748 28500 18754 28552
rect 20533 28543 20591 28549
rect 20533 28509 20545 28543
rect 20579 28540 20591 28543
rect 20622 28540 20628 28552
rect 20579 28512 20628 28540
rect 20579 28509 20591 28512
rect 20533 28503 20591 28509
rect 20622 28500 20628 28512
rect 20680 28500 20686 28552
rect 20732 28549 20760 28580
rect 21560 28552 21588 28580
rect 20717 28543 20775 28549
rect 20717 28509 20729 28543
rect 20763 28509 20775 28543
rect 20717 28503 20775 28509
rect 20809 28543 20867 28549
rect 20809 28509 20821 28543
rect 20855 28509 20867 28543
rect 20809 28503 20867 28509
rect 20901 28543 20959 28549
rect 20901 28509 20913 28543
rect 20947 28540 20959 28543
rect 21450 28540 21456 28552
rect 20947 28512 21456 28540
rect 20947 28509 20959 28512
rect 20901 28503 20959 28509
rect 18187 28444 18368 28472
rect 18187 28441 18199 28444
rect 18141 28435 18199 28441
rect 18414 28432 18420 28484
rect 18472 28432 18478 28484
rect 18509 28475 18567 28481
rect 18509 28441 18521 28475
rect 18555 28441 18567 28475
rect 20824 28472 20852 28503
rect 21450 28500 21456 28512
rect 21508 28500 21514 28552
rect 21542 28500 21548 28552
rect 21600 28500 21606 28552
rect 22649 28543 22707 28549
rect 22649 28509 22661 28543
rect 22695 28509 22707 28543
rect 22649 28503 22707 28509
rect 21082 28472 21088 28484
rect 20824 28444 21088 28472
rect 18509 28435 18567 28441
rect 17494 28364 17500 28416
rect 17552 28404 17558 28416
rect 17931 28407 17989 28413
rect 17931 28404 17943 28407
rect 17552 28376 17943 28404
rect 17552 28364 17558 28376
rect 17931 28373 17943 28376
rect 17977 28373 17989 28407
rect 18524 28404 18552 28435
rect 21082 28432 21088 28444
rect 21140 28432 21146 28484
rect 21177 28475 21235 28481
rect 21177 28441 21189 28475
rect 21223 28472 21235 28475
rect 22382 28475 22440 28481
rect 22382 28472 22394 28475
rect 21223 28444 22394 28472
rect 21223 28441 21235 28444
rect 21177 28435 21235 28441
rect 22382 28441 22394 28444
rect 22428 28441 22440 28475
rect 22664 28472 22692 28503
rect 23014 28500 23020 28552
rect 23072 28500 23078 28552
rect 23201 28543 23259 28549
rect 23201 28509 23213 28543
rect 23247 28540 23259 28543
rect 23676 28540 23704 28704
rect 23860 28676 23888 28707
rect 25038 28676 25044 28688
rect 23860 28648 25044 28676
rect 25038 28636 25044 28648
rect 25096 28636 25102 28688
rect 25130 28636 25136 28688
rect 25188 28636 25194 28688
rect 25148 28608 25176 28636
rect 25516 28620 25544 28716
rect 25774 28704 25780 28756
rect 25832 28744 25838 28756
rect 25869 28747 25927 28753
rect 25869 28744 25881 28747
rect 25832 28716 25881 28744
rect 25832 28704 25838 28716
rect 25869 28713 25881 28716
rect 25915 28713 25927 28747
rect 25869 28707 25927 28713
rect 27890 28704 27896 28756
rect 27948 28704 27954 28756
rect 25148 28580 25360 28608
rect 25332 28552 25360 28580
rect 25498 28568 25504 28620
rect 25556 28568 25562 28620
rect 27525 28611 27583 28617
rect 27525 28577 27537 28611
rect 27571 28608 27583 28611
rect 27706 28608 27712 28620
rect 27571 28580 27712 28608
rect 27571 28577 27583 28580
rect 27525 28571 27583 28577
rect 27706 28568 27712 28580
rect 27764 28608 27770 28620
rect 27908 28608 27936 28704
rect 27764 28580 27936 28608
rect 28077 28611 28135 28617
rect 27764 28568 27770 28580
rect 28077 28577 28089 28611
rect 28123 28608 28135 28611
rect 28994 28608 29000 28620
rect 28123 28580 29000 28608
rect 28123 28577 28135 28580
rect 28077 28571 28135 28577
rect 28994 28568 29000 28580
rect 29052 28568 29058 28620
rect 24673 28543 24731 28549
rect 24673 28540 24685 28543
rect 23247 28512 23704 28540
rect 24044 28512 24685 28540
rect 23247 28509 23259 28512
rect 23201 28503 23259 28509
rect 24044 28484 24072 28512
rect 24673 28509 24685 28512
rect 24719 28509 24731 28543
rect 24673 28503 24731 28509
rect 25130 28500 25136 28552
rect 25188 28500 25194 28552
rect 25314 28500 25320 28552
rect 25372 28500 25378 28552
rect 25409 28543 25467 28549
rect 25409 28509 25421 28543
rect 25455 28509 25467 28543
rect 25409 28503 25467 28509
rect 22664 28444 23244 28472
rect 22382 28435 22440 28441
rect 23216 28416 23244 28444
rect 24026 28432 24032 28484
rect 24084 28432 24090 28484
rect 25424 28472 25452 28503
rect 25682 28500 25688 28552
rect 25740 28500 25746 28552
rect 27249 28543 27307 28549
rect 27249 28540 27261 28543
rect 27172 28512 27261 28540
rect 25498 28472 25504 28484
rect 25424 28444 25504 28472
rect 25498 28432 25504 28444
rect 25556 28432 25562 28484
rect 27172 28416 27200 28512
rect 27249 28509 27261 28512
rect 27295 28509 27307 28543
rect 27249 28503 27307 28509
rect 27338 28500 27344 28552
rect 27396 28500 27402 28552
rect 27801 28543 27859 28549
rect 27801 28540 27813 28543
rect 27632 28512 27813 28540
rect 27632 28416 27660 28512
rect 27801 28509 27813 28512
rect 27847 28509 27859 28543
rect 27801 28503 27859 28509
rect 27893 28543 27951 28549
rect 27893 28509 27905 28543
rect 27939 28509 27951 28543
rect 27893 28503 27951 28509
rect 30009 28543 30067 28549
rect 30009 28509 30021 28543
rect 30055 28540 30067 28543
rect 31018 28540 31024 28552
rect 30055 28512 31024 28540
rect 30055 28509 30067 28512
rect 30009 28503 30067 28509
rect 27908 28416 27936 28503
rect 31018 28500 31024 28512
rect 31076 28540 31082 28552
rect 31846 28549 31852 28552
rect 31573 28543 31631 28549
rect 31573 28540 31585 28543
rect 31076 28512 31585 28540
rect 31076 28500 31082 28512
rect 31573 28509 31585 28512
rect 31619 28509 31631 28543
rect 31840 28540 31852 28549
rect 31807 28512 31852 28540
rect 31573 28503 31631 28509
rect 31840 28503 31852 28512
rect 31846 28500 31852 28503
rect 31904 28500 31910 28552
rect 30276 28475 30334 28481
rect 30276 28441 30288 28475
rect 30322 28472 30334 28475
rect 30374 28472 30380 28484
rect 30322 28444 30380 28472
rect 30322 28441 30334 28444
rect 30276 28435 30334 28441
rect 30374 28432 30380 28444
rect 30432 28432 30438 28484
rect 18598 28404 18604 28416
rect 18524 28376 18604 28404
rect 17931 28367 17989 28373
rect 18598 28364 18604 28376
rect 18656 28364 18662 28416
rect 23106 28364 23112 28416
rect 23164 28364 23170 28416
rect 23198 28364 23204 28416
rect 23256 28364 23262 28416
rect 23842 28413 23848 28416
rect 23819 28407 23848 28413
rect 23819 28373 23831 28407
rect 23819 28367 23848 28373
rect 23842 28364 23848 28367
rect 23900 28364 23906 28416
rect 27154 28364 27160 28416
rect 27212 28364 27218 28416
rect 27522 28364 27528 28416
rect 27580 28364 27586 28416
rect 27614 28364 27620 28416
rect 27672 28364 27678 28416
rect 27890 28364 27896 28416
rect 27948 28364 27954 28416
rect 28074 28364 28080 28416
rect 28132 28364 28138 28416
rect 31386 28364 31392 28416
rect 31444 28364 31450 28416
rect 32122 28364 32128 28416
rect 32180 28404 32186 28416
rect 32953 28407 33011 28413
rect 32953 28404 32965 28407
rect 32180 28376 32965 28404
rect 32180 28364 32186 28376
rect 32953 28373 32965 28376
rect 32999 28373 33011 28407
rect 32953 28367 33011 28373
rect 1104 28314 35027 28336
rect 1104 28262 9390 28314
rect 9442 28262 9454 28314
rect 9506 28262 9518 28314
rect 9570 28262 9582 28314
rect 9634 28262 9646 28314
rect 9698 28262 17831 28314
rect 17883 28262 17895 28314
rect 17947 28262 17959 28314
rect 18011 28262 18023 28314
rect 18075 28262 18087 28314
rect 18139 28262 26272 28314
rect 26324 28262 26336 28314
rect 26388 28262 26400 28314
rect 26452 28262 26464 28314
rect 26516 28262 26528 28314
rect 26580 28262 34713 28314
rect 34765 28262 34777 28314
rect 34829 28262 34841 28314
rect 34893 28262 34905 28314
rect 34957 28262 34969 28314
rect 35021 28262 35027 28314
rect 1104 28240 35027 28262
rect 16850 28160 16856 28212
rect 16908 28160 16914 28212
rect 18414 28160 18420 28212
rect 18472 28200 18478 28212
rect 18601 28203 18659 28209
rect 18601 28200 18613 28203
rect 18472 28172 18613 28200
rect 18472 28160 18478 28172
rect 18601 28169 18613 28172
rect 18647 28169 18659 28203
rect 18601 28163 18659 28169
rect 23658 28160 23664 28212
rect 23716 28200 23722 28212
rect 24026 28200 24032 28212
rect 23716 28172 24032 28200
rect 23716 28160 23722 28172
rect 24026 28160 24032 28172
rect 24084 28160 24090 28212
rect 25038 28160 25044 28212
rect 25096 28200 25102 28212
rect 25133 28203 25191 28209
rect 25133 28200 25145 28203
rect 25096 28172 25145 28200
rect 25096 28160 25102 28172
rect 25133 28169 25145 28172
rect 25179 28169 25191 28203
rect 25133 28163 25191 28169
rect 25498 28160 25504 28212
rect 25556 28200 25562 28212
rect 26789 28203 26847 28209
rect 26789 28200 26801 28203
rect 25556 28172 26801 28200
rect 25556 28160 25562 28172
rect 26789 28169 26801 28172
rect 26835 28169 26847 28203
rect 26789 28163 26847 28169
rect 17405 28135 17463 28141
rect 17405 28101 17417 28135
rect 17451 28132 17463 28135
rect 17451 28104 17908 28132
rect 17451 28101 17463 28104
rect 17405 28095 17463 28101
rect 17034 28024 17040 28076
rect 17092 28024 17098 28076
rect 17221 28067 17279 28073
rect 17221 28033 17233 28067
rect 17267 28064 17279 28067
rect 17420 28064 17448 28095
rect 17267 28036 17448 28064
rect 17267 28033 17279 28036
rect 17221 28027 17279 28033
rect 17494 28024 17500 28076
rect 17552 28064 17558 28076
rect 17880 28073 17908 28104
rect 22296 28104 23336 28132
rect 17589 28067 17647 28073
rect 17589 28064 17601 28067
rect 17552 28036 17601 28064
rect 17552 28024 17558 28036
rect 17589 28033 17601 28036
rect 17635 28033 17647 28067
rect 17589 28027 17647 28033
rect 17865 28067 17923 28073
rect 17865 28033 17877 28067
rect 17911 28033 17923 28067
rect 17865 28027 17923 28033
rect 18049 28067 18107 28073
rect 18049 28033 18061 28067
rect 18095 28064 18107 28067
rect 18138 28064 18144 28076
rect 18095 28036 18144 28064
rect 18095 28033 18107 28036
rect 18049 28027 18107 28033
rect 18138 28024 18144 28036
rect 18196 28024 18202 28076
rect 18233 28067 18291 28073
rect 18233 28033 18245 28067
rect 18279 28064 18291 28067
rect 18322 28064 18328 28076
rect 18279 28036 18328 28064
rect 18279 28033 18291 28036
rect 18233 28027 18291 28033
rect 17313 27999 17371 28005
rect 17313 27965 17325 27999
rect 17359 27965 17371 27999
rect 17313 27959 17371 27965
rect 17773 27999 17831 28005
rect 17773 27965 17785 27999
rect 17819 27996 17831 27999
rect 17954 27996 17960 28008
rect 17819 27968 17960 27996
rect 17819 27965 17831 27968
rect 17773 27959 17831 27965
rect 17328 27928 17356 27959
rect 17954 27956 17960 27968
rect 18012 27996 18018 28008
rect 18248 27996 18276 28027
rect 18322 28024 18328 28036
rect 18380 28024 18386 28076
rect 18417 28067 18475 28073
rect 18417 28033 18429 28067
rect 18463 28064 18475 28067
rect 18966 28064 18972 28076
rect 18463 28036 18972 28064
rect 18463 28033 18475 28036
rect 18417 28027 18475 28033
rect 18966 28024 18972 28036
rect 19024 28024 19030 28076
rect 19334 28024 19340 28076
rect 19392 28024 19398 28076
rect 22296 28073 22324 28104
rect 23308 28076 23336 28104
rect 22281 28067 22339 28073
rect 22281 28033 22293 28067
rect 22327 28033 22339 28067
rect 22281 28027 22339 28033
rect 22548 28067 22606 28073
rect 22548 28033 22560 28067
rect 22594 28064 22606 28067
rect 22922 28064 22928 28076
rect 22594 28036 22928 28064
rect 22594 28033 22606 28036
rect 22548 28027 22606 28033
rect 22922 28024 22928 28036
rect 22980 28024 22986 28076
rect 23290 28024 23296 28076
rect 23348 28064 23354 28076
rect 23566 28064 23572 28076
rect 23348 28036 23572 28064
rect 23348 28024 23354 28036
rect 23566 28024 23572 28036
rect 23624 28064 23630 28076
rect 24026 28073 24032 28076
rect 23753 28067 23811 28073
rect 23753 28064 23765 28067
rect 23624 28036 23765 28064
rect 23624 28024 23630 28036
rect 23753 28033 23765 28036
rect 23799 28033 23811 28067
rect 23753 28027 23811 28033
rect 24020 28027 24032 28073
rect 24026 28024 24032 28027
rect 24084 28024 24090 28076
rect 25676 28067 25734 28073
rect 25676 28033 25688 28067
rect 25722 28064 25734 28067
rect 25958 28064 25964 28076
rect 25722 28036 25964 28064
rect 25722 28033 25734 28036
rect 25676 28027 25734 28033
rect 25958 28024 25964 28036
rect 26016 28024 26022 28076
rect 26804 28064 26832 28163
rect 27522 28160 27528 28212
rect 27580 28160 27586 28212
rect 27706 28160 27712 28212
rect 27764 28160 27770 28212
rect 28169 28203 28227 28209
rect 28169 28169 28181 28203
rect 28215 28200 28227 28203
rect 28810 28200 28816 28212
rect 28215 28172 28816 28200
rect 28215 28169 28227 28172
rect 28169 28163 28227 28169
rect 28810 28160 28816 28172
rect 28868 28160 28874 28212
rect 28994 28160 29000 28212
rect 29052 28160 29058 28212
rect 30374 28160 30380 28212
rect 30432 28160 30438 28212
rect 31202 28200 31208 28212
rect 30852 28172 31208 28200
rect 27154 28064 27160 28076
rect 26804 28036 27160 28064
rect 27154 28024 27160 28036
rect 27212 28024 27218 28076
rect 27540 28064 27568 28160
rect 27724 28132 27752 28160
rect 29012 28132 29040 28160
rect 27724 28104 28948 28132
rect 29012 28104 29408 28132
rect 28920 28073 28948 28104
rect 27709 28067 27767 28073
rect 27709 28064 27721 28067
rect 27540 28036 27721 28064
rect 27709 28033 27721 28036
rect 27755 28033 27767 28067
rect 27985 28067 28043 28073
rect 27985 28064 27997 28067
rect 27709 28027 27767 28033
rect 27816 28036 27997 28064
rect 18012 27968 18276 27996
rect 18012 27956 18018 27968
rect 18690 27956 18696 28008
rect 18748 27956 18754 28008
rect 19429 27999 19487 28005
rect 19429 27965 19441 27999
rect 19475 27996 19487 27999
rect 20070 27996 20076 28008
rect 19475 27968 20076 27996
rect 19475 27965 19487 27968
rect 19429 27959 19487 27965
rect 20070 27956 20076 27968
rect 20128 27956 20134 28008
rect 25406 27956 25412 28008
rect 25464 27956 25470 28008
rect 27249 27999 27307 28005
rect 27249 27965 27261 27999
rect 27295 27965 27307 27999
rect 27249 27959 27307 27965
rect 18708 27928 18736 27956
rect 17328 27900 18736 27928
rect 19705 27931 19763 27937
rect 19705 27897 19717 27931
rect 19751 27928 19763 27931
rect 20254 27928 20260 27940
rect 19751 27900 20260 27928
rect 19751 27897 19763 27900
rect 19705 27891 19763 27897
rect 20254 27888 20260 27900
rect 20312 27888 20318 27940
rect 18046 27820 18052 27872
rect 18104 27820 18110 27872
rect 27264 27860 27292 27959
rect 27614 27956 27620 28008
rect 27672 27996 27678 28008
rect 27816 27996 27844 28036
rect 27985 28033 27997 28036
rect 28031 28064 28043 28067
rect 28445 28067 28503 28073
rect 28445 28064 28457 28067
rect 28031 28036 28457 28064
rect 28031 28033 28043 28036
rect 27985 28027 28043 28033
rect 28445 28033 28457 28036
rect 28491 28033 28503 28067
rect 28445 28027 28503 28033
rect 28905 28067 28963 28073
rect 28905 28033 28917 28067
rect 28951 28033 28963 28067
rect 28905 28027 28963 28033
rect 28994 28024 29000 28076
rect 29052 28064 29058 28076
rect 29089 28067 29147 28073
rect 29089 28064 29101 28067
rect 29052 28036 29101 28064
rect 29052 28024 29058 28036
rect 29089 28033 29101 28036
rect 29135 28033 29147 28067
rect 29089 28027 29147 28033
rect 29178 28024 29184 28076
rect 29236 28024 29242 28076
rect 29380 28073 29408 28104
rect 30852 28073 30880 28172
rect 31202 28160 31208 28172
rect 31260 28160 31266 28212
rect 31754 28160 31760 28212
rect 31812 28200 31818 28212
rect 32309 28203 32367 28209
rect 32309 28200 32321 28203
rect 31812 28172 32321 28200
rect 31812 28160 31818 28172
rect 32309 28169 32321 28172
rect 32355 28200 32367 28203
rect 32398 28200 32404 28212
rect 32355 28172 32404 28200
rect 32355 28169 32367 28172
rect 32309 28163 32367 28169
rect 32398 28160 32404 28172
rect 32456 28160 32462 28212
rect 31386 28132 31392 28144
rect 30944 28104 31392 28132
rect 30944 28076 30972 28104
rect 31386 28092 31392 28104
rect 31444 28132 31450 28144
rect 31481 28135 31539 28141
rect 31481 28132 31493 28135
rect 31444 28104 31493 28132
rect 31444 28092 31450 28104
rect 31481 28101 31493 28104
rect 31527 28132 31539 28135
rect 32493 28135 32551 28141
rect 32493 28132 32505 28135
rect 31527 28104 32505 28132
rect 31527 28101 31539 28104
rect 31481 28095 31539 28101
rect 32493 28101 32505 28104
rect 32539 28101 32551 28135
rect 32493 28095 32551 28101
rect 29365 28067 29423 28073
rect 29365 28033 29377 28067
rect 29411 28033 29423 28067
rect 29365 28027 29423 28033
rect 30561 28067 30619 28073
rect 30561 28033 30573 28067
rect 30607 28064 30619 28067
rect 30653 28067 30711 28073
rect 30653 28064 30665 28067
rect 30607 28036 30665 28064
rect 30607 28033 30619 28036
rect 30561 28027 30619 28033
rect 30653 28033 30665 28036
rect 30699 28033 30711 28067
rect 30653 28027 30711 28033
rect 30837 28067 30895 28073
rect 30837 28033 30849 28067
rect 30883 28033 30895 28067
rect 30837 28027 30895 28033
rect 30926 28024 30932 28076
rect 30984 28024 30990 28076
rect 31021 28067 31079 28073
rect 31021 28033 31033 28067
rect 31067 28033 31079 28067
rect 31021 28027 31079 28033
rect 27672 27968 27844 27996
rect 27672 27956 27678 27968
rect 27890 27956 27896 28008
rect 27948 27996 27954 28008
rect 28537 27999 28595 28005
rect 28537 27996 28549 27999
rect 27948 27968 28549 27996
rect 27948 27956 27954 27968
rect 28537 27965 28549 27968
rect 28583 27996 28595 27999
rect 29273 27999 29331 28005
rect 29273 27996 29285 27999
rect 28583 27968 29285 27996
rect 28583 27965 28595 27968
rect 28537 27959 28595 27965
rect 29273 27965 29285 27968
rect 29319 27965 29331 27999
rect 31036 27996 31064 28027
rect 31110 28024 31116 28076
rect 31168 28024 31174 28076
rect 31757 28067 31815 28073
rect 31757 28064 31769 28067
rect 31588 28036 31769 28064
rect 31588 27996 31616 28036
rect 31757 28033 31769 28036
rect 31803 28064 31815 28067
rect 32122 28064 32128 28076
rect 31803 28036 32128 28064
rect 31803 28033 31815 28036
rect 31757 28027 31815 28033
rect 32122 28024 32128 28036
rect 32180 28024 32186 28076
rect 32398 28024 32404 28076
rect 32456 28024 32462 28076
rect 31036 27968 31616 27996
rect 31665 27999 31723 28005
rect 29273 27959 29331 27965
rect 31665 27965 31677 27999
rect 31711 27996 31723 27999
rect 32416 27996 32444 28024
rect 31711 27968 32444 27996
rect 31711 27965 31723 27968
rect 31665 27959 31723 27965
rect 27430 27888 27436 27940
rect 27488 27928 27494 27940
rect 27525 27931 27583 27937
rect 27525 27928 27537 27931
rect 27488 27900 27537 27928
rect 27488 27888 27494 27900
rect 27525 27897 27537 27900
rect 27571 27928 27583 27931
rect 27801 27931 27859 27937
rect 27801 27928 27813 27931
rect 27571 27900 27813 27928
rect 27571 27897 27583 27900
rect 27525 27891 27583 27897
rect 27801 27897 27813 27900
rect 27847 27928 27859 27931
rect 27982 27928 27988 27940
rect 27847 27900 27988 27928
rect 27847 27897 27859 27900
rect 27801 27891 27859 27897
rect 27982 27888 27988 27900
rect 28040 27888 28046 27940
rect 28813 27931 28871 27937
rect 28813 27897 28825 27931
rect 28859 27928 28871 27931
rect 29362 27928 29368 27940
rect 28859 27900 29368 27928
rect 28859 27897 28871 27900
rect 28813 27891 28871 27897
rect 29362 27888 29368 27900
rect 29420 27888 29426 27940
rect 27706 27860 27712 27872
rect 27264 27832 27712 27860
rect 27706 27820 27712 27832
rect 27764 27820 27770 27872
rect 31294 27820 31300 27872
rect 31352 27820 31358 27872
rect 31662 27820 31668 27872
rect 31720 27820 31726 27872
rect 31941 27863 31999 27869
rect 31941 27829 31953 27863
rect 31987 27860 31999 27863
rect 32490 27860 32496 27872
rect 31987 27832 32496 27860
rect 31987 27829 31999 27832
rect 31941 27823 31999 27829
rect 32490 27820 32496 27832
rect 32548 27820 32554 27872
rect 32677 27863 32735 27869
rect 32677 27829 32689 27863
rect 32723 27860 32735 27863
rect 32766 27860 32772 27872
rect 32723 27832 32772 27860
rect 32723 27829 32735 27832
rect 32677 27823 32735 27829
rect 32766 27820 32772 27832
rect 32824 27820 32830 27872
rect 1104 27770 34868 27792
rect 1104 27718 5170 27770
rect 5222 27718 5234 27770
rect 5286 27718 5298 27770
rect 5350 27718 5362 27770
rect 5414 27718 5426 27770
rect 5478 27718 13611 27770
rect 13663 27718 13675 27770
rect 13727 27718 13739 27770
rect 13791 27718 13803 27770
rect 13855 27718 13867 27770
rect 13919 27718 22052 27770
rect 22104 27718 22116 27770
rect 22168 27718 22180 27770
rect 22232 27718 22244 27770
rect 22296 27718 22308 27770
rect 22360 27718 30493 27770
rect 30545 27718 30557 27770
rect 30609 27718 30621 27770
rect 30673 27718 30685 27770
rect 30737 27718 30749 27770
rect 30801 27718 34868 27770
rect 1104 27696 34868 27718
rect 17954 27616 17960 27668
rect 18012 27616 18018 27668
rect 18138 27616 18144 27668
rect 18196 27656 18202 27668
rect 18233 27659 18291 27665
rect 18233 27656 18245 27659
rect 18196 27628 18245 27656
rect 18196 27616 18202 27628
rect 18233 27625 18245 27628
rect 18279 27625 18291 27659
rect 21082 27656 21088 27668
rect 18233 27619 18291 27625
rect 19812 27628 21088 27656
rect 18046 27548 18052 27600
rect 18104 27548 18110 27600
rect 18064 27520 18092 27548
rect 17604 27492 18092 27520
rect 18325 27523 18383 27529
rect 16577 27455 16635 27461
rect 16577 27421 16589 27455
rect 16623 27452 16635 27455
rect 16666 27452 16672 27464
rect 16623 27424 16672 27452
rect 16623 27421 16635 27424
rect 16577 27415 16635 27421
rect 16666 27412 16672 27424
rect 16724 27412 16730 27464
rect 16844 27455 16902 27461
rect 16844 27421 16856 27455
rect 16890 27452 16902 27455
rect 17604 27452 17632 27492
rect 18325 27489 18337 27523
rect 18371 27520 18383 27523
rect 18874 27520 18880 27532
rect 18371 27492 18880 27520
rect 18371 27489 18383 27492
rect 18325 27483 18383 27489
rect 18874 27480 18880 27492
rect 18932 27480 18938 27532
rect 16890 27424 17632 27452
rect 16890 27421 16902 27424
rect 16844 27415 16902 27421
rect 17954 27412 17960 27464
rect 18012 27452 18018 27464
rect 19812 27461 19840 27628
rect 21082 27616 21088 27628
rect 21140 27656 21146 27668
rect 21818 27656 21824 27668
rect 21140 27628 21824 27656
rect 21140 27616 21146 27628
rect 21818 27616 21824 27628
rect 21876 27616 21882 27668
rect 22922 27616 22928 27668
rect 22980 27616 22986 27668
rect 24026 27616 24032 27668
rect 24084 27656 24090 27668
rect 24213 27659 24271 27665
rect 24213 27656 24225 27659
rect 24084 27628 24225 27656
rect 24084 27616 24090 27628
rect 24213 27625 24225 27628
rect 24259 27625 24271 27659
rect 25038 27656 25044 27668
rect 24213 27619 24271 27625
rect 24688 27628 25044 27656
rect 20622 27588 20628 27600
rect 20088 27560 20628 27588
rect 20088 27461 20116 27560
rect 20622 27548 20628 27560
rect 20680 27548 20686 27600
rect 23750 27548 23756 27600
rect 23808 27588 23814 27600
rect 24581 27591 24639 27597
rect 24581 27588 24593 27591
rect 23808 27560 24593 27588
rect 23808 27548 23814 27560
rect 24581 27557 24593 27560
rect 24627 27557 24639 27591
rect 24581 27551 24639 27557
rect 20548 27492 20852 27520
rect 18049 27455 18107 27461
rect 18049 27452 18061 27455
rect 18012 27424 18061 27452
rect 18012 27412 18018 27424
rect 18049 27421 18061 27424
rect 18095 27421 18107 27455
rect 18049 27415 18107 27421
rect 18141 27455 18199 27461
rect 18141 27421 18153 27455
rect 18187 27452 18199 27455
rect 19061 27455 19119 27461
rect 18187 27424 18552 27452
rect 18187 27421 18199 27424
rect 18141 27415 18199 27421
rect 18064 27384 18092 27415
rect 18414 27384 18420 27396
rect 18064 27356 18420 27384
rect 18414 27344 18420 27356
rect 18472 27344 18478 27396
rect 17494 27276 17500 27328
rect 17552 27316 17558 27328
rect 18524 27316 18552 27424
rect 19061 27421 19073 27455
rect 19107 27452 19119 27455
rect 19705 27455 19763 27461
rect 19705 27452 19717 27455
rect 19107 27424 19717 27452
rect 19107 27421 19119 27424
rect 19061 27415 19119 27421
rect 19352 27328 19380 27424
rect 19705 27421 19717 27424
rect 19751 27421 19763 27455
rect 19705 27415 19763 27421
rect 19797 27455 19855 27461
rect 19797 27421 19809 27455
rect 19843 27421 19855 27455
rect 19797 27415 19855 27421
rect 19889 27455 19947 27461
rect 19889 27421 19901 27455
rect 19935 27421 19947 27455
rect 19889 27415 19947 27421
rect 20073 27455 20131 27461
rect 20073 27421 20085 27455
rect 20119 27421 20131 27455
rect 20073 27415 20131 27421
rect 19904 27384 19932 27415
rect 20254 27412 20260 27464
rect 20312 27412 20318 27464
rect 20349 27455 20407 27461
rect 20349 27421 20361 27455
rect 20395 27421 20407 27455
rect 20548 27452 20576 27492
rect 20824 27461 20852 27492
rect 20990 27480 20996 27532
rect 21048 27480 21054 27532
rect 23293 27523 23351 27529
rect 23293 27489 23305 27523
rect 23339 27520 23351 27523
rect 23569 27523 23627 27529
rect 23569 27520 23581 27523
rect 23339 27492 23581 27520
rect 23339 27489 23351 27492
rect 23293 27483 23351 27489
rect 23569 27489 23581 27492
rect 23615 27520 23627 27523
rect 24397 27523 24455 27529
rect 24397 27520 24409 27523
rect 23615 27492 24072 27520
rect 23615 27489 23627 27492
rect 23569 27483 23627 27489
rect 20609 27455 20667 27461
rect 20609 27452 20621 27455
rect 20548 27424 20621 27452
rect 20349 27415 20407 27421
rect 20609 27421 20621 27424
rect 20655 27421 20667 27455
rect 20609 27415 20667 27421
rect 20717 27455 20775 27461
rect 20717 27421 20729 27455
rect 20763 27421 20775 27455
rect 20717 27415 20775 27421
rect 20809 27455 20867 27461
rect 20809 27421 20821 27455
rect 20855 27452 20867 27455
rect 21082 27452 21088 27464
rect 20855 27424 21088 27452
rect 20855 27421 20867 27424
rect 20809 27415 20867 27421
rect 20165 27387 20223 27393
rect 20165 27384 20177 27387
rect 19904 27356 20177 27384
rect 20165 27353 20177 27356
rect 20211 27353 20223 27387
rect 20165 27347 20223 27353
rect 17552 27288 18552 27316
rect 17552 27276 17558 27288
rect 18966 27276 18972 27328
rect 19024 27276 19030 27328
rect 19334 27276 19340 27328
rect 19392 27276 19398 27328
rect 19426 27276 19432 27328
rect 19484 27276 19490 27328
rect 20272 27316 20300 27412
rect 20364 27384 20392 27415
rect 20438 27384 20444 27396
rect 20364 27356 20444 27384
rect 20438 27344 20444 27356
rect 20496 27344 20502 27396
rect 20732 27384 20760 27415
rect 21082 27412 21088 27424
rect 21140 27412 21146 27464
rect 23106 27412 23112 27464
rect 23164 27412 23170 27464
rect 23385 27455 23443 27461
rect 23385 27421 23397 27455
rect 23431 27452 23443 27455
rect 23658 27452 23664 27464
rect 23431 27424 23664 27452
rect 23431 27421 23443 27424
rect 23385 27415 23443 27421
rect 23658 27412 23664 27424
rect 23716 27412 23722 27464
rect 24044 27461 24072 27492
rect 24136 27492 24409 27520
rect 23753 27455 23811 27461
rect 23753 27421 23765 27455
rect 23799 27421 23811 27455
rect 23753 27415 23811 27421
rect 23937 27455 23995 27461
rect 23937 27421 23949 27455
rect 23983 27421 23995 27455
rect 23937 27415 23995 27421
rect 24029 27455 24087 27461
rect 24029 27421 24041 27455
rect 24075 27421 24087 27455
rect 24029 27415 24087 27421
rect 20548 27356 20760 27384
rect 20346 27316 20352 27328
rect 20272 27288 20352 27316
rect 20346 27276 20352 27288
rect 20404 27316 20410 27328
rect 20548 27325 20576 27356
rect 23768 27328 23796 27415
rect 20533 27319 20591 27325
rect 20533 27316 20545 27319
rect 20404 27288 20545 27316
rect 20404 27276 20410 27288
rect 20533 27285 20545 27288
rect 20579 27285 20591 27319
rect 20533 27279 20591 27285
rect 20806 27276 20812 27328
rect 20864 27316 20870 27328
rect 20993 27319 21051 27325
rect 20993 27316 21005 27319
rect 20864 27288 21005 27316
rect 20864 27276 20870 27288
rect 20993 27285 21005 27288
rect 21039 27285 21051 27319
rect 20993 27279 21051 27285
rect 23750 27276 23756 27328
rect 23808 27276 23814 27328
rect 23952 27316 23980 27415
rect 24136 27396 24164 27492
rect 24397 27489 24409 27492
rect 24443 27489 24455 27523
rect 24397 27483 24455 27489
rect 24688 27461 24716 27628
rect 25038 27616 25044 27628
rect 25096 27616 25102 27668
rect 25130 27616 25136 27668
rect 25188 27656 25194 27668
rect 25225 27659 25283 27665
rect 25225 27656 25237 27659
rect 25188 27628 25237 27656
rect 25188 27616 25194 27628
rect 25225 27625 25237 27628
rect 25271 27625 25283 27659
rect 25225 27619 25283 27625
rect 25958 27616 25964 27668
rect 26016 27616 26022 27668
rect 27801 27659 27859 27665
rect 27801 27625 27813 27659
rect 27847 27656 27859 27659
rect 28074 27656 28080 27668
rect 27847 27628 28080 27656
rect 27847 27625 27859 27628
rect 27801 27619 27859 27625
rect 27890 27588 27896 27600
rect 27724 27560 27896 27588
rect 25133 27523 25191 27529
rect 25133 27489 25145 27523
rect 25179 27520 25191 27523
rect 27621 27523 27679 27529
rect 25179 27492 25636 27520
rect 25179 27489 25191 27492
rect 25133 27483 25191 27489
rect 24213 27455 24271 27461
rect 24213 27421 24225 27455
rect 24259 27421 24271 27455
rect 24213 27415 24271 27421
rect 24673 27455 24731 27461
rect 24673 27421 24685 27455
rect 24719 27421 24731 27455
rect 24673 27415 24731 27421
rect 24118 27344 24124 27396
rect 24176 27344 24182 27396
rect 24228 27384 24256 27415
rect 24397 27387 24455 27393
rect 24397 27384 24409 27387
rect 24228 27356 24409 27384
rect 24397 27353 24409 27356
rect 24443 27353 24455 27387
rect 24397 27347 24455 27353
rect 24688 27316 24716 27415
rect 25314 27412 25320 27464
rect 25372 27452 25378 27464
rect 25409 27455 25467 27461
rect 25409 27452 25421 27455
rect 25372 27424 25421 27452
rect 25372 27412 25378 27424
rect 25409 27421 25421 27424
rect 25455 27421 25467 27455
rect 25409 27415 25467 27421
rect 25498 27412 25504 27464
rect 25556 27412 25562 27464
rect 25608 27461 25636 27492
rect 26344 27492 27016 27520
rect 25593 27455 25651 27461
rect 25593 27421 25605 27455
rect 25639 27421 25651 27455
rect 25593 27415 25651 27421
rect 25774 27412 25780 27464
rect 25832 27412 25838 27464
rect 26344 27461 26372 27492
rect 26988 27464 27016 27492
rect 27621 27489 27633 27523
rect 27667 27520 27679 27523
rect 27724 27520 27752 27560
rect 27890 27548 27896 27560
rect 27948 27548 27954 27600
rect 27667 27492 27752 27520
rect 27667 27489 27679 27492
rect 27621 27483 27679 27489
rect 26237 27455 26295 27461
rect 26237 27421 26249 27455
rect 26283 27421 26295 27455
rect 26237 27415 26295 27421
rect 26329 27455 26387 27461
rect 26329 27421 26341 27455
rect 26375 27421 26387 27455
rect 26329 27415 26387 27421
rect 26421 27455 26479 27461
rect 26421 27421 26433 27455
rect 26467 27421 26479 27455
rect 26421 27415 26479 27421
rect 26605 27455 26663 27461
rect 26605 27421 26617 27455
rect 26651 27452 26663 27455
rect 26878 27452 26884 27464
rect 26651 27424 26884 27452
rect 26651 27421 26663 27424
rect 26605 27415 26663 27421
rect 24762 27344 24768 27396
rect 24820 27344 24826 27396
rect 24946 27344 24952 27396
rect 25004 27344 25010 27396
rect 25516 27384 25544 27412
rect 26252 27384 26280 27415
rect 25516 27356 26280 27384
rect 26436 27384 26464 27415
rect 26878 27412 26884 27424
rect 26936 27412 26942 27464
rect 26970 27412 26976 27464
rect 27028 27412 27034 27464
rect 27249 27455 27307 27461
rect 27249 27421 27261 27455
rect 27295 27421 27307 27455
rect 27249 27415 27307 27421
rect 27065 27387 27123 27393
rect 27065 27384 27077 27387
rect 26436 27356 27077 27384
rect 27065 27353 27077 27356
rect 27111 27353 27123 27387
rect 27264 27384 27292 27415
rect 27430 27412 27436 27464
rect 27488 27412 27494 27464
rect 27525 27455 27583 27461
rect 27525 27421 27537 27455
rect 27571 27452 27583 27455
rect 27571 27424 27844 27452
rect 27571 27421 27583 27424
rect 27525 27415 27583 27421
rect 27617 27387 27675 27393
rect 27617 27384 27629 27387
rect 27264 27356 27629 27384
rect 27065 27347 27123 27353
rect 27617 27353 27629 27356
rect 27663 27353 27675 27387
rect 27617 27347 27675 27353
rect 27706 27344 27712 27396
rect 27764 27344 27770 27396
rect 27816 27384 27844 27424
rect 27890 27412 27896 27464
rect 27948 27412 27954 27464
rect 28000 27384 28028 27628
rect 28074 27616 28080 27628
rect 28132 27616 28138 27668
rect 32398 27616 32404 27668
rect 32456 27616 32462 27668
rect 28994 27548 29000 27600
rect 29052 27588 29058 27600
rect 29549 27591 29607 27597
rect 29549 27588 29561 27591
rect 29052 27560 29561 27588
rect 29052 27548 29058 27560
rect 29549 27557 29561 27560
rect 29595 27557 29607 27591
rect 29549 27551 29607 27557
rect 29012 27520 29040 27548
rect 29012 27492 29132 27520
rect 28258 27412 28264 27464
rect 28316 27452 28322 27464
rect 28718 27452 28724 27464
rect 28316 27424 28724 27452
rect 28316 27412 28322 27424
rect 28718 27412 28724 27424
rect 28776 27412 28782 27464
rect 28902 27412 28908 27464
rect 28960 27412 28966 27464
rect 29104 27461 29132 27492
rect 28997 27455 29055 27461
rect 28997 27421 29009 27455
rect 29043 27421 29055 27455
rect 28997 27415 29055 27421
rect 29089 27455 29147 27461
rect 29089 27421 29101 27455
rect 29135 27421 29147 27455
rect 29089 27415 29147 27421
rect 30929 27455 30987 27461
rect 30929 27421 30941 27455
rect 30975 27421 30987 27455
rect 30929 27415 30987 27421
rect 27816 27356 28028 27384
rect 28353 27387 28411 27393
rect 28353 27353 28365 27387
rect 28399 27384 28411 27387
rect 28810 27384 28816 27396
rect 28399 27356 28816 27384
rect 28399 27353 28411 27356
rect 28353 27347 28411 27353
rect 28810 27344 28816 27356
rect 28868 27344 28874 27396
rect 29012 27384 29040 27415
rect 29365 27387 29423 27393
rect 29012 27356 29132 27384
rect 23952 27288 24716 27316
rect 27724 27316 27752 27344
rect 29104 27328 29132 27356
rect 29365 27353 29377 27387
rect 29411 27384 29423 27387
rect 30662 27387 30720 27393
rect 30662 27384 30674 27387
rect 29411 27356 30674 27384
rect 29411 27353 29423 27356
rect 29365 27347 29423 27353
rect 30662 27353 30674 27356
rect 30708 27353 30720 27387
rect 30944 27384 30972 27415
rect 31018 27412 31024 27464
rect 31076 27412 31082 27464
rect 31294 27461 31300 27464
rect 31288 27452 31300 27461
rect 31255 27424 31300 27452
rect 31288 27415 31300 27424
rect 31294 27412 31300 27415
rect 31352 27412 31358 27464
rect 30944 27356 31524 27384
rect 30662 27347 30720 27353
rect 31496 27328 31524 27356
rect 28077 27319 28135 27325
rect 28077 27316 28089 27319
rect 27724 27288 28089 27316
rect 28077 27285 28089 27288
rect 28123 27285 28135 27319
rect 28077 27279 28135 27285
rect 29086 27276 29092 27328
rect 29144 27276 29150 27328
rect 31478 27276 31484 27328
rect 31536 27276 31542 27328
rect 1104 27226 35027 27248
rect 1104 27174 9390 27226
rect 9442 27174 9454 27226
rect 9506 27174 9518 27226
rect 9570 27174 9582 27226
rect 9634 27174 9646 27226
rect 9698 27174 17831 27226
rect 17883 27174 17895 27226
rect 17947 27174 17959 27226
rect 18011 27174 18023 27226
rect 18075 27174 18087 27226
rect 18139 27174 26272 27226
rect 26324 27174 26336 27226
rect 26388 27174 26400 27226
rect 26452 27174 26464 27226
rect 26516 27174 26528 27226
rect 26580 27174 34713 27226
rect 34765 27174 34777 27226
rect 34829 27174 34841 27226
rect 34893 27174 34905 27226
rect 34957 27174 34969 27226
rect 35021 27174 35027 27226
rect 1104 27152 35027 27174
rect 16850 27072 16856 27124
rect 16908 27112 16914 27124
rect 17129 27115 17187 27121
rect 17129 27112 17141 27115
rect 16908 27084 17141 27112
rect 16908 27072 16914 27084
rect 17129 27081 17141 27084
rect 17175 27081 17187 27115
rect 17129 27075 17187 27081
rect 18230 27072 18236 27124
rect 18288 27072 18294 27124
rect 18325 27115 18383 27121
rect 18325 27081 18337 27115
rect 18371 27112 18383 27115
rect 19334 27112 19340 27124
rect 18371 27084 19340 27112
rect 18371 27081 18383 27084
rect 18325 27075 18383 27081
rect 19334 27072 19340 27084
rect 19392 27072 19398 27124
rect 20717 27115 20775 27121
rect 19904 27084 20576 27112
rect 17957 27047 18015 27053
rect 17957 27013 17969 27047
rect 18003 27044 18015 27047
rect 18966 27044 18972 27056
rect 18003 27016 18972 27044
rect 18003 27013 18015 27016
rect 17957 27007 18015 27013
rect 18966 27004 18972 27016
rect 19024 27004 19030 27056
rect 17129 26979 17187 26985
rect 17129 26945 17141 26979
rect 17175 26976 17187 26979
rect 17310 26976 17316 26988
rect 17175 26948 17316 26976
rect 17175 26945 17187 26948
rect 17129 26939 17187 26945
rect 17310 26936 17316 26948
rect 17368 26936 17374 26988
rect 17589 26979 17647 26985
rect 17589 26945 17601 26979
rect 17635 26945 17647 26979
rect 17589 26939 17647 26945
rect 16853 26911 16911 26917
rect 16853 26877 16865 26911
rect 16899 26877 16911 26911
rect 17604 26908 17632 26939
rect 17678 26936 17684 26988
rect 17736 26936 17742 26988
rect 17862 26936 17868 26988
rect 17920 26936 17926 26988
rect 18095 26979 18153 26985
rect 18095 26945 18107 26979
rect 18141 26976 18153 26979
rect 18414 26976 18420 26988
rect 18141 26948 18420 26976
rect 18141 26945 18153 26948
rect 18095 26939 18153 26945
rect 18414 26936 18420 26948
rect 18472 26936 18478 26988
rect 19352 26976 19380 27072
rect 19426 27004 19432 27056
rect 19484 27053 19490 27056
rect 19484 27044 19496 27053
rect 19484 27016 19529 27044
rect 19484 27007 19496 27016
rect 19484 27004 19490 27007
rect 19797 26979 19855 26985
rect 19797 26976 19809 26979
rect 19352 26948 19809 26976
rect 19797 26945 19809 26948
rect 19843 26945 19855 26979
rect 19797 26939 19855 26945
rect 18230 26908 18236 26920
rect 17604 26880 18236 26908
rect 16853 26871 16911 26877
rect 16868 26772 16896 26871
rect 18230 26868 18236 26880
rect 18288 26868 18294 26920
rect 19702 26868 19708 26920
rect 19760 26908 19766 26920
rect 19904 26908 19932 27084
rect 20073 27047 20131 27053
rect 20073 27013 20085 27047
rect 20119 27044 20131 27047
rect 20119 27016 20300 27044
rect 20119 27013 20131 27016
rect 20073 27007 20131 27013
rect 20272 26985 20300 27016
rect 20346 27004 20352 27056
rect 20404 27004 20410 27056
rect 20548 27044 20576 27084
rect 20717 27081 20729 27115
rect 20763 27112 20775 27115
rect 20898 27112 20904 27124
rect 20763 27084 20904 27112
rect 20763 27081 20775 27084
rect 20717 27075 20775 27081
rect 20898 27072 20904 27084
rect 20956 27072 20962 27124
rect 21082 27072 21088 27124
rect 21140 27072 21146 27124
rect 21266 27072 21272 27124
rect 21324 27112 21330 27124
rect 23385 27115 23443 27121
rect 23385 27112 23397 27115
rect 21324 27084 23152 27112
rect 21324 27072 21330 27084
rect 20548 27016 21496 27044
rect 20257 26979 20315 26985
rect 20257 26945 20269 26979
rect 20303 26945 20315 26979
rect 20257 26939 20315 26945
rect 19760 26880 19932 26908
rect 19760 26868 19766 26880
rect 20070 26868 20076 26920
rect 20128 26868 20134 26920
rect 20364 26917 20392 27004
rect 20530 26936 20536 26988
rect 20588 26976 20594 26988
rect 20809 26979 20867 26985
rect 20809 26976 20821 26979
rect 20588 26948 20821 26976
rect 20588 26936 20594 26948
rect 20809 26945 20821 26948
rect 20855 26945 20867 26979
rect 21174 26976 21180 26988
rect 20809 26939 20867 26945
rect 20916 26948 21180 26976
rect 20349 26911 20407 26917
rect 20349 26877 20361 26911
rect 20395 26877 20407 26911
rect 20349 26871 20407 26877
rect 20441 26911 20499 26917
rect 20441 26877 20453 26911
rect 20487 26908 20499 26911
rect 20714 26908 20720 26920
rect 20487 26880 20720 26908
rect 20487 26877 20499 26880
rect 20441 26871 20499 26877
rect 20714 26868 20720 26880
rect 20772 26868 20778 26920
rect 17037 26843 17095 26849
rect 17037 26809 17049 26843
rect 17083 26840 17095 26843
rect 17494 26840 17500 26852
rect 17083 26812 17500 26840
rect 17083 26809 17095 26812
rect 17037 26803 17095 26809
rect 17494 26800 17500 26812
rect 17552 26800 17558 26852
rect 20916 26840 20944 26948
rect 21174 26936 21180 26948
rect 21232 26936 21238 26988
rect 21358 26936 21364 26988
rect 21416 26936 21422 26988
rect 21468 26976 21496 27016
rect 21468 26948 22094 26976
rect 21085 26911 21143 26917
rect 21085 26877 21097 26911
rect 21131 26908 21143 26911
rect 21266 26908 21272 26920
rect 21131 26880 21272 26908
rect 21131 26877 21143 26880
rect 21085 26871 21143 26877
rect 21266 26868 21272 26880
rect 21324 26868 21330 26920
rect 19904 26812 20944 26840
rect 16942 26772 16948 26784
rect 16868 26744 16948 26772
rect 16942 26732 16948 26744
rect 17000 26772 17006 26784
rect 18506 26772 18512 26784
rect 17000 26744 18512 26772
rect 17000 26732 17006 26744
rect 18506 26732 18512 26744
rect 18564 26732 18570 26784
rect 19426 26732 19432 26784
rect 19484 26772 19490 26784
rect 19904 26781 19932 26812
rect 19889 26775 19947 26781
rect 19889 26772 19901 26775
rect 19484 26744 19901 26772
rect 19484 26732 19490 26744
rect 19889 26741 19901 26744
rect 19935 26741 19947 26775
rect 19889 26735 19947 26741
rect 20714 26732 20720 26784
rect 20772 26772 20778 26784
rect 20901 26775 20959 26781
rect 20901 26772 20913 26775
rect 20772 26744 20913 26772
rect 20772 26732 20778 26744
rect 20901 26741 20913 26744
rect 20947 26772 20959 26775
rect 21082 26772 21088 26784
rect 20947 26744 21088 26772
rect 20947 26741 20959 26744
rect 20901 26735 20959 26741
rect 21082 26732 21088 26744
rect 21140 26732 21146 26784
rect 21174 26732 21180 26784
rect 21232 26772 21238 26784
rect 21726 26772 21732 26784
rect 21232 26744 21732 26772
rect 21232 26732 21238 26744
rect 21726 26732 21732 26744
rect 21784 26772 21790 26784
rect 21821 26775 21879 26781
rect 21821 26772 21833 26775
rect 21784 26744 21833 26772
rect 21784 26732 21790 26744
rect 21821 26741 21833 26744
rect 21867 26741 21879 26775
rect 22066 26772 22094 26948
rect 22462 26936 22468 26988
rect 22520 26976 22526 26988
rect 22934 26979 22992 26985
rect 22934 26976 22946 26979
rect 22520 26948 22946 26976
rect 22520 26936 22526 26948
rect 22934 26945 22946 26948
rect 22980 26945 22992 26979
rect 22934 26939 22992 26945
rect 23124 26908 23152 27084
rect 23216 27084 23397 27112
rect 23216 26988 23244 27084
rect 23385 27081 23397 27084
rect 23431 27081 23443 27115
rect 23385 27075 23443 27081
rect 23566 27072 23572 27124
rect 23624 27112 23630 27124
rect 23661 27115 23719 27121
rect 23661 27112 23673 27115
rect 23624 27084 23673 27112
rect 23624 27072 23630 27084
rect 23661 27081 23673 27084
rect 23707 27081 23719 27115
rect 23661 27075 23719 27081
rect 24762 27072 24768 27124
rect 24820 27112 24826 27124
rect 24949 27115 25007 27121
rect 24949 27112 24961 27115
rect 24820 27084 24961 27112
rect 24820 27072 24826 27084
rect 24949 27081 24961 27084
rect 24995 27081 25007 27115
rect 24949 27075 25007 27081
rect 23198 26936 23204 26988
rect 23256 26936 23262 26988
rect 23584 26985 23612 27072
rect 24118 27044 24124 27056
rect 23768 27016 24124 27044
rect 23569 26979 23627 26985
rect 23569 26945 23581 26979
rect 23615 26945 23627 26979
rect 23569 26939 23627 26945
rect 23768 26908 23796 27016
rect 24118 27004 24124 27016
rect 24176 27044 24182 27056
rect 24486 27044 24492 27056
rect 24176 27016 24492 27044
rect 24176 27004 24182 27016
rect 24486 27004 24492 27016
rect 24544 27004 24550 27056
rect 24964 27044 24992 27075
rect 25774 27072 25780 27124
rect 25832 27112 25838 27124
rect 25869 27115 25927 27121
rect 25869 27112 25881 27115
rect 25832 27084 25881 27112
rect 25832 27072 25838 27084
rect 25869 27081 25881 27084
rect 25915 27081 25927 27115
rect 25869 27075 25927 27081
rect 28902 27072 28908 27124
rect 28960 27072 28966 27124
rect 29089 27115 29147 27121
rect 29089 27081 29101 27115
rect 29135 27112 29147 27115
rect 29178 27112 29184 27124
rect 29135 27084 29184 27112
rect 29135 27081 29147 27084
rect 29089 27075 29147 27081
rect 29178 27072 29184 27084
rect 29236 27072 29242 27124
rect 29362 27072 29368 27124
rect 29420 27072 29426 27124
rect 31110 27072 31116 27124
rect 31168 27112 31174 27124
rect 31205 27115 31263 27121
rect 31205 27112 31217 27115
rect 31168 27084 31217 27112
rect 31168 27072 31174 27084
rect 31205 27081 31217 27084
rect 31251 27081 31263 27115
rect 32398 27112 32404 27124
rect 31205 27075 31263 27081
rect 31726 27084 32404 27112
rect 28920 27044 28948 27072
rect 29273 27047 29331 27053
rect 29273 27044 29285 27047
rect 24964 27016 25728 27044
rect 28920 27016 29285 27044
rect 23845 26979 23903 26985
rect 23845 26945 23857 26979
rect 23891 26945 23903 26979
rect 23845 26939 23903 26945
rect 23124 26880 23796 26908
rect 23198 26800 23204 26852
rect 23256 26800 23262 26852
rect 23860 26840 23888 26939
rect 24762 26936 24768 26988
rect 24820 26976 24826 26988
rect 24857 26979 24915 26985
rect 24857 26976 24869 26979
rect 24820 26948 24869 26976
rect 24820 26936 24826 26948
rect 24857 26945 24869 26948
rect 24903 26945 24915 26979
rect 24857 26939 24915 26945
rect 24946 26936 24952 26988
rect 25004 26936 25010 26988
rect 25314 26936 25320 26988
rect 25372 26936 25378 26988
rect 25498 26936 25504 26988
rect 25556 26936 25562 26988
rect 25700 26985 25728 27016
rect 29273 27013 29285 27016
rect 29319 27013 29331 27047
rect 29273 27007 29331 27013
rect 25593 26979 25651 26985
rect 25593 26945 25605 26979
rect 25639 26945 25651 26979
rect 25593 26939 25651 26945
rect 25685 26979 25743 26985
rect 25685 26945 25697 26979
rect 25731 26945 25743 26979
rect 25685 26939 25743 26945
rect 28721 26979 28779 26985
rect 28721 26945 28733 26979
rect 28767 26976 28779 26979
rect 28810 26976 28816 26988
rect 28767 26948 28816 26976
rect 28767 26945 28779 26948
rect 28721 26939 28779 26945
rect 24964 26908 24992 26936
rect 25608 26908 25636 26939
rect 28810 26936 28816 26948
rect 28868 26936 28874 26988
rect 28905 26979 28963 26985
rect 28905 26945 28917 26979
rect 28951 26976 28963 26979
rect 28994 26976 29000 26988
rect 28951 26948 29000 26976
rect 28951 26945 28963 26948
rect 28905 26939 28963 26945
rect 27338 26908 27344 26920
rect 24964 26880 27344 26908
rect 27338 26868 27344 26880
rect 27396 26908 27402 26920
rect 28920 26908 28948 26939
rect 28994 26936 29000 26948
rect 29052 26936 29058 26988
rect 29380 26985 29408 27072
rect 31726 27044 31754 27084
rect 32398 27072 32404 27084
rect 32456 27072 32462 27124
rect 31680 27016 31754 27044
rect 29181 26979 29239 26985
rect 29181 26945 29193 26979
rect 29227 26945 29239 26979
rect 29181 26939 29239 26945
rect 29365 26979 29423 26985
rect 29365 26945 29377 26979
rect 29411 26945 29423 26979
rect 29365 26939 29423 26945
rect 27396 26880 28948 26908
rect 27396 26868 27402 26880
rect 29086 26868 29092 26920
rect 29144 26908 29150 26920
rect 29196 26908 29224 26939
rect 30926 26936 30932 26988
rect 30984 26936 30990 26988
rect 31021 26979 31079 26985
rect 31021 26945 31033 26979
rect 31067 26976 31079 26979
rect 31202 26976 31208 26988
rect 31067 26948 31208 26976
rect 31067 26945 31079 26948
rect 31021 26939 31079 26945
rect 31202 26936 31208 26948
rect 31260 26936 31266 26988
rect 31680 26985 31708 27016
rect 31665 26979 31723 26985
rect 31665 26945 31677 26979
rect 31711 26945 31723 26979
rect 31665 26939 31723 26945
rect 31757 26979 31815 26985
rect 31757 26945 31769 26979
rect 31803 26945 31815 26979
rect 31757 26939 31815 26945
rect 31941 26979 31999 26985
rect 31941 26945 31953 26979
rect 31987 26976 31999 26979
rect 32493 26979 32551 26985
rect 32493 26976 32505 26979
rect 31987 26948 32505 26976
rect 31987 26945 31999 26948
rect 31941 26939 31999 26945
rect 32493 26945 32505 26948
rect 32539 26945 32551 26979
rect 32493 26939 32551 26945
rect 29144 26880 29224 26908
rect 31220 26908 31248 26936
rect 31772 26908 31800 26939
rect 31220 26880 31800 26908
rect 29144 26868 29150 26880
rect 33042 26840 33048 26852
rect 23860 26812 33048 26840
rect 33042 26800 33048 26812
rect 33100 26800 33106 26852
rect 22830 26772 22836 26784
rect 22066 26744 22836 26772
rect 21821 26735 21879 26741
rect 22830 26732 22836 26744
rect 22888 26772 22894 26784
rect 23216 26772 23244 26800
rect 22888 26744 23244 26772
rect 22888 26732 22894 26744
rect 32214 26732 32220 26784
rect 32272 26772 32278 26784
rect 32309 26775 32367 26781
rect 32309 26772 32321 26775
rect 32272 26744 32321 26772
rect 32272 26732 32278 26744
rect 32309 26741 32321 26744
rect 32355 26741 32367 26775
rect 32309 26735 32367 26741
rect 1104 26682 34868 26704
rect 1104 26630 5170 26682
rect 5222 26630 5234 26682
rect 5286 26630 5298 26682
rect 5350 26630 5362 26682
rect 5414 26630 5426 26682
rect 5478 26630 13611 26682
rect 13663 26630 13675 26682
rect 13727 26630 13739 26682
rect 13791 26630 13803 26682
rect 13855 26630 13867 26682
rect 13919 26630 22052 26682
rect 22104 26630 22116 26682
rect 22168 26630 22180 26682
rect 22232 26630 22244 26682
rect 22296 26630 22308 26682
rect 22360 26630 30493 26682
rect 30545 26630 30557 26682
rect 30609 26630 30621 26682
rect 30673 26630 30685 26682
rect 30737 26630 30749 26682
rect 30801 26630 34868 26682
rect 1104 26608 34868 26630
rect 17678 26528 17684 26580
rect 17736 26568 17742 26580
rect 17862 26568 17868 26580
rect 17736 26540 17868 26568
rect 17736 26528 17742 26540
rect 17862 26528 17868 26540
rect 17920 26528 17926 26580
rect 18506 26528 18512 26580
rect 18564 26568 18570 26580
rect 19702 26568 19708 26580
rect 18564 26540 19708 26568
rect 18564 26528 18570 26540
rect 19702 26528 19708 26540
rect 19760 26528 19766 26580
rect 20070 26528 20076 26580
rect 20128 26568 20134 26580
rect 20165 26571 20223 26577
rect 20165 26568 20177 26571
rect 20128 26540 20177 26568
rect 20128 26528 20134 26540
rect 20165 26537 20177 26540
rect 20211 26537 20223 26571
rect 20165 26531 20223 26537
rect 20898 26528 20904 26580
rect 20956 26528 20962 26580
rect 21177 26571 21235 26577
rect 21177 26568 21189 26571
rect 21100 26540 21189 26568
rect 21100 26512 21128 26540
rect 21177 26537 21189 26540
rect 21223 26537 21235 26571
rect 21177 26531 21235 26537
rect 22005 26571 22063 26577
rect 22005 26537 22017 26571
rect 22051 26568 22063 26571
rect 22462 26568 22468 26580
rect 22051 26540 22468 26568
rect 22051 26537 22063 26540
rect 22005 26531 22063 26537
rect 22462 26528 22468 26540
rect 22520 26528 22526 26580
rect 23750 26568 23756 26580
rect 22664 26540 23756 26568
rect 18874 26460 18880 26512
rect 18932 26500 18938 26512
rect 20806 26500 20812 26512
rect 18932 26472 20812 26500
rect 18932 26460 18938 26472
rect 20806 26460 20812 26472
rect 20864 26460 20870 26512
rect 21082 26460 21088 26512
rect 21140 26460 21146 26512
rect 21652 26472 21864 26500
rect 20714 26392 20720 26444
rect 20772 26392 20778 26444
rect 21652 26432 21680 26472
rect 21560 26404 21680 26432
rect 21836 26432 21864 26472
rect 21910 26460 21916 26512
rect 21968 26500 21974 26512
rect 22664 26509 22692 26540
rect 23750 26528 23756 26540
rect 23808 26568 23814 26580
rect 24397 26571 24455 26577
rect 24397 26568 24409 26571
rect 23808 26540 24409 26568
rect 23808 26528 23814 26540
rect 24397 26537 24409 26540
rect 24443 26537 24455 26571
rect 24397 26531 24455 26537
rect 24578 26528 24584 26580
rect 24636 26528 24642 26580
rect 25225 26571 25283 26577
rect 25225 26537 25237 26571
rect 25271 26568 25283 26571
rect 25314 26568 25320 26580
rect 25271 26540 25320 26568
rect 25271 26537 25283 26540
rect 25225 26531 25283 26537
rect 25314 26528 25320 26540
rect 25372 26528 25378 26580
rect 25498 26528 25504 26580
rect 25556 26568 25562 26580
rect 25869 26571 25927 26577
rect 25869 26568 25881 26571
rect 25556 26540 25881 26568
rect 25556 26528 25562 26540
rect 25869 26537 25881 26540
rect 25915 26537 25927 26571
rect 25869 26531 25927 26537
rect 26970 26528 26976 26580
rect 27028 26568 27034 26580
rect 27430 26568 27436 26580
rect 27028 26540 27436 26568
rect 27028 26528 27034 26540
rect 27430 26528 27436 26540
rect 27488 26568 27494 26580
rect 28997 26571 29055 26577
rect 28997 26568 29009 26571
rect 27488 26540 29009 26568
rect 27488 26528 27494 26540
rect 28997 26537 29009 26540
rect 29043 26568 29055 26571
rect 29086 26568 29092 26580
rect 29043 26540 29092 26568
rect 29043 26537 29055 26540
rect 28997 26531 29055 26537
rect 29086 26528 29092 26540
rect 29144 26528 29150 26580
rect 22649 26503 22707 26509
rect 21968 26472 22324 26500
rect 21968 26460 21974 26472
rect 22189 26435 22247 26441
rect 22189 26432 22201 26435
rect 21836 26404 22201 26432
rect 16301 26367 16359 26373
rect 16301 26333 16313 26367
rect 16347 26333 16359 26367
rect 16301 26327 16359 26333
rect 16568 26367 16626 26373
rect 16568 26333 16580 26367
rect 16614 26364 16626 26367
rect 16850 26364 16856 26376
rect 16614 26336 16856 26364
rect 16614 26333 16626 26336
rect 16568 26327 16626 26333
rect 16316 26296 16344 26327
rect 16850 26324 16856 26336
rect 16908 26324 16914 26376
rect 17586 26324 17592 26376
rect 17644 26364 17650 26376
rect 19337 26367 19395 26373
rect 19337 26364 19349 26367
rect 17644 26336 19349 26364
rect 17644 26324 17650 26336
rect 19337 26333 19349 26336
rect 19383 26333 19395 26367
rect 19337 26327 19395 26333
rect 19426 26324 19432 26376
rect 19484 26324 19490 26376
rect 20530 26324 20536 26376
rect 20588 26364 20594 26376
rect 20625 26367 20683 26373
rect 20625 26364 20637 26367
rect 20588 26336 20637 26364
rect 20588 26324 20594 26336
rect 20625 26333 20637 26336
rect 20671 26333 20683 26367
rect 20625 26327 20683 26333
rect 20898 26324 20904 26376
rect 20956 26364 20962 26376
rect 21077 26369 21135 26375
rect 21077 26366 21089 26369
rect 21008 26364 21089 26366
rect 20956 26338 21089 26364
rect 20956 26336 21036 26338
rect 20956 26324 20962 26336
rect 21077 26335 21089 26338
rect 21123 26335 21135 26369
rect 21077 26329 21135 26335
rect 21266 26324 21272 26376
rect 21324 26324 21330 26376
rect 21358 26324 21364 26376
rect 21416 26324 21422 26376
rect 21560 26373 21588 26404
rect 22189 26401 22201 26404
rect 22235 26401 22247 26435
rect 22189 26395 22247 26401
rect 21545 26367 21603 26373
rect 21545 26333 21557 26367
rect 21591 26333 21603 26367
rect 21545 26327 21603 26333
rect 21637 26367 21695 26373
rect 21637 26333 21649 26367
rect 21683 26333 21695 26367
rect 21637 26327 21695 26333
rect 16666 26296 16672 26308
rect 16316 26268 16672 26296
rect 16666 26256 16672 26268
rect 16724 26296 16730 26308
rect 18506 26296 18512 26308
rect 16724 26268 18512 26296
rect 16724 26256 16730 26268
rect 18506 26256 18512 26268
rect 18564 26256 18570 26308
rect 20254 26256 20260 26308
rect 20312 26256 20318 26308
rect 21652 26296 21680 26327
rect 21726 26324 21732 26376
rect 21784 26324 21790 26376
rect 22296 26373 22324 26472
rect 22649 26469 22661 26503
rect 22695 26469 22707 26503
rect 22649 26463 22707 26469
rect 22741 26503 22799 26509
rect 22741 26469 22753 26503
rect 22787 26469 22799 26503
rect 24605 26500 24633 26528
rect 24605 26472 26372 26500
rect 22741 26463 22799 26469
rect 22756 26432 22784 26463
rect 22756 26404 22968 26432
rect 22097 26367 22155 26373
rect 22097 26333 22109 26367
rect 22143 26333 22155 26367
rect 22097 26327 22155 26333
rect 22281 26367 22339 26373
rect 22281 26333 22293 26367
rect 22327 26333 22339 26367
rect 22281 26327 22339 26333
rect 22741 26367 22799 26373
rect 22741 26333 22753 26367
rect 22787 26333 22799 26367
rect 22741 26327 22799 26333
rect 21818 26296 21824 26308
rect 21652 26268 21824 26296
rect 21818 26256 21824 26268
rect 21876 26296 21882 26308
rect 22112 26296 22140 26327
rect 21876 26268 22140 26296
rect 21876 26256 21882 26268
rect 22462 26256 22468 26308
rect 22520 26256 22526 26308
rect 22756 26296 22784 26327
rect 22830 26324 22836 26376
rect 22888 26324 22894 26376
rect 22940 26364 22968 26404
rect 24964 26404 25636 26432
rect 23089 26367 23147 26373
rect 23089 26364 23101 26367
rect 22940 26336 23101 26364
rect 23089 26333 23101 26336
rect 23135 26333 23147 26367
rect 24857 26367 24915 26373
rect 24857 26364 24869 26367
rect 23089 26327 23147 26333
rect 23584 26336 24869 26364
rect 23474 26296 23480 26308
rect 22756 26268 23480 26296
rect 23474 26256 23480 26268
rect 23532 26256 23538 26308
rect 23584 26240 23612 26336
rect 24857 26333 24869 26336
rect 24903 26333 24915 26367
rect 24857 26327 24915 26333
rect 24762 26296 24768 26308
rect 24228 26268 24768 26296
rect 24228 26240 24256 26268
rect 24762 26256 24768 26268
rect 24820 26256 24826 26308
rect 17402 26188 17408 26240
rect 17460 26228 17466 26240
rect 21266 26228 21272 26240
rect 17460 26200 21272 26228
rect 17460 26188 17466 26200
rect 21266 26188 21272 26200
rect 21324 26188 21330 26240
rect 23566 26188 23572 26240
rect 23624 26188 23630 26240
rect 24210 26188 24216 26240
rect 24268 26188 24274 26240
rect 24565 26231 24623 26237
rect 24565 26197 24577 26231
rect 24611 26228 24623 26231
rect 24872 26228 24900 26327
rect 24964 26240 24992 26404
rect 25608 26373 25636 26404
rect 25409 26367 25467 26373
rect 25409 26333 25421 26367
rect 25455 26333 25467 26367
rect 25409 26327 25467 26333
rect 25593 26367 25651 26373
rect 25593 26333 25605 26367
rect 25639 26333 25651 26367
rect 25593 26327 25651 26333
rect 25777 26367 25835 26373
rect 25777 26333 25789 26367
rect 25823 26364 25835 26367
rect 26142 26364 26148 26376
rect 25823 26336 26148 26364
rect 25823 26333 25835 26336
rect 25777 26327 25835 26333
rect 24611 26200 24900 26228
rect 24611 26197 24623 26200
rect 24565 26191 24623 26197
rect 24946 26188 24952 26240
rect 25004 26188 25010 26240
rect 25424 26228 25452 26327
rect 26142 26324 26148 26336
rect 26200 26324 26206 26376
rect 26234 26324 26240 26376
rect 26292 26324 26298 26376
rect 26344 26373 26372 26472
rect 26878 26460 26884 26512
rect 26936 26500 26942 26512
rect 28718 26500 28724 26512
rect 26936 26472 28724 26500
rect 26936 26460 26942 26472
rect 27172 26373 27200 26472
rect 28718 26460 28724 26472
rect 28776 26460 28782 26512
rect 29546 26460 29552 26512
rect 29604 26500 29610 26512
rect 29825 26503 29883 26509
rect 29825 26500 29837 26503
rect 29604 26472 29837 26500
rect 29604 26460 29610 26472
rect 29825 26469 29837 26472
rect 29871 26469 29883 26503
rect 29825 26463 29883 26469
rect 32950 26460 32956 26512
rect 33008 26500 33014 26512
rect 33321 26503 33379 26509
rect 33321 26500 33333 26503
rect 33008 26472 33333 26500
rect 33008 26460 33014 26472
rect 33321 26469 33333 26472
rect 33367 26469 33379 26503
rect 33321 26463 33379 26469
rect 27246 26392 27252 26444
rect 27304 26432 27310 26444
rect 27798 26432 27804 26444
rect 27304 26404 27804 26432
rect 27304 26392 27310 26404
rect 27798 26392 27804 26404
rect 27856 26432 27862 26444
rect 30834 26432 30840 26444
rect 27856 26404 28856 26432
rect 27856 26392 27862 26404
rect 28828 26376 28856 26404
rect 29564 26404 30840 26432
rect 26329 26367 26387 26373
rect 26329 26333 26341 26367
rect 26375 26333 26387 26367
rect 26329 26327 26387 26333
rect 27157 26367 27215 26373
rect 27157 26333 27169 26367
rect 27203 26333 27215 26367
rect 27157 26327 27215 26333
rect 27338 26324 27344 26376
rect 27396 26324 27402 26376
rect 27430 26324 27436 26376
rect 27488 26324 27494 26376
rect 27525 26367 27583 26373
rect 27525 26333 27537 26367
rect 27571 26364 27583 26367
rect 28077 26367 28135 26373
rect 28077 26364 28089 26367
rect 27571 26336 28089 26364
rect 27571 26333 27583 26336
rect 27525 26327 27583 26333
rect 28077 26333 28089 26336
rect 28123 26364 28135 26367
rect 28626 26364 28632 26376
rect 28123 26336 28632 26364
rect 28123 26333 28135 26336
rect 28077 26327 28135 26333
rect 25501 26299 25559 26305
rect 25501 26265 25513 26299
rect 25547 26296 25559 26299
rect 26053 26299 26111 26305
rect 26053 26296 26065 26299
rect 25547 26268 26065 26296
rect 25547 26265 25559 26268
rect 25501 26259 25559 26265
rect 26053 26265 26065 26268
rect 26099 26296 26111 26299
rect 27540 26296 27568 26327
rect 28626 26324 28632 26336
rect 28684 26324 28690 26376
rect 28810 26324 28816 26376
rect 28868 26324 28874 26376
rect 29564 26373 29592 26404
rect 29840 26376 29868 26404
rect 30834 26392 30840 26404
rect 30892 26392 30898 26444
rect 29549 26367 29607 26373
rect 29549 26333 29561 26367
rect 29595 26333 29607 26367
rect 29549 26327 29607 26333
rect 29822 26324 29828 26376
rect 29880 26324 29886 26376
rect 31018 26324 31024 26376
rect 31076 26364 31082 26376
rect 31754 26364 31760 26376
rect 31076 26336 31760 26364
rect 31076 26324 31082 26336
rect 31754 26324 31760 26336
rect 31812 26364 31818 26376
rect 32214 26373 32220 26376
rect 31941 26367 31999 26373
rect 31941 26364 31953 26367
rect 31812 26336 31953 26364
rect 31812 26324 31818 26336
rect 31941 26333 31953 26336
rect 31987 26333 31999 26367
rect 32208 26364 32220 26373
rect 32175 26336 32220 26364
rect 31941 26327 31999 26333
rect 32208 26327 32220 26336
rect 32214 26324 32220 26327
rect 32272 26324 32278 26376
rect 27893 26299 27951 26305
rect 27893 26296 27905 26299
rect 26099 26268 27568 26296
rect 27724 26268 27905 26296
rect 26099 26265 26111 26268
rect 26053 26259 26111 26265
rect 27724 26240 27752 26268
rect 27893 26265 27905 26268
rect 27939 26265 27951 26299
rect 27893 26259 27951 26265
rect 28261 26299 28319 26305
rect 28261 26265 28273 26299
rect 28307 26296 28319 26299
rect 28902 26296 28908 26308
rect 28307 26268 28908 26296
rect 28307 26265 28319 26268
rect 28261 26259 28319 26265
rect 28902 26256 28908 26268
rect 28960 26256 28966 26308
rect 25682 26228 25688 26240
rect 25424 26200 25688 26228
rect 25682 26188 25688 26200
rect 25740 26228 25746 26240
rect 26234 26228 26240 26240
rect 25740 26200 26240 26228
rect 25740 26188 25746 26200
rect 26234 26188 26240 26200
rect 26292 26228 26298 26240
rect 26421 26231 26479 26237
rect 26421 26228 26433 26231
rect 26292 26200 26433 26228
rect 26292 26188 26298 26200
rect 26421 26197 26433 26200
rect 26467 26197 26479 26231
rect 26421 26191 26479 26197
rect 26694 26188 26700 26240
rect 26752 26228 26758 26240
rect 27706 26228 27712 26240
rect 26752 26200 27712 26228
rect 26752 26188 26758 26200
rect 27706 26188 27712 26200
rect 27764 26188 27770 26240
rect 27798 26188 27804 26240
rect 27856 26188 27862 26240
rect 30006 26188 30012 26240
rect 30064 26188 30070 26240
rect 1104 26138 35027 26160
rect 1104 26086 9390 26138
rect 9442 26086 9454 26138
rect 9506 26086 9518 26138
rect 9570 26086 9582 26138
rect 9634 26086 9646 26138
rect 9698 26086 17831 26138
rect 17883 26086 17895 26138
rect 17947 26086 17959 26138
rect 18011 26086 18023 26138
rect 18075 26086 18087 26138
rect 18139 26086 26272 26138
rect 26324 26086 26336 26138
rect 26388 26086 26400 26138
rect 26452 26086 26464 26138
rect 26516 26086 26528 26138
rect 26580 26086 34713 26138
rect 34765 26086 34777 26138
rect 34829 26086 34841 26138
rect 34893 26086 34905 26138
rect 34957 26086 34969 26138
rect 35021 26086 35027 26138
rect 1104 26064 35027 26086
rect 17494 25984 17500 26036
rect 17552 25984 17558 26036
rect 17665 26027 17723 26033
rect 17665 26024 17677 26027
rect 17604 25996 17677 26024
rect 17604 25956 17632 25996
rect 17665 25993 17677 25996
rect 17711 26024 17723 26027
rect 17711 25996 18828 26024
rect 17711 25993 17723 25996
rect 17665 25987 17723 25993
rect 17144 25928 17632 25956
rect 17144 25900 17172 25928
rect 17770 25916 17776 25968
rect 17828 25956 17834 25968
rect 17865 25959 17923 25965
rect 17865 25956 17877 25959
rect 17828 25928 17877 25956
rect 17828 25916 17834 25928
rect 17865 25925 17877 25928
rect 17911 25925 17923 25959
rect 17865 25919 17923 25925
rect 18340 25928 18736 25956
rect 17126 25848 17132 25900
rect 17184 25848 17190 25900
rect 17221 25891 17279 25897
rect 17221 25857 17233 25891
rect 17267 25857 17279 25891
rect 17221 25851 17279 25857
rect 17405 25891 17463 25897
rect 17405 25857 17417 25891
rect 17451 25888 17463 25891
rect 17788 25888 17816 25916
rect 17451 25860 17816 25888
rect 17451 25857 17463 25860
rect 17405 25851 17463 25857
rect 17236 25696 17264 25851
rect 17310 25780 17316 25832
rect 17368 25820 17374 25832
rect 17788 25820 17816 25860
rect 17954 25848 17960 25900
rect 18012 25888 18018 25900
rect 18340 25897 18368 25928
rect 18049 25891 18107 25897
rect 18049 25888 18061 25891
rect 18012 25860 18061 25888
rect 18012 25848 18018 25860
rect 18049 25857 18061 25860
rect 18095 25857 18107 25891
rect 18049 25851 18107 25857
rect 18325 25891 18383 25897
rect 18325 25857 18337 25891
rect 18371 25857 18383 25891
rect 18325 25851 18383 25857
rect 18417 25891 18475 25897
rect 18417 25857 18429 25891
rect 18463 25857 18475 25891
rect 18417 25851 18475 25857
rect 18141 25823 18199 25829
rect 18141 25820 18153 25823
rect 17368 25792 17448 25820
rect 17788 25792 18153 25820
rect 17368 25780 17374 25792
rect 17420 25761 17448 25792
rect 18141 25789 18153 25792
rect 18187 25789 18199 25823
rect 18141 25783 18199 25789
rect 18432 25764 18460 25851
rect 18708 25820 18736 25928
rect 18800 25894 18828 25996
rect 20898 25984 20904 26036
rect 20956 26024 20962 26036
rect 21085 26027 21143 26033
rect 21085 26024 21097 26027
rect 20956 25996 21097 26024
rect 20956 25984 20962 25996
rect 21085 25993 21097 25996
rect 21131 25993 21143 26027
rect 23753 26027 23811 26033
rect 21085 25987 21143 25993
rect 22066 25996 22968 26024
rect 19076 25928 19334 25956
rect 19076 25897 19104 25928
rect 18877 25894 18935 25897
rect 18800 25891 18935 25894
rect 18800 25866 18889 25891
rect 18877 25857 18889 25866
rect 18923 25857 18935 25891
rect 18877 25851 18935 25857
rect 19061 25891 19119 25897
rect 19061 25857 19073 25891
rect 19107 25857 19119 25891
rect 19061 25851 19119 25857
rect 19076 25820 19104 25851
rect 19150 25848 19156 25900
rect 19208 25848 19214 25900
rect 18708 25792 19104 25820
rect 19306 25820 19334 25928
rect 21174 25916 21180 25968
rect 21232 25956 21238 25968
rect 21269 25959 21327 25965
rect 21269 25956 21281 25959
rect 21232 25928 21281 25956
rect 21232 25916 21238 25928
rect 21269 25925 21281 25928
rect 21315 25925 21327 25959
rect 22066 25956 22094 25996
rect 22940 25956 22968 25996
rect 23753 25993 23765 26027
rect 23799 26024 23811 26027
rect 24121 26027 24179 26033
rect 24121 26024 24133 26027
rect 23799 25996 24133 26024
rect 23799 25993 23811 25996
rect 23753 25987 23811 25993
rect 24121 25993 24133 25996
rect 24167 26024 24179 26027
rect 24578 26024 24584 26036
rect 24167 25996 24584 26024
rect 24167 25993 24179 25996
rect 24121 25987 24179 25993
rect 24578 25984 24584 25996
rect 24636 25984 24642 26036
rect 25516 25996 25912 26024
rect 23937 25959 23995 25965
rect 21269 25919 21327 25925
rect 21376 25928 22094 25956
rect 22204 25928 22876 25956
rect 22940 25928 23888 25956
rect 19978 25848 19984 25900
rect 20036 25888 20042 25900
rect 21376 25888 21404 25928
rect 20036 25860 21404 25888
rect 20036 25848 20042 25860
rect 21450 25848 21456 25900
rect 21508 25848 21514 25900
rect 22204 25897 22232 25928
rect 22848 25900 22876 25928
rect 22189 25891 22247 25897
rect 22189 25857 22201 25891
rect 22235 25857 22247 25891
rect 22189 25851 22247 25857
rect 22456 25891 22514 25897
rect 22456 25857 22468 25891
rect 22502 25888 22514 25891
rect 22738 25888 22744 25900
rect 22502 25860 22744 25888
rect 22502 25857 22514 25860
rect 22456 25851 22514 25857
rect 22738 25848 22744 25860
rect 22796 25848 22802 25900
rect 22830 25848 22836 25900
rect 22888 25848 22894 25900
rect 23566 25848 23572 25900
rect 23624 25888 23630 25900
rect 23661 25891 23719 25897
rect 23661 25888 23673 25891
rect 23624 25860 23673 25888
rect 23624 25848 23630 25860
rect 23661 25857 23673 25860
rect 23707 25857 23719 25891
rect 23860 25888 23888 25928
rect 23937 25925 23949 25959
rect 23983 25956 23995 25959
rect 24210 25956 24216 25968
rect 23983 25928 24216 25956
rect 23983 25925 23995 25928
rect 23937 25919 23995 25925
rect 24210 25916 24216 25928
rect 24268 25916 24274 25968
rect 24302 25916 24308 25968
rect 24360 25956 24366 25968
rect 25038 25956 25044 25968
rect 24360 25928 25044 25956
rect 24360 25916 24366 25928
rect 25038 25916 25044 25928
rect 25096 25956 25102 25968
rect 25516 25956 25544 25996
rect 25884 25965 25912 25996
rect 26694 25984 26700 26036
rect 26752 25984 26758 26036
rect 27249 26027 27307 26033
rect 27249 25993 27261 26027
rect 27295 26024 27307 26027
rect 27338 26024 27344 26036
rect 27295 25996 27344 26024
rect 27295 25993 27307 25996
rect 27249 25987 27307 25993
rect 27338 25984 27344 25996
rect 27396 25984 27402 26036
rect 27614 25984 27620 26036
rect 27672 25984 27678 26036
rect 28337 26027 28395 26033
rect 28337 26024 28349 26027
rect 27816 25996 28349 26024
rect 25096 25928 25544 25956
rect 25869 25959 25927 25965
rect 25096 25916 25102 25928
rect 25869 25925 25881 25959
rect 25915 25956 25927 25959
rect 25961 25959 26019 25965
rect 25961 25956 25973 25959
rect 25915 25928 25973 25956
rect 25915 25925 25927 25928
rect 25869 25919 25927 25925
rect 25961 25925 25973 25928
rect 26007 25925 26019 25959
rect 25961 25919 26019 25925
rect 26142 25916 26148 25968
rect 26200 25956 26206 25968
rect 26200 25928 26556 25956
rect 26200 25916 26206 25928
rect 24320 25888 24348 25916
rect 23860 25860 24348 25888
rect 23661 25851 23719 25857
rect 24670 25848 24676 25900
rect 24728 25888 24734 25900
rect 25234 25891 25292 25897
rect 25234 25888 25246 25891
rect 24728 25860 25246 25888
rect 24728 25848 24734 25860
rect 25234 25857 25246 25860
rect 25280 25857 25292 25891
rect 25234 25851 25292 25857
rect 25406 25848 25412 25900
rect 25464 25888 25470 25900
rect 25501 25891 25559 25897
rect 25501 25888 25513 25891
rect 25464 25860 25513 25888
rect 25464 25848 25470 25860
rect 25501 25857 25513 25860
rect 25547 25857 25559 25891
rect 25501 25851 25559 25857
rect 25593 25891 25651 25897
rect 25593 25857 25605 25891
rect 25639 25857 25651 25891
rect 25593 25851 25651 25857
rect 19306 25792 19840 25820
rect 17405 25755 17463 25761
rect 17405 25721 17417 25755
rect 17451 25721 17463 25755
rect 18414 25752 18420 25764
rect 17405 25715 17463 25721
rect 17696 25724 18420 25752
rect 17218 25644 17224 25696
rect 17276 25684 17282 25696
rect 17696 25693 17724 25724
rect 18414 25712 18420 25724
rect 18472 25752 18478 25764
rect 19150 25752 19156 25764
rect 18472 25724 19156 25752
rect 18472 25712 18478 25724
rect 19150 25712 19156 25724
rect 19208 25712 19214 25764
rect 19812 25696 19840 25792
rect 19886 25780 19892 25832
rect 19944 25820 19950 25832
rect 20990 25820 20996 25832
rect 19944 25792 20996 25820
rect 19944 25780 19950 25792
rect 20990 25780 20996 25792
rect 21048 25820 21054 25832
rect 21542 25820 21548 25832
rect 21048 25792 21548 25820
rect 21048 25780 21054 25792
rect 21542 25780 21548 25792
rect 21600 25780 21606 25832
rect 23474 25780 23480 25832
rect 23532 25820 23538 25832
rect 23532 25792 23980 25820
rect 23532 25780 23538 25792
rect 23952 25761 23980 25792
rect 23937 25755 23995 25761
rect 23937 25721 23949 25755
rect 23983 25721 23995 25755
rect 23937 25715 23995 25721
rect 17681 25687 17739 25693
rect 17681 25684 17693 25687
rect 17276 25656 17693 25684
rect 17276 25644 17282 25656
rect 17681 25653 17693 25656
rect 17727 25653 17739 25687
rect 17681 25647 17739 25653
rect 18322 25644 18328 25696
rect 18380 25684 18386 25696
rect 18601 25687 18659 25693
rect 18601 25684 18613 25687
rect 18380 25656 18613 25684
rect 18380 25644 18386 25656
rect 18601 25653 18613 25656
rect 18647 25653 18659 25687
rect 18601 25647 18659 25653
rect 18690 25644 18696 25696
rect 18748 25644 18754 25696
rect 19794 25644 19800 25696
rect 19852 25644 19858 25696
rect 23566 25644 23572 25696
rect 23624 25644 23630 25696
rect 24854 25644 24860 25696
rect 24912 25684 24918 25696
rect 25608 25684 25636 25851
rect 25682 25848 25688 25900
rect 25740 25848 25746 25900
rect 26528 25897 26556 25928
rect 26804 25928 27384 25956
rect 26237 25891 26295 25897
rect 26237 25857 26249 25891
rect 26283 25857 26295 25891
rect 26237 25851 26295 25857
rect 26513 25891 26571 25897
rect 26513 25857 26525 25891
rect 26559 25888 26571 25891
rect 26694 25888 26700 25900
rect 26559 25860 26700 25888
rect 26559 25857 26571 25860
rect 26513 25851 26571 25857
rect 24912 25656 25636 25684
rect 24912 25644 24918 25656
rect 25866 25644 25872 25696
rect 25924 25644 25930 25696
rect 25961 25687 26019 25693
rect 25961 25653 25973 25687
rect 26007 25684 26019 25687
rect 26050 25684 26056 25696
rect 26007 25656 26056 25684
rect 26007 25653 26019 25656
rect 25961 25647 26019 25653
rect 26050 25644 26056 25656
rect 26108 25644 26114 25696
rect 26252 25684 26280 25851
rect 26694 25848 26700 25860
rect 26752 25848 26758 25900
rect 26804 25897 26832 25928
rect 27356 25897 27384 25928
rect 26789 25891 26847 25897
rect 26789 25857 26801 25891
rect 26835 25857 26847 25891
rect 26789 25851 26847 25857
rect 26973 25891 27031 25897
rect 26973 25857 26985 25891
rect 27019 25857 27031 25891
rect 26973 25851 27031 25857
rect 27341 25891 27399 25897
rect 27341 25857 27353 25891
rect 27387 25888 27399 25891
rect 27816 25888 27844 25996
rect 28337 25993 28349 25996
rect 28383 26024 28395 26027
rect 28629 26027 28687 26033
rect 28629 26024 28641 26027
rect 28383 25996 28641 26024
rect 28383 25993 28395 25996
rect 28337 25987 28395 25993
rect 28629 25993 28641 25996
rect 28675 25993 28687 26027
rect 28629 25987 28687 25993
rect 28810 25984 28816 26036
rect 28868 26024 28874 26036
rect 29365 26027 29423 26033
rect 29365 26024 29377 26027
rect 28868 25996 29377 26024
rect 28868 25984 28874 25996
rect 29365 25993 29377 25996
rect 29411 25993 29423 26027
rect 29365 25987 29423 25993
rect 29546 25984 29552 26036
rect 29604 26024 29610 26036
rect 29604 25996 31156 26024
rect 29604 25984 29610 25996
rect 28537 25959 28595 25965
rect 28537 25925 28549 25959
rect 28583 25925 28595 25959
rect 28537 25919 28595 25925
rect 29472 25928 29684 25956
rect 27387 25860 27844 25888
rect 27387 25857 27399 25860
rect 27341 25851 27399 25857
rect 26513 25755 26571 25761
rect 26513 25721 26525 25755
rect 26559 25752 26571 25755
rect 26988 25752 27016 25851
rect 27890 25848 27896 25900
rect 27948 25888 27954 25900
rect 28552 25888 28580 25919
rect 27948 25860 28580 25888
rect 27948 25848 27954 25860
rect 28626 25848 28632 25900
rect 28684 25848 28690 25900
rect 28813 25891 28871 25897
rect 28813 25857 28825 25891
rect 28859 25857 28871 25891
rect 28813 25851 28871 25857
rect 27249 25823 27307 25829
rect 27249 25789 27261 25823
rect 27295 25820 27307 25823
rect 27430 25820 27436 25832
rect 27295 25792 27436 25820
rect 27295 25789 27307 25792
rect 27249 25783 27307 25789
rect 27430 25780 27436 25792
rect 27488 25780 27494 25832
rect 27706 25780 27712 25832
rect 27764 25820 27770 25832
rect 27985 25823 28043 25829
rect 27985 25820 27997 25823
rect 27764 25792 27997 25820
rect 27764 25780 27770 25792
rect 27985 25789 27997 25792
rect 28031 25789 28043 25823
rect 28828 25820 28856 25851
rect 28902 25820 28908 25832
rect 28828 25792 28908 25820
rect 27985 25783 28043 25789
rect 26559 25724 27016 25752
rect 27065 25755 27123 25761
rect 26559 25721 26571 25724
rect 26513 25715 26571 25721
rect 27065 25721 27077 25755
rect 27111 25752 27123 25755
rect 28000 25752 28028 25783
rect 28902 25780 28908 25792
rect 28960 25780 28966 25832
rect 27111 25724 27568 25752
rect 28000 25724 28396 25752
rect 27111 25721 27123 25724
rect 27065 25715 27123 25721
rect 27246 25684 27252 25696
rect 26252 25656 27252 25684
rect 27246 25644 27252 25656
rect 27304 25644 27310 25696
rect 27540 25684 27568 25724
rect 28368 25693 28396 25724
rect 28169 25687 28227 25693
rect 28169 25684 28181 25687
rect 27540 25656 28181 25684
rect 28169 25653 28181 25656
rect 28215 25653 28227 25687
rect 28169 25647 28227 25653
rect 28353 25687 28411 25693
rect 28353 25653 28365 25687
rect 28399 25653 28411 25687
rect 28353 25647 28411 25653
rect 29362 25644 29368 25696
rect 29420 25684 29426 25696
rect 29472 25684 29500 25928
rect 29656 25897 29684 25928
rect 29840 25928 30328 25956
rect 29549 25891 29607 25897
rect 29549 25857 29561 25891
rect 29595 25857 29607 25891
rect 29549 25851 29607 25857
rect 29641 25891 29699 25897
rect 29641 25857 29653 25891
rect 29687 25857 29699 25891
rect 29641 25851 29699 25857
rect 29564 25752 29592 25851
rect 29730 25780 29736 25832
rect 29788 25820 29794 25832
rect 29840 25829 29868 25928
rect 29917 25891 29975 25897
rect 29917 25857 29929 25891
rect 29963 25888 29975 25891
rect 30006 25888 30012 25900
rect 29963 25860 30012 25888
rect 29963 25857 29975 25860
rect 29917 25851 29975 25857
rect 30006 25848 30012 25860
rect 30064 25848 30070 25900
rect 30098 25848 30104 25900
rect 30156 25888 30162 25900
rect 30300 25897 30328 25928
rect 30193 25891 30251 25897
rect 30193 25888 30205 25891
rect 30156 25860 30205 25888
rect 30156 25848 30162 25860
rect 30193 25857 30205 25860
rect 30239 25857 30251 25891
rect 30193 25851 30251 25857
rect 30285 25891 30343 25897
rect 30285 25857 30297 25891
rect 30331 25857 30343 25891
rect 30285 25851 30343 25857
rect 30561 25891 30619 25897
rect 30561 25857 30573 25891
rect 30607 25857 30619 25891
rect 30561 25851 30619 25857
rect 30929 25891 30987 25897
rect 30929 25857 30941 25891
rect 30975 25888 30987 25891
rect 31021 25891 31079 25897
rect 31021 25888 31033 25891
rect 30975 25860 31033 25888
rect 30975 25857 30987 25860
rect 30929 25851 30987 25857
rect 31021 25857 31033 25860
rect 31067 25857 31079 25891
rect 31021 25851 31079 25857
rect 29825 25823 29883 25829
rect 29825 25820 29837 25823
rect 29788 25792 29837 25820
rect 29788 25780 29794 25792
rect 29825 25789 29837 25792
rect 29871 25789 29883 25823
rect 30024 25820 30052 25848
rect 30576 25820 30604 25851
rect 30024 25792 30604 25820
rect 31128 25820 31156 25996
rect 31202 25984 31208 26036
rect 31260 25984 31266 26036
rect 32582 25984 32588 26036
rect 32640 25984 32646 26036
rect 31220 25897 31248 25984
rect 31404 25928 31754 25956
rect 31404 25897 31432 25928
rect 31205 25891 31263 25897
rect 31205 25857 31217 25891
rect 31251 25857 31263 25891
rect 31205 25851 31263 25857
rect 31389 25891 31447 25897
rect 31389 25857 31401 25891
rect 31435 25857 31447 25891
rect 31389 25851 31447 25857
rect 31478 25848 31484 25900
rect 31536 25848 31542 25900
rect 31726 25888 31754 25928
rect 32401 25891 32459 25897
rect 32401 25888 32413 25891
rect 31726 25860 32413 25888
rect 32401 25857 32413 25860
rect 32447 25888 32459 25891
rect 32950 25888 32956 25900
rect 32447 25860 32956 25888
rect 32447 25857 32459 25860
rect 32401 25851 32459 25857
rect 32950 25848 32956 25860
rect 33008 25848 33014 25900
rect 32306 25820 32312 25832
rect 31128 25792 32312 25820
rect 29825 25783 29883 25789
rect 32306 25780 32312 25792
rect 32364 25780 32370 25832
rect 32674 25780 32680 25832
rect 32732 25780 32738 25832
rect 32766 25780 32772 25832
rect 32824 25780 32830 25832
rect 30374 25752 30380 25764
rect 29564 25724 30380 25752
rect 30374 25712 30380 25724
rect 30432 25752 30438 25764
rect 30469 25755 30527 25761
rect 30469 25752 30481 25755
rect 30432 25724 30481 25752
rect 30432 25712 30438 25724
rect 30469 25721 30481 25724
rect 30515 25721 30527 25755
rect 30469 25715 30527 25721
rect 29914 25684 29920 25696
rect 29420 25656 29920 25684
rect 29420 25644 29426 25656
rect 29914 25644 29920 25656
rect 29972 25644 29978 25696
rect 30009 25687 30067 25693
rect 30009 25653 30021 25687
rect 30055 25684 30067 25687
rect 30098 25684 30104 25696
rect 30055 25656 30104 25684
rect 30055 25653 30067 25656
rect 30009 25647 30067 25653
rect 30098 25644 30104 25656
rect 30156 25644 30162 25696
rect 30745 25687 30803 25693
rect 30745 25653 30757 25687
rect 30791 25684 30803 25687
rect 30834 25684 30840 25696
rect 30791 25656 30840 25684
rect 30791 25653 30803 25656
rect 30745 25647 30803 25653
rect 30834 25644 30840 25656
rect 30892 25644 30898 25696
rect 31570 25644 31576 25696
rect 31628 25684 31634 25696
rect 31665 25687 31723 25693
rect 31665 25684 31677 25687
rect 31628 25656 31677 25684
rect 31628 25644 31634 25656
rect 31665 25653 31677 25656
rect 31711 25684 31723 25687
rect 31754 25684 31760 25696
rect 31711 25656 31760 25684
rect 31711 25653 31723 25656
rect 31665 25647 31723 25653
rect 31754 25644 31760 25656
rect 31812 25644 31818 25696
rect 32122 25644 32128 25696
rect 32180 25644 32186 25696
rect 1104 25594 34868 25616
rect 1104 25542 5170 25594
rect 5222 25542 5234 25594
rect 5286 25542 5298 25594
rect 5350 25542 5362 25594
rect 5414 25542 5426 25594
rect 5478 25542 13611 25594
rect 13663 25542 13675 25594
rect 13727 25542 13739 25594
rect 13791 25542 13803 25594
rect 13855 25542 13867 25594
rect 13919 25542 22052 25594
rect 22104 25542 22116 25594
rect 22168 25542 22180 25594
rect 22232 25542 22244 25594
rect 22296 25542 22308 25594
rect 22360 25542 30493 25594
rect 30545 25542 30557 25594
rect 30609 25542 30621 25594
rect 30673 25542 30685 25594
rect 30737 25542 30749 25594
rect 30801 25542 34868 25594
rect 1104 25520 34868 25542
rect 17126 25440 17132 25492
rect 17184 25440 17190 25492
rect 18049 25483 18107 25489
rect 18049 25449 18061 25483
rect 18095 25480 18107 25483
rect 18230 25480 18236 25492
rect 18095 25452 18236 25480
rect 18095 25449 18107 25452
rect 18049 25443 18107 25449
rect 18230 25440 18236 25452
rect 18288 25440 18294 25492
rect 18322 25440 18328 25492
rect 18380 25440 18386 25492
rect 18417 25483 18475 25489
rect 18417 25449 18429 25483
rect 18463 25480 18475 25483
rect 18690 25480 18696 25492
rect 18463 25452 18696 25480
rect 18463 25449 18475 25452
rect 18417 25443 18475 25449
rect 18690 25440 18696 25452
rect 18748 25440 18754 25492
rect 19794 25440 19800 25492
rect 19852 25440 19858 25492
rect 19886 25440 19892 25492
rect 19944 25440 19950 25492
rect 19978 25440 19984 25492
rect 20036 25440 20042 25492
rect 20088 25452 21036 25480
rect 17144 25344 17172 25440
rect 17310 25372 17316 25424
rect 17368 25412 17374 25424
rect 17497 25415 17555 25421
rect 17497 25412 17509 25415
rect 17368 25384 17509 25412
rect 17368 25372 17374 25384
rect 17497 25381 17509 25384
rect 17543 25381 17555 25415
rect 17497 25375 17555 25381
rect 16868 25316 17172 25344
rect 16868 25285 16896 25316
rect 16853 25279 16911 25285
rect 16853 25245 16865 25279
rect 16899 25245 16911 25279
rect 16853 25239 16911 25245
rect 16942 25236 16948 25288
rect 17000 25276 17006 25288
rect 17037 25279 17095 25285
rect 17037 25276 17049 25279
rect 17000 25248 17049 25276
rect 17000 25236 17006 25248
rect 17037 25245 17049 25248
rect 17083 25245 17095 25279
rect 17144 25276 17172 25316
rect 17221 25279 17279 25285
rect 17221 25276 17233 25279
rect 17144 25248 17233 25276
rect 17037 25239 17095 25245
rect 17221 25245 17233 25248
rect 17267 25245 17279 25279
rect 17221 25239 17279 25245
rect 18233 25279 18291 25285
rect 18233 25245 18245 25279
rect 18279 25276 18291 25279
rect 18340 25276 18368 25440
rect 19334 25372 19340 25424
rect 19392 25372 19398 25424
rect 19904 25412 19932 25440
rect 19628 25384 19932 25412
rect 18279 25248 18368 25276
rect 18509 25279 18567 25285
rect 18279 25245 18291 25248
rect 18233 25239 18291 25245
rect 18509 25245 18521 25279
rect 18555 25276 18567 25279
rect 18969 25279 19027 25285
rect 18969 25276 18981 25279
rect 18555 25248 18981 25276
rect 18555 25245 18567 25248
rect 18509 25239 18567 25245
rect 18969 25245 18981 25248
rect 19015 25245 19027 25279
rect 18969 25239 19027 25245
rect 19061 25279 19119 25285
rect 19061 25245 19073 25279
rect 19107 25276 19119 25279
rect 19518 25276 19524 25288
rect 19107 25248 19524 25276
rect 19107 25245 19119 25248
rect 19061 25239 19119 25245
rect 19518 25236 19524 25248
rect 19576 25236 19582 25288
rect 19628 25285 19656 25384
rect 19996 25344 20024 25440
rect 19812 25316 20024 25344
rect 19613 25279 19671 25285
rect 19613 25245 19625 25279
rect 19659 25245 19671 25279
rect 19613 25239 19671 25245
rect 17497 25211 17555 25217
rect 17497 25177 17509 25211
rect 17543 25208 17555 25211
rect 19337 25211 19395 25217
rect 17543 25180 18276 25208
rect 17543 25177 17555 25180
rect 17497 25171 17555 25177
rect 18248 25152 18276 25180
rect 19337 25177 19349 25211
rect 19383 25208 19395 25211
rect 19812 25208 19840 25316
rect 19889 25279 19947 25285
rect 19889 25245 19901 25279
rect 19935 25276 19947 25279
rect 19981 25279 20039 25285
rect 19981 25276 19993 25279
rect 19935 25248 19993 25276
rect 19935 25245 19947 25248
rect 19889 25239 19947 25245
rect 19981 25245 19993 25248
rect 20027 25276 20039 25279
rect 20088 25276 20116 25452
rect 21008 25424 21036 25452
rect 22738 25440 22744 25492
rect 22796 25480 22802 25492
rect 22833 25483 22891 25489
rect 22833 25480 22845 25483
rect 22796 25452 22845 25480
rect 22796 25440 22802 25452
rect 22833 25449 22845 25452
rect 22879 25449 22891 25483
rect 22833 25443 22891 25449
rect 24670 25440 24676 25492
rect 24728 25440 24734 25492
rect 25866 25480 25872 25492
rect 24872 25452 25872 25480
rect 20625 25415 20683 25421
rect 20625 25381 20637 25415
rect 20671 25412 20683 25415
rect 20898 25412 20904 25424
rect 20671 25384 20904 25412
rect 20671 25381 20683 25384
rect 20625 25375 20683 25381
rect 20898 25372 20904 25384
rect 20956 25372 20962 25424
rect 20990 25372 20996 25424
rect 21048 25372 21054 25424
rect 21266 25372 21272 25424
rect 21324 25412 21330 25424
rect 21324 25384 22968 25412
rect 21324 25372 21330 25384
rect 20254 25344 20260 25356
rect 20180 25316 20260 25344
rect 20180 25285 20208 25316
rect 20254 25304 20260 25316
rect 20312 25344 20318 25356
rect 20312 25316 21128 25344
rect 20312 25304 20318 25316
rect 20027 25248 20116 25276
rect 20165 25279 20223 25285
rect 20027 25245 20039 25248
rect 19981 25239 20039 25245
rect 20165 25245 20177 25279
rect 20211 25245 20223 25279
rect 20165 25239 20223 25245
rect 20349 25279 20407 25285
rect 20349 25245 20361 25279
rect 20395 25245 20407 25279
rect 20349 25239 20407 25245
rect 20254 25208 20260 25220
rect 19383 25180 20260 25208
rect 19383 25177 19395 25180
rect 19337 25171 19395 25177
rect 20254 25168 20260 25180
rect 20312 25168 20318 25220
rect 20364 25152 20392 25239
rect 20438 25236 20444 25288
rect 20496 25276 20502 25288
rect 20625 25279 20683 25285
rect 20625 25276 20637 25279
rect 20496 25248 20637 25276
rect 20496 25236 20502 25248
rect 20625 25245 20637 25248
rect 20671 25245 20683 25279
rect 20625 25239 20683 25245
rect 20901 25211 20959 25217
rect 20901 25177 20913 25211
rect 20947 25208 20959 25211
rect 20990 25208 20996 25220
rect 20947 25180 20996 25208
rect 20947 25177 20959 25180
rect 20901 25171 20959 25177
rect 20990 25168 20996 25180
rect 21048 25168 21054 25220
rect 21100 25217 21128 25316
rect 21818 25236 21824 25288
rect 21876 25276 21882 25288
rect 22462 25276 22468 25288
rect 21876 25248 22468 25276
rect 21876 25236 21882 25248
rect 22462 25236 22468 25248
rect 22520 25276 22526 25288
rect 22649 25279 22707 25285
rect 22649 25276 22661 25279
rect 22520 25248 22661 25276
rect 22520 25236 22526 25248
rect 22649 25245 22661 25248
rect 22695 25245 22707 25279
rect 22649 25239 22707 25245
rect 22833 25279 22891 25285
rect 22833 25245 22845 25279
rect 22879 25245 22891 25279
rect 22940 25276 22968 25384
rect 23017 25347 23075 25353
rect 23017 25313 23029 25347
rect 23063 25344 23075 25347
rect 23934 25344 23940 25356
rect 23063 25316 23940 25344
rect 23063 25313 23075 25316
rect 23017 25307 23075 25313
rect 23934 25304 23940 25316
rect 23992 25304 23998 25356
rect 23201 25279 23259 25285
rect 23201 25276 23213 25279
rect 22940 25248 23213 25276
rect 22833 25239 22891 25245
rect 23201 25245 23213 25248
rect 23247 25245 23259 25279
rect 23201 25239 23259 25245
rect 21085 25211 21143 25217
rect 21085 25177 21097 25211
rect 21131 25208 21143 25211
rect 21450 25208 21456 25220
rect 21131 25180 21456 25208
rect 21131 25177 21143 25180
rect 21085 25171 21143 25177
rect 21450 25168 21456 25180
rect 21508 25208 21514 25220
rect 22738 25208 22744 25220
rect 21508 25180 22744 25208
rect 21508 25168 21514 25180
rect 22738 25168 22744 25180
rect 22796 25168 22802 25220
rect 22848 25208 22876 25239
rect 23566 25208 23572 25220
rect 22848 25180 23572 25208
rect 23566 25168 23572 25180
rect 23624 25168 23630 25220
rect 23952 25208 23980 25304
rect 24872 25285 24900 25452
rect 25866 25440 25872 25452
rect 25924 25440 25930 25492
rect 26694 25440 26700 25492
rect 26752 25480 26758 25492
rect 27065 25483 27123 25489
rect 27065 25480 27077 25483
rect 26752 25452 27077 25480
rect 26752 25440 26758 25452
rect 27065 25449 27077 25452
rect 27111 25480 27123 25483
rect 27890 25480 27896 25492
rect 27111 25452 27896 25480
rect 27111 25449 27123 25452
rect 27065 25443 27123 25449
rect 27890 25440 27896 25452
rect 27948 25440 27954 25492
rect 28537 25483 28595 25489
rect 28537 25449 28549 25483
rect 28583 25480 28595 25483
rect 28626 25480 28632 25492
rect 28583 25452 28632 25480
rect 28583 25449 28595 25452
rect 28537 25443 28595 25449
rect 28626 25440 28632 25452
rect 28684 25440 28690 25492
rect 29362 25440 29368 25492
rect 29420 25440 29426 25492
rect 29730 25440 29736 25492
rect 29788 25480 29794 25492
rect 30009 25483 30067 25489
rect 30009 25480 30021 25483
rect 29788 25452 30021 25480
rect 29788 25440 29794 25452
rect 30009 25449 30021 25452
rect 30055 25449 30067 25483
rect 30009 25443 30067 25449
rect 30098 25440 30104 25492
rect 30156 25440 30162 25492
rect 32306 25440 32312 25492
rect 32364 25480 32370 25492
rect 33045 25483 33103 25489
rect 33045 25480 33057 25483
rect 32364 25452 33057 25480
rect 32364 25440 32370 25452
rect 33045 25449 33057 25452
rect 33091 25449 33103 25483
rect 33045 25443 33103 25449
rect 24946 25372 24952 25424
rect 25004 25412 25010 25424
rect 25041 25415 25099 25421
rect 25041 25412 25053 25415
rect 25004 25384 25053 25412
rect 25004 25372 25010 25384
rect 25041 25381 25053 25384
rect 25087 25381 25099 25415
rect 25682 25412 25688 25424
rect 25041 25375 25099 25381
rect 25148 25384 25688 25412
rect 25148 25353 25176 25384
rect 25682 25372 25688 25384
rect 25740 25372 25746 25424
rect 29822 25372 29828 25424
rect 29880 25372 29886 25424
rect 25133 25347 25191 25353
rect 25133 25313 25145 25347
rect 25179 25313 25191 25347
rect 25133 25307 25191 25313
rect 28902 25304 28908 25356
rect 28960 25344 28966 25356
rect 30116 25344 30144 25440
rect 28960 25316 30144 25344
rect 28960 25304 28966 25316
rect 24857 25279 24915 25285
rect 24857 25245 24869 25279
rect 24903 25245 24915 25279
rect 24857 25239 24915 25245
rect 25406 25236 25412 25288
rect 25464 25276 25470 25288
rect 25685 25279 25743 25285
rect 25685 25276 25697 25279
rect 25464 25248 25697 25276
rect 25464 25236 25470 25248
rect 25685 25245 25697 25248
rect 25731 25276 25743 25279
rect 27157 25279 27215 25285
rect 27157 25276 27169 25279
rect 25731 25248 27169 25276
rect 25731 25245 25743 25248
rect 25685 25239 25743 25245
rect 27157 25245 27169 25248
rect 27203 25245 27215 25279
rect 27157 25239 27215 25245
rect 27424 25279 27482 25285
rect 27424 25245 27436 25279
rect 27470 25276 27482 25279
rect 27798 25276 27804 25288
rect 27470 25248 27804 25276
rect 27470 25245 27482 25248
rect 27424 25239 27482 25245
rect 25498 25208 25504 25220
rect 23952 25180 25504 25208
rect 25498 25168 25504 25180
rect 25556 25168 25562 25220
rect 25958 25217 25964 25220
rect 25952 25171 25964 25217
rect 25958 25168 25964 25171
rect 26016 25168 26022 25220
rect 27172 25208 27200 25239
rect 27798 25236 27804 25248
rect 27856 25236 27862 25288
rect 29178 25236 29184 25288
rect 29236 25236 29242 25288
rect 29362 25236 29368 25288
rect 29420 25285 29426 25288
rect 29420 25279 29435 25285
rect 29423 25245 29435 25279
rect 29420 25239 29435 25245
rect 29420 25236 29426 25239
rect 30098 25236 30104 25288
rect 30156 25276 30162 25288
rect 30193 25279 30251 25285
rect 30193 25276 30205 25279
rect 30156 25248 30205 25276
rect 30156 25236 30162 25248
rect 30193 25245 30205 25248
rect 30239 25245 30251 25279
rect 30193 25239 30251 25245
rect 30460 25279 30518 25285
rect 30460 25245 30472 25279
rect 30506 25276 30518 25279
rect 30834 25276 30840 25288
rect 30506 25248 30840 25276
rect 30506 25245 30518 25248
rect 30460 25239 30518 25245
rect 29086 25208 29092 25220
rect 27172 25180 29092 25208
rect 29086 25168 29092 25180
rect 29144 25168 29150 25220
rect 29546 25168 29552 25220
rect 29604 25168 29610 25220
rect 30208 25208 30236 25239
rect 30834 25236 30840 25248
rect 30892 25236 30898 25288
rect 31570 25236 31576 25288
rect 31628 25276 31634 25288
rect 31665 25279 31723 25285
rect 31665 25276 31677 25279
rect 31628 25248 31677 25276
rect 31628 25236 31634 25248
rect 31665 25245 31677 25248
rect 31711 25245 31723 25279
rect 31665 25239 31723 25245
rect 31680 25208 31708 25239
rect 30208 25180 31708 25208
rect 31754 25168 31760 25220
rect 31812 25208 31818 25220
rect 31910 25211 31968 25217
rect 31910 25208 31922 25211
rect 31812 25180 31922 25208
rect 31812 25168 31818 25180
rect 31910 25177 31922 25180
rect 31956 25177 31968 25211
rect 31910 25171 31968 25177
rect 16942 25100 16948 25152
rect 17000 25100 17006 25152
rect 17218 25100 17224 25152
rect 17276 25140 17282 25152
rect 17313 25143 17371 25149
rect 17313 25140 17325 25143
rect 17276 25112 17325 25140
rect 17276 25100 17282 25112
rect 17313 25109 17325 25112
rect 17359 25109 17371 25143
rect 17313 25103 17371 25109
rect 18230 25100 18236 25152
rect 18288 25100 18294 25152
rect 20073 25143 20131 25149
rect 20073 25109 20085 25143
rect 20119 25140 20131 25143
rect 20346 25140 20352 25152
rect 20119 25112 20352 25140
rect 20119 25109 20131 25112
rect 20073 25103 20131 25109
rect 20346 25100 20352 25112
rect 20404 25100 20410 25152
rect 20441 25143 20499 25149
rect 20441 25109 20453 25143
rect 20487 25140 20499 25143
rect 20714 25140 20720 25152
rect 20487 25112 20720 25140
rect 20487 25109 20499 25112
rect 20441 25103 20499 25109
rect 20714 25100 20720 25112
rect 20772 25140 20778 25152
rect 21266 25140 21272 25152
rect 20772 25112 21272 25140
rect 20772 25100 20778 25112
rect 21266 25100 21272 25112
rect 21324 25100 21330 25152
rect 23385 25143 23443 25149
rect 23385 25109 23397 25143
rect 23431 25140 23443 25143
rect 23750 25140 23756 25152
rect 23431 25112 23756 25140
rect 23431 25109 23443 25112
rect 23385 25103 23443 25109
rect 23750 25100 23756 25112
rect 23808 25100 23814 25152
rect 31570 25100 31576 25152
rect 31628 25100 31634 25152
rect 1104 25050 35027 25072
rect 1104 24998 9390 25050
rect 9442 24998 9454 25050
rect 9506 24998 9518 25050
rect 9570 24998 9582 25050
rect 9634 24998 9646 25050
rect 9698 24998 17831 25050
rect 17883 24998 17895 25050
rect 17947 24998 17959 25050
rect 18011 24998 18023 25050
rect 18075 24998 18087 25050
rect 18139 24998 26272 25050
rect 26324 24998 26336 25050
rect 26388 24998 26400 25050
rect 26452 24998 26464 25050
rect 26516 24998 26528 25050
rect 26580 24998 34713 25050
rect 34765 24998 34777 25050
rect 34829 24998 34841 25050
rect 34893 24998 34905 25050
rect 34957 24998 34969 25050
rect 35021 24998 35027 25050
rect 1104 24976 35027 24998
rect 17126 24896 17132 24948
rect 17184 24936 17190 24948
rect 18049 24939 18107 24945
rect 18049 24936 18061 24939
rect 17184 24908 18061 24936
rect 17184 24896 17190 24908
rect 18049 24905 18061 24908
rect 18095 24905 18107 24939
rect 18049 24899 18107 24905
rect 18141 24939 18199 24945
rect 18141 24905 18153 24939
rect 18187 24936 18199 24939
rect 18230 24936 18236 24948
rect 18187 24908 18236 24936
rect 18187 24905 18199 24908
rect 18141 24899 18199 24905
rect 16942 24877 16948 24880
rect 16936 24868 16948 24877
rect 16903 24840 16948 24868
rect 16936 24831 16948 24840
rect 16942 24828 16948 24831
rect 17000 24828 17006 24880
rect 16669 24803 16727 24809
rect 16669 24769 16681 24803
rect 16715 24769 16727 24803
rect 18064 24800 18092 24899
rect 18230 24896 18236 24908
rect 18288 24896 18294 24948
rect 18414 24896 18420 24948
rect 18472 24896 18478 24948
rect 19518 24896 19524 24948
rect 19576 24936 19582 24948
rect 19889 24939 19947 24945
rect 19889 24936 19901 24939
rect 19576 24908 19901 24936
rect 19576 24896 19582 24908
rect 19889 24905 19901 24908
rect 19935 24936 19947 24939
rect 20438 24936 20444 24948
rect 19935 24908 20444 24936
rect 19935 24905 19947 24908
rect 19889 24899 19947 24905
rect 20438 24896 20444 24908
rect 20496 24896 20502 24948
rect 20530 24896 20536 24948
rect 20588 24896 20594 24948
rect 20824 24908 21496 24936
rect 18432 24809 18460 24896
rect 18325 24803 18383 24809
rect 18325 24800 18337 24803
rect 18064 24772 18337 24800
rect 16669 24763 16727 24769
rect 18325 24769 18337 24772
rect 18371 24769 18383 24803
rect 18325 24763 18383 24769
rect 18417 24803 18475 24809
rect 18417 24769 18429 24803
rect 18463 24769 18475 24803
rect 18417 24763 18475 24769
rect 18776 24803 18834 24809
rect 18776 24769 18788 24803
rect 18822 24800 18834 24803
rect 19242 24800 19248 24812
rect 18822 24772 19248 24800
rect 18822 24769 18834 24772
rect 18776 24763 18834 24769
rect 16684 24596 16712 24763
rect 19242 24760 19248 24772
rect 19300 24760 19306 24812
rect 20456 24800 20484 24896
rect 20824 24809 20852 24908
rect 21468 24877 21496 24908
rect 21910 24896 21916 24948
rect 21968 24936 21974 24948
rect 22005 24939 22063 24945
rect 22005 24936 22017 24939
rect 21968 24908 22017 24936
rect 21968 24896 21974 24908
rect 22005 24905 22017 24908
rect 22051 24905 22063 24939
rect 22005 24899 22063 24905
rect 23750 24896 23756 24948
rect 23808 24896 23814 24948
rect 25038 24896 25044 24948
rect 25096 24896 25102 24948
rect 25869 24939 25927 24945
rect 25869 24905 25881 24939
rect 25915 24936 25927 24939
rect 25958 24936 25964 24948
rect 25915 24908 25964 24936
rect 25915 24905 25927 24908
rect 25869 24899 25927 24905
rect 25958 24896 25964 24908
rect 26016 24896 26022 24948
rect 28552 24908 29141 24936
rect 21453 24871 21511 24877
rect 21223 24837 21281 24843
rect 21223 24834 21235 24837
rect 20809 24803 20867 24809
rect 20809 24800 20821 24803
rect 20456 24772 20821 24800
rect 20809 24769 20821 24772
rect 20855 24769 20867 24803
rect 20809 24763 20867 24769
rect 21100 24806 21235 24834
rect 18230 24743 18236 24744
rect 18156 24741 18236 24743
rect 18141 24735 18236 24741
rect 18141 24701 18153 24735
rect 18187 24715 18236 24735
rect 18187 24701 18199 24715
rect 18141 24695 18199 24701
rect 18230 24692 18236 24715
rect 18288 24692 18294 24744
rect 18506 24692 18512 24744
rect 18564 24692 18570 24744
rect 20257 24735 20315 24741
rect 20257 24701 20269 24735
rect 20303 24701 20315 24735
rect 20257 24695 20315 24701
rect 18524 24664 18552 24692
rect 18248 24636 18552 24664
rect 20272 24664 20300 24695
rect 20714 24692 20720 24744
rect 20772 24732 20778 24744
rect 20901 24735 20959 24741
rect 20901 24732 20913 24735
rect 20772 24704 20913 24732
rect 20772 24692 20778 24704
rect 20901 24701 20913 24704
rect 20947 24701 20959 24735
rect 20901 24695 20959 24701
rect 20346 24664 20352 24676
rect 20272 24636 20352 24664
rect 16942 24596 16948 24608
rect 16684 24568 16948 24596
rect 16942 24556 16948 24568
rect 17000 24596 17006 24608
rect 18248 24596 18276 24636
rect 20346 24624 20352 24636
rect 20404 24664 20410 24676
rect 21100 24664 21128 24806
rect 21223 24803 21235 24806
rect 21269 24803 21281 24837
rect 21453 24837 21465 24871
rect 21499 24837 21511 24871
rect 21453 24831 21511 24837
rect 21223 24797 21281 24803
rect 21542 24760 21548 24812
rect 21600 24800 21606 24812
rect 21821 24803 21879 24809
rect 21821 24800 21833 24803
rect 21600 24772 21833 24800
rect 21600 24760 21606 24772
rect 21821 24769 21833 24772
rect 21867 24769 21879 24803
rect 21821 24763 21879 24769
rect 22554 24760 22560 24812
rect 22612 24800 22618 24812
rect 22833 24803 22891 24809
rect 22833 24800 22845 24803
rect 22612 24772 22845 24800
rect 22612 24760 22618 24772
rect 22833 24769 22845 24772
rect 22879 24800 22891 24803
rect 23768 24800 23796 24896
rect 24121 24803 24179 24809
rect 24121 24800 24133 24803
rect 22879 24772 23428 24800
rect 23768 24772 24133 24800
rect 22879 24769 22891 24772
rect 22833 24763 22891 24769
rect 23017 24735 23075 24741
rect 23017 24701 23029 24735
rect 23063 24732 23075 24735
rect 23400 24732 23428 24772
rect 24121 24769 24133 24772
rect 24167 24769 24179 24803
rect 24121 24763 24179 24769
rect 24946 24760 24952 24812
rect 25004 24760 25010 24812
rect 26050 24760 26056 24812
rect 26108 24760 26114 24812
rect 26329 24803 26387 24809
rect 26329 24769 26341 24803
rect 26375 24800 26387 24803
rect 26694 24800 26700 24812
rect 26375 24772 26700 24800
rect 26375 24769 26387 24772
rect 26329 24763 26387 24769
rect 26694 24760 26700 24772
rect 26752 24760 26758 24812
rect 27430 24760 27436 24812
rect 27488 24760 27494 24812
rect 28353 24803 28411 24809
rect 28353 24800 28365 24803
rect 28092 24772 28365 24800
rect 26237 24735 26295 24741
rect 23063 24704 23244 24732
rect 23400 24704 25176 24732
rect 23063 24701 23075 24704
rect 23017 24695 23075 24701
rect 20404 24636 21128 24664
rect 20404 24624 20410 24636
rect 23216 24608 23244 24704
rect 25148 24608 25176 24704
rect 26237 24701 26249 24735
rect 26283 24732 26295 24735
rect 27448 24732 27476 24760
rect 26283 24704 27476 24732
rect 26283 24701 26295 24704
rect 26237 24695 26295 24701
rect 26142 24624 26148 24676
rect 26200 24664 26206 24676
rect 28092 24664 28120 24772
rect 28353 24769 28365 24772
rect 28399 24769 28411 24803
rect 28353 24763 28411 24769
rect 28169 24735 28227 24741
rect 28169 24701 28181 24735
rect 28215 24732 28227 24735
rect 28552 24732 28580 24908
rect 29113 24868 29141 24908
rect 29178 24896 29184 24948
rect 29236 24936 29242 24948
rect 30009 24939 30067 24945
rect 30009 24936 30021 24939
rect 29236 24908 30021 24936
rect 29236 24896 29242 24908
rect 30009 24905 30021 24908
rect 30055 24905 30067 24939
rect 30009 24899 30067 24905
rect 29546 24868 29552 24880
rect 28644 24840 29049 24868
rect 29113 24840 29552 24868
rect 28644 24809 28672 24840
rect 28902 24809 28908 24812
rect 28629 24803 28687 24809
rect 28629 24769 28641 24803
rect 28675 24769 28687 24803
rect 28629 24763 28687 24769
rect 28896 24763 28908 24809
rect 28902 24760 28908 24763
rect 28960 24760 28966 24812
rect 29021 24800 29049 24840
rect 29546 24828 29552 24840
rect 29604 24828 29610 24880
rect 30024 24800 30052 24899
rect 30374 24896 30380 24948
rect 30432 24936 30438 24948
rect 30469 24939 30527 24945
rect 30469 24936 30481 24939
rect 30432 24908 30481 24936
rect 30432 24896 30438 24908
rect 30469 24905 30481 24908
rect 30515 24905 30527 24939
rect 30469 24899 30527 24905
rect 31754 24896 31760 24948
rect 31812 24896 31818 24948
rect 32125 24871 32183 24877
rect 30760 24840 31524 24868
rect 30760 24809 30788 24840
rect 30101 24803 30159 24809
rect 30101 24800 30113 24803
rect 29021 24772 29684 24800
rect 30024 24772 30113 24800
rect 28215 24704 28580 24732
rect 28215 24701 28227 24704
rect 28169 24695 28227 24701
rect 29656 24664 29684 24772
rect 30101 24769 30113 24772
rect 30147 24769 30159 24803
rect 30101 24763 30159 24769
rect 30285 24803 30343 24809
rect 30285 24769 30297 24803
rect 30331 24769 30343 24803
rect 30285 24763 30343 24769
rect 30745 24803 30803 24809
rect 30745 24769 30757 24803
rect 30791 24769 30803 24803
rect 30745 24763 30803 24769
rect 29730 24692 29736 24744
rect 29788 24732 29794 24744
rect 30303 24732 30331 24763
rect 30834 24760 30840 24812
rect 30892 24800 30898 24812
rect 30892 24772 31064 24800
rect 30892 24760 30898 24772
rect 30926 24732 30932 24744
rect 29788 24704 30932 24732
rect 29788 24692 29794 24704
rect 30926 24692 30932 24704
rect 30984 24692 30990 24744
rect 31036 24732 31064 24772
rect 31110 24760 31116 24812
rect 31168 24760 31174 24812
rect 31202 24760 31208 24812
rect 31260 24760 31266 24812
rect 31496 24809 31524 24840
rect 32125 24837 32137 24871
rect 32171 24837 32183 24871
rect 32125 24831 32183 24837
rect 31297 24803 31355 24809
rect 31297 24769 31309 24803
rect 31343 24769 31355 24803
rect 31297 24763 31355 24769
rect 31389 24803 31447 24809
rect 31389 24769 31401 24803
rect 31435 24769 31447 24803
rect 31389 24763 31447 24769
rect 31481 24803 31539 24809
rect 31481 24769 31493 24803
rect 31527 24800 31539 24803
rect 31570 24800 31576 24812
rect 31527 24772 31576 24800
rect 31527 24769 31539 24772
rect 31481 24763 31539 24769
rect 31220 24732 31248 24760
rect 31036 24704 31248 24732
rect 31202 24664 31208 24676
rect 26200 24636 28672 24664
rect 29656 24636 31208 24664
rect 26200 24624 26206 24636
rect 17000 24568 18276 24596
rect 17000 24556 17006 24568
rect 21082 24556 21088 24608
rect 21140 24556 21146 24608
rect 21266 24556 21272 24608
rect 21324 24556 21330 24608
rect 22646 24556 22652 24608
rect 22704 24596 22710 24608
rect 23106 24596 23112 24608
rect 22704 24568 23112 24596
rect 22704 24556 22710 24568
rect 23106 24556 23112 24568
rect 23164 24556 23170 24608
rect 23198 24556 23204 24608
rect 23256 24556 23262 24608
rect 24302 24556 24308 24608
rect 24360 24556 24366 24608
rect 25130 24556 25136 24608
rect 25188 24556 25194 24608
rect 28534 24556 28540 24608
rect 28592 24556 28598 24608
rect 28644 24596 28672 24636
rect 31202 24624 31208 24636
rect 31260 24624 31266 24676
rect 31312 24664 31340 24763
rect 31404 24732 31432 24763
rect 31570 24760 31576 24772
rect 31628 24760 31634 24812
rect 32140 24732 32168 24831
rect 32306 24760 32312 24812
rect 32364 24800 32370 24812
rect 32401 24803 32459 24809
rect 32401 24800 32413 24803
rect 32364 24772 32413 24800
rect 32364 24760 32370 24772
rect 32401 24769 32413 24772
rect 32447 24769 32459 24803
rect 32401 24763 32459 24769
rect 32490 24760 32496 24812
rect 32548 24760 32554 24812
rect 32585 24803 32643 24809
rect 32585 24769 32597 24803
rect 32631 24800 32643 24803
rect 32674 24800 32680 24812
rect 32631 24772 32680 24800
rect 32631 24769 32643 24772
rect 32585 24763 32643 24769
rect 31404 24704 32168 24732
rect 32214 24692 32220 24744
rect 32272 24732 32278 24744
rect 32600 24732 32628 24763
rect 32674 24760 32680 24772
rect 32732 24760 32738 24812
rect 32858 24760 32864 24812
rect 32916 24760 32922 24812
rect 33042 24760 33048 24812
rect 33100 24800 33106 24812
rect 33137 24803 33195 24809
rect 33137 24800 33149 24803
rect 33100 24772 33149 24800
rect 33100 24760 33106 24772
rect 33137 24769 33149 24772
rect 33183 24769 33195 24803
rect 33137 24763 33195 24769
rect 32272 24704 32628 24732
rect 32272 24692 32278 24704
rect 32122 24664 32128 24676
rect 31312 24636 32128 24664
rect 32122 24624 32128 24636
rect 32180 24624 32186 24676
rect 32953 24667 33011 24673
rect 32953 24664 32965 24667
rect 32416 24636 32965 24664
rect 29546 24596 29552 24608
rect 28644 24568 29552 24596
rect 29546 24556 29552 24568
rect 29604 24556 29610 24608
rect 31018 24556 31024 24608
rect 31076 24556 31082 24608
rect 31220 24596 31248 24624
rect 31478 24596 31484 24608
rect 31220 24568 31484 24596
rect 31478 24556 31484 24568
rect 31536 24596 31542 24608
rect 32416 24596 32444 24636
rect 32953 24633 32965 24636
rect 32999 24633 33011 24667
rect 32953 24627 33011 24633
rect 31536 24568 32444 24596
rect 31536 24556 31542 24568
rect 32674 24556 32680 24608
rect 32732 24596 32738 24608
rect 33318 24596 33324 24608
rect 32732 24568 33324 24596
rect 32732 24556 32738 24568
rect 33318 24556 33324 24568
rect 33376 24556 33382 24608
rect 1104 24506 34868 24528
rect 1104 24454 5170 24506
rect 5222 24454 5234 24506
rect 5286 24454 5298 24506
rect 5350 24454 5362 24506
rect 5414 24454 5426 24506
rect 5478 24454 13611 24506
rect 13663 24454 13675 24506
rect 13727 24454 13739 24506
rect 13791 24454 13803 24506
rect 13855 24454 13867 24506
rect 13919 24454 22052 24506
rect 22104 24454 22116 24506
rect 22168 24454 22180 24506
rect 22232 24454 22244 24506
rect 22296 24454 22308 24506
rect 22360 24454 30493 24506
rect 30545 24454 30557 24506
rect 30609 24454 30621 24506
rect 30673 24454 30685 24506
rect 30737 24454 30749 24506
rect 30801 24454 34868 24506
rect 1104 24432 34868 24454
rect 18414 24352 18420 24404
rect 18472 24352 18478 24404
rect 19242 24352 19248 24404
rect 19300 24352 19306 24404
rect 20993 24395 21051 24401
rect 20993 24361 21005 24395
rect 21039 24392 21051 24395
rect 21082 24392 21088 24404
rect 21039 24364 21088 24392
rect 21039 24361 21051 24364
rect 20993 24355 21051 24361
rect 21082 24352 21088 24364
rect 21140 24352 21146 24404
rect 21542 24352 21548 24404
rect 21600 24392 21606 24404
rect 22373 24395 22431 24401
rect 22373 24392 22385 24395
rect 21600 24364 22385 24392
rect 21600 24352 21606 24364
rect 22373 24361 22385 24364
rect 22419 24361 22431 24395
rect 22373 24355 22431 24361
rect 22554 24352 22560 24404
rect 22612 24352 22618 24404
rect 22738 24352 22744 24404
rect 22796 24392 22802 24404
rect 23017 24395 23075 24401
rect 23017 24392 23029 24395
rect 22796 24364 23029 24392
rect 22796 24352 22802 24364
rect 23017 24361 23029 24364
rect 23063 24361 23075 24395
rect 23017 24355 23075 24361
rect 23106 24352 23112 24404
rect 23164 24392 23170 24404
rect 23477 24395 23535 24401
rect 23477 24392 23489 24395
rect 23164 24364 23489 24392
rect 23164 24352 23170 24364
rect 23477 24361 23489 24364
rect 23523 24361 23535 24395
rect 23477 24355 23535 24361
rect 24302 24352 24308 24404
rect 24360 24352 24366 24404
rect 28534 24352 28540 24404
rect 28592 24352 28598 24404
rect 28902 24352 28908 24404
rect 28960 24392 28966 24404
rect 29089 24395 29147 24401
rect 29089 24392 29101 24395
rect 28960 24364 29101 24392
rect 28960 24352 28966 24364
rect 29089 24361 29101 24364
rect 29135 24361 29147 24395
rect 29089 24355 29147 24361
rect 30009 24395 30067 24401
rect 30009 24361 30021 24395
rect 30055 24392 30067 24395
rect 30834 24392 30840 24404
rect 30055 24364 30840 24392
rect 30055 24361 30067 24364
rect 30009 24355 30067 24361
rect 30834 24352 30840 24364
rect 30892 24352 30898 24404
rect 31018 24352 31024 24404
rect 31076 24352 31082 24404
rect 31202 24352 31208 24404
rect 31260 24352 31266 24404
rect 33318 24352 33324 24404
rect 33376 24352 33382 24404
rect 19613 24327 19671 24333
rect 19613 24293 19625 24327
rect 19659 24324 19671 24327
rect 19659 24296 20576 24324
rect 19659 24293 19671 24296
rect 19613 24287 19671 24293
rect 16942 24216 16948 24268
rect 17000 24256 17006 24268
rect 17037 24259 17095 24265
rect 17037 24256 17049 24259
rect 17000 24228 17049 24256
rect 17000 24216 17006 24228
rect 17037 24225 17049 24228
rect 17083 24225 17095 24259
rect 17037 24219 17095 24225
rect 18230 24216 18236 24268
rect 18288 24256 18294 24268
rect 18874 24256 18880 24268
rect 18288 24228 18880 24256
rect 18288 24216 18294 24228
rect 18874 24216 18880 24228
rect 18932 24216 18938 24268
rect 19518 24216 19524 24268
rect 19576 24256 19582 24268
rect 19705 24259 19763 24265
rect 19705 24256 19717 24259
rect 19576 24228 19717 24256
rect 19576 24216 19582 24228
rect 19705 24225 19717 24228
rect 19751 24225 19763 24259
rect 19705 24219 19763 24225
rect 20548 24256 20576 24296
rect 21910 24284 21916 24336
rect 21968 24284 21974 24336
rect 22572 24324 22600 24352
rect 22204 24296 22600 24324
rect 20742 24256 20944 24264
rect 21177 24259 21235 24265
rect 21177 24256 21189 24259
rect 20548 24236 21189 24256
rect 20548 24228 20770 24236
rect 20916 24228 21189 24236
rect 17310 24197 17316 24200
rect 17304 24188 17316 24197
rect 17271 24160 17316 24188
rect 17304 24151 17316 24160
rect 17310 24148 17316 24151
rect 17368 24148 17374 24200
rect 19334 24148 19340 24200
rect 19392 24188 19398 24200
rect 20548 24197 20576 24228
rect 21177 24225 21189 24228
rect 21223 24256 21235 24259
rect 21928 24256 21956 24284
rect 21223 24228 21956 24256
rect 21223 24225 21235 24228
rect 21177 24219 21235 24225
rect 19429 24191 19487 24197
rect 19429 24188 19441 24191
rect 19392 24160 19441 24188
rect 19392 24148 19398 24160
rect 19429 24157 19441 24160
rect 19475 24157 19487 24191
rect 19429 24151 19487 24157
rect 20441 24191 20499 24197
rect 20441 24157 20453 24191
rect 20487 24157 20499 24191
rect 20441 24151 20499 24157
rect 20533 24191 20591 24197
rect 20533 24157 20545 24191
rect 20579 24157 20591 24191
rect 20533 24151 20591 24157
rect 20625 24191 20683 24197
rect 20625 24157 20637 24191
rect 20671 24157 20683 24191
rect 20625 24151 20683 24157
rect 20162 24012 20168 24064
rect 20220 24012 20226 24064
rect 20456 24052 20484 24151
rect 20640 24120 20668 24151
rect 20714 24148 20720 24200
rect 20772 24188 20778 24200
rect 20809 24191 20867 24197
rect 20809 24188 20821 24191
rect 20772 24160 20821 24188
rect 20772 24148 20778 24160
rect 20809 24157 20821 24160
rect 20855 24157 20867 24191
rect 20809 24151 20867 24157
rect 20898 24148 20904 24200
rect 20956 24148 20962 24200
rect 22204 24197 22232 24296
rect 22646 24284 22652 24336
rect 22704 24284 22710 24336
rect 22833 24327 22891 24333
rect 22833 24293 22845 24327
rect 22879 24293 22891 24327
rect 22833 24287 22891 24293
rect 22664 24256 22692 24284
rect 22572 24228 22692 24256
rect 22848 24256 22876 24287
rect 22949 24256 23060 24264
rect 24320 24256 24348 24352
rect 22848 24236 23336 24256
rect 22848 24228 22977 24236
rect 23032 24228 23336 24236
rect 24320 24228 24808 24256
rect 22572 24197 22600 24228
rect 22005 24191 22063 24197
rect 22005 24157 22017 24191
rect 22051 24157 22063 24191
rect 22005 24151 22063 24157
rect 22189 24191 22247 24197
rect 22189 24157 22201 24191
rect 22235 24157 22247 24191
rect 22189 24151 22247 24157
rect 22557 24191 22615 24197
rect 22557 24157 22569 24191
rect 22603 24157 22615 24191
rect 22557 24151 22615 24157
rect 22649 24191 22707 24197
rect 22649 24157 22661 24191
rect 22695 24157 22707 24191
rect 22649 24151 22707 24157
rect 21177 24123 21235 24129
rect 21177 24120 21189 24123
rect 20640 24092 21189 24120
rect 21177 24089 21189 24092
rect 21223 24089 21235 24123
rect 21177 24083 21235 24089
rect 20990 24052 20996 24064
rect 20456 24024 20996 24052
rect 20990 24012 20996 24024
rect 21048 24052 21054 24064
rect 21450 24052 21456 24064
rect 21048 24024 21456 24052
rect 21048 24012 21054 24024
rect 21450 24012 21456 24024
rect 21508 24012 21514 24064
rect 22020 24052 22048 24151
rect 22097 24123 22155 24129
rect 22097 24089 22109 24123
rect 22143 24120 22155 24123
rect 22664 24120 22692 24151
rect 22922 24148 22928 24200
rect 22980 24148 22986 24200
rect 23308 24197 23336 24228
rect 23201 24191 23259 24197
rect 23201 24188 23213 24191
rect 23032 24160 23213 24188
rect 23032 24120 23060 24160
rect 23201 24157 23213 24160
rect 23247 24157 23259 24191
rect 23201 24151 23259 24157
rect 23293 24191 23351 24197
rect 23293 24157 23305 24191
rect 23339 24157 23351 24191
rect 23293 24151 23351 24157
rect 22143 24092 23060 24120
rect 22143 24089 22155 24092
rect 22097 24083 22155 24089
rect 22738 24052 22744 24064
rect 22020 24024 22744 24052
rect 22738 24012 22744 24024
rect 22796 24012 22802 24064
rect 23106 24012 23112 24064
rect 23164 24052 23170 24064
rect 23308 24052 23336 24151
rect 23566 24148 23572 24200
rect 23624 24148 23630 24200
rect 23842 24148 23848 24200
rect 23900 24148 23906 24200
rect 23937 24191 23995 24197
rect 23937 24157 23949 24191
rect 23983 24157 23995 24191
rect 23937 24151 23995 24157
rect 23952 24120 23980 24151
rect 24670 24148 24676 24200
rect 24728 24148 24734 24200
rect 24780 24188 24808 24228
rect 24929 24191 24987 24197
rect 24929 24188 24941 24191
rect 24780 24160 24941 24188
rect 24929 24157 24941 24160
rect 24975 24157 24987 24191
rect 28552 24188 28580 24352
rect 31036 24256 31064 24352
rect 31220 24324 31248 24352
rect 31220 24296 31754 24324
rect 31726 24256 31754 24296
rect 31941 24259 31999 24265
rect 31941 24256 31953 24259
rect 31036 24228 31524 24256
rect 31726 24228 31953 24256
rect 31496 24197 31524 24228
rect 31941 24225 31953 24228
rect 31987 24225 31999 24259
rect 31941 24219 31999 24225
rect 29273 24191 29331 24197
rect 29273 24188 29285 24191
rect 28552 24160 29285 24188
rect 24929 24151 24987 24157
rect 29273 24157 29285 24160
rect 29319 24157 29331 24191
rect 29273 24151 29331 24157
rect 31205 24191 31263 24197
rect 31205 24157 31217 24191
rect 31251 24157 31263 24191
rect 31205 24151 31263 24157
rect 31481 24191 31539 24197
rect 31481 24157 31493 24191
rect 31527 24157 31539 24191
rect 31481 24151 31539 24157
rect 23952 24092 25452 24120
rect 25424 24064 25452 24092
rect 29546 24080 29552 24132
rect 29604 24120 29610 24132
rect 29917 24123 29975 24129
rect 29917 24120 29929 24123
rect 29604 24092 29929 24120
rect 29604 24080 29610 24092
rect 29917 24089 29929 24092
rect 29963 24089 29975 24123
rect 31220 24120 31248 24151
rect 32030 24120 32036 24132
rect 31220 24092 32036 24120
rect 29917 24083 29975 24089
rect 32030 24080 32036 24092
rect 32088 24080 32094 24132
rect 32208 24123 32266 24129
rect 32208 24089 32220 24123
rect 32254 24120 32266 24123
rect 32582 24120 32588 24132
rect 32254 24092 32588 24120
rect 32254 24089 32266 24092
rect 32208 24083 32266 24089
rect 32582 24080 32588 24092
rect 32640 24080 32646 24132
rect 23164 24024 23336 24052
rect 23164 24012 23170 24024
rect 24118 24012 24124 24064
rect 24176 24012 24182 24064
rect 25406 24012 25412 24064
rect 25464 24012 25470 24064
rect 26050 24012 26056 24064
rect 26108 24012 26114 24064
rect 31018 24012 31024 24064
rect 31076 24012 31082 24064
rect 31294 24012 31300 24064
rect 31352 24012 31358 24064
rect 1104 23962 35027 23984
rect 1104 23910 9390 23962
rect 9442 23910 9454 23962
rect 9506 23910 9518 23962
rect 9570 23910 9582 23962
rect 9634 23910 9646 23962
rect 9698 23910 17831 23962
rect 17883 23910 17895 23962
rect 17947 23910 17959 23962
rect 18011 23910 18023 23962
rect 18075 23910 18087 23962
rect 18139 23910 26272 23962
rect 26324 23910 26336 23962
rect 26388 23910 26400 23962
rect 26452 23910 26464 23962
rect 26516 23910 26528 23962
rect 26580 23910 34713 23962
rect 34765 23910 34777 23962
rect 34829 23910 34841 23962
rect 34893 23910 34905 23962
rect 34957 23910 34969 23962
rect 35021 23910 35027 23962
rect 1104 23888 35027 23910
rect 20162 23808 20168 23860
rect 20220 23808 20226 23860
rect 21450 23808 21456 23860
rect 21508 23808 21514 23860
rect 22738 23808 22744 23860
rect 22796 23848 22802 23860
rect 23198 23848 23204 23860
rect 22796 23820 23204 23848
rect 22796 23808 22802 23820
rect 23198 23808 23204 23820
rect 23256 23808 23262 23860
rect 23566 23848 23572 23860
rect 23308 23820 23572 23848
rect 20180 23780 20208 23808
rect 20318 23783 20376 23789
rect 20318 23780 20330 23783
rect 20180 23752 20330 23780
rect 20318 23749 20330 23752
rect 20364 23749 20376 23783
rect 20318 23743 20376 23749
rect 22922 23740 22928 23792
rect 22980 23780 22986 23792
rect 23308 23780 23336 23820
rect 23566 23808 23572 23820
rect 23624 23808 23630 23860
rect 25130 23808 25136 23860
rect 25188 23808 25194 23860
rect 25590 23808 25596 23860
rect 25648 23848 25654 23860
rect 25869 23851 25927 23857
rect 25869 23848 25881 23851
rect 25648 23820 25881 23848
rect 25648 23808 25654 23820
rect 25869 23817 25881 23820
rect 25915 23817 25927 23851
rect 25869 23811 25927 23817
rect 26789 23851 26847 23857
rect 26789 23817 26801 23851
rect 26835 23817 26847 23851
rect 26789 23811 26847 23817
rect 25317 23783 25375 23789
rect 25317 23780 25329 23783
rect 22980 23752 23336 23780
rect 23492 23752 25329 23780
rect 22980 23740 22986 23752
rect 20073 23715 20131 23721
rect 20073 23681 20085 23715
rect 20119 23712 20131 23715
rect 21821 23715 21879 23721
rect 21821 23712 21833 23715
rect 20119 23684 21833 23712
rect 20119 23681 20131 23684
rect 20073 23675 20131 23681
rect 21821 23681 21833 23684
rect 21867 23681 21879 23715
rect 21821 23675 21879 23681
rect 22088 23715 22146 23721
rect 22088 23681 22100 23715
rect 22134 23712 22146 23715
rect 22370 23712 22376 23724
rect 22134 23684 22376 23712
rect 22134 23681 22146 23684
rect 22088 23675 22146 23681
rect 21836 23508 21864 23675
rect 22370 23672 22376 23684
rect 22428 23672 22434 23724
rect 23492 23721 23520 23752
rect 25317 23749 25329 23752
rect 25363 23780 25375 23783
rect 25406 23780 25412 23792
rect 25363 23752 25412 23780
rect 25363 23749 25375 23752
rect 25317 23743 25375 23749
rect 25406 23740 25412 23752
rect 25464 23780 25470 23792
rect 26142 23780 26148 23792
rect 25464 23752 26148 23780
rect 25464 23740 25470 23752
rect 26142 23740 26148 23752
rect 26200 23740 26206 23792
rect 26804 23780 26832 23811
rect 29822 23808 29828 23860
rect 29880 23808 29886 23860
rect 31018 23848 31024 23860
rect 30576 23820 31024 23848
rect 27218 23783 27276 23789
rect 27218 23780 27230 23783
rect 26804 23752 27230 23780
rect 27218 23749 27230 23752
rect 27264 23749 27276 23783
rect 29840 23780 29868 23808
rect 27218 23743 27276 23749
rect 29564 23752 29868 23780
rect 23477 23715 23535 23721
rect 23477 23681 23489 23715
rect 23523 23681 23535 23715
rect 23477 23675 23535 23681
rect 24020 23715 24078 23721
rect 24020 23681 24032 23715
rect 24066 23712 24078 23715
rect 24394 23712 24400 23724
rect 24066 23684 24400 23712
rect 24066 23681 24078 23684
rect 24020 23675 24078 23681
rect 24394 23672 24400 23684
rect 24452 23672 24458 23724
rect 24486 23672 24492 23724
rect 24544 23712 24550 23724
rect 25685 23715 25743 23721
rect 25685 23712 25697 23715
rect 24544 23684 25697 23712
rect 24544 23672 24550 23684
rect 25685 23681 25697 23684
rect 25731 23681 25743 23715
rect 25685 23675 25743 23681
rect 26510 23672 26516 23724
rect 26568 23672 26574 23724
rect 26605 23715 26663 23721
rect 26605 23681 26617 23715
rect 26651 23712 26663 23715
rect 26786 23712 26792 23724
rect 26651 23684 26792 23712
rect 26651 23681 26663 23684
rect 26605 23675 26663 23681
rect 26786 23672 26792 23684
rect 26844 23672 26850 23724
rect 26973 23715 27031 23721
rect 26973 23681 26985 23715
rect 27019 23712 27031 23715
rect 29270 23712 29276 23724
rect 27019 23684 29276 23712
rect 27019 23681 27031 23684
rect 26973 23675 27031 23681
rect 23658 23604 23664 23656
rect 23716 23604 23722 23656
rect 23753 23647 23811 23653
rect 23753 23613 23765 23647
rect 23799 23613 23811 23647
rect 23753 23607 23811 23613
rect 23382 23536 23388 23588
rect 23440 23576 23446 23588
rect 23768 23576 23796 23607
rect 24854 23604 24860 23656
rect 24912 23644 24918 23656
rect 25866 23644 25872 23656
rect 24912 23616 25872 23644
rect 24912 23604 24918 23616
rect 25866 23604 25872 23616
rect 25924 23644 25930 23656
rect 26988 23644 27016 23675
rect 29270 23672 29276 23684
rect 29328 23672 29334 23724
rect 29564 23721 29592 23752
rect 29549 23715 29607 23721
rect 29549 23681 29561 23715
rect 29595 23681 29607 23715
rect 29549 23675 29607 23681
rect 29638 23672 29644 23724
rect 29696 23672 29702 23724
rect 29825 23715 29883 23721
rect 29825 23681 29837 23715
rect 29871 23712 29883 23715
rect 30101 23715 30159 23721
rect 30101 23712 30113 23715
rect 29871 23684 30113 23712
rect 29871 23681 29883 23684
rect 29825 23675 29883 23681
rect 30101 23681 30113 23684
rect 30147 23681 30159 23715
rect 30101 23675 30159 23681
rect 30190 23672 30196 23724
rect 30248 23712 30254 23724
rect 30576 23721 30604 23820
rect 31018 23808 31024 23820
rect 31076 23808 31082 23860
rect 31294 23808 31300 23860
rect 31352 23808 31358 23860
rect 32582 23808 32588 23860
rect 32640 23808 32646 23860
rect 30828 23783 30886 23789
rect 30828 23749 30840 23783
rect 30874 23780 30886 23783
rect 31312 23780 31340 23808
rect 30874 23752 31340 23780
rect 30874 23749 30886 23752
rect 30828 23743 30886 23749
rect 30561 23715 30619 23721
rect 30561 23712 30573 23715
rect 30248 23684 30573 23712
rect 30248 23672 30254 23684
rect 30561 23681 30573 23684
rect 30607 23681 30619 23715
rect 30561 23675 30619 23681
rect 31938 23672 31944 23724
rect 31996 23712 32002 23724
rect 32309 23715 32367 23721
rect 32309 23712 32321 23715
rect 31996 23684 32321 23712
rect 31996 23672 32002 23684
rect 32309 23681 32321 23684
rect 32355 23681 32367 23715
rect 32309 23675 32367 23681
rect 32493 23715 32551 23721
rect 32493 23681 32505 23715
rect 32539 23712 32551 23715
rect 32769 23715 32827 23721
rect 32769 23712 32781 23715
rect 32539 23684 32781 23712
rect 32539 23681 32551 23684
rect 32493 23675 32551 23681
rect 32769 23681 32781 23684
rect 32815 23681 32827 23715
rect 32769 23675 32827 23681
rect 32125 23647 32183 23653
rect 32125 23644 32137 23647
rect 25924 23616 27016 23644
rect 31956 23616 32137 23644
rect 25924 23604 25930 23616
rect 31956 23585 31984 23616
rect 32125 23613 32137 23616
rect 32171 23644 32183 23647
rect 32214 23644 32220 23656
rect 32171 23616 32220 23644
rect 32171 23613 32183 23616
rect 32125 23607 32183 23613
rect 32214 23604 32220 23616
rect 32272 23604 32278 23656
rect 23440 23548 23796 23576
rect 31941 23579 31999 23585
rect 23440 23536 23446 23548
rect 31941 23545 31953 23579
rect 31987 23545 31999 23579
rect 31941 23539 31999 23545
rect 22922 23508 22928 23520
rect 21836 23480 22928 23508
rect 22922 23468 22928 23480
rect 22980 23468 22986 23520
rect 23290 23468 23296 23520
rect 23348 23468 23354 23520
rect 26326 23468 26332 23520
rect 26384 23468 26390 23520
rect 27890 23468 27896 23520
rect 27948 23508 27954 23520
rect 28353 23511 28411 23517
rect 28353 23508 28365 23511
rect 27948 23480 28365 23508
rect 27948 23468 27954 23480
rect 28353 23477 28365 23480
rect 28399 23477 28411 23511
rect 28353 23471 28411 23477
rect 29914 23468 29920 23520
rect 29972 23468 29978 23520
rect 1104 23418 34868 23440
rect 1104 23366 5170 23418
rect 5222 23366 5234 23418
rect 5286 23366 5298 23418
rect 5350 23366 5362 23418
rect 5414 23366 5426 23418
rect 5478 23366 13611 23418
rect 13663 23366 13675 23418
rect 13727 23366 13739 23418
rect 13791 23366 13803 23418
rect 13855 23366 13867 23418
rect 13919 23366 22052 23418
rect 22104 23366 22116 23418
rect 22168 23366 22180 23418
rect 22232 23366 22244 23418
rect 22296 23366 22308 23418
rect 22360 23366 30493 23418
rect 30545 23366 30557 23418
rect 30609 23366 30621 23418
rect 30673 23366 30685 23418
rect 30737 23366 30749 23418
rect 30801 23366 34868 23418
rect 1104 23344 34868 23366
rect 22281 23307 22339 23313
rect 22281 23273 22293 23307
rect 22327 23304 22339 23307
rect 22370 23304 22376 23316
rect 22327 23276 22376 23304
rect 22327 23273 22339 23276
rect 22281 23267 22339 23273
rect 22370 23264 22376 23276
rect 22428 23264 22434 23316
rect 23017 23307 23075 23313
rect 23017 23273 23029 23307
rect 23063 23304 23075 23307
rect 23106 23304 23112 23316
rect 23063 23276 23112 23304
rect 23063 23273 23075 23276
rect 23017 23267 23075 23273
rect 23106 23264 23112 23276
rect 23164 23264 23170 23316
rect 23566 23264 23572 23316
rect 23624 23264 23630 23316
rect 24394 23264 24400 23316
rect 24452 23264 24458 23316
rect 25498 23264 25504 23316
rect 25556 23264 25562 23316
rect 26050 23264 26056 23316
rect 26108 23304 26114 23316
rect 27525 23307 27583 23313
rect 27525 23304 27537 23307
rect 26108 23276 27537 23304
rect 26108 23264 26114 23276
rect 27525 23273 27537 23276
rect 27571 23273 27583 23307
rect 30190 23304 30196 23316
rect 27525 23267 27583 23273
rect 29288 23276 30196 23304
rect 23201 23239 23259 23245
rect 23201 23205 23213 23239
rect 23247 23205 23259 23239
rect 23201 23199 23259 23205
rect 23216 23168 23244 23199
rect 23750 23196 23756 23248
rect 23808 23236 23814 23248
rect 23808 23208 24992 23236
rect 23808 23196 23814 23208
rect 23842 23168 23848 23180
rect 23216 23140 23848 23168
rect 23842 23128 23848 23140
rect 23900 23168 23906 23180
rect 24964 23168 24992 23208
rect 29288 23180 29316 23276
rect 30190 23264 30196 23276
rect 30248 23264 30254 23316
rect 30926 23264 30932 23316
rect 30984 23264 30990 23316
rect 23900 23140 24072 23168
rect 24964 23140 26004 23168
rect 23900 23128 23906 23140
rect 17034 23060 17040 23112
rect 17092 23100 17098 23112
rect 17313 23103 17371 23109
rect 17313 23100 17325 23103
rect 17092 23072 17325 23100
rect 17092 23060 17098 23072
rect 17313 23069 17325 23072
rect 17359 23069 17371 23103
rect 17313 23063 17371 23069
rect 17497 23103 17555 23109
rect 17497 23069 17509 23103
rect 17543 23100 17555 23103
rect 18322 23100 18328 23112
rect 17543 23072 18328 23100
rect 17543 23069 17555 23072
rect 17497 23063 17555 23069
rect 18322 23060 18328 23072
rect 18380 23060 18386 23112
rect 20622 23060 20628 23112
rect 20680 23060 20686 23112
rect 20714 23060 20720 23112
rect 20772 23060 20778 23112
rect 20898 23060 20904 23112
rect 20956 23100 20962 23112
rect 21726 23100 21732 23112
rect 20956 23072 21732 23100
rect 20956 23060 20962 23072
rect 21726 23060 21732 23072
rect 21784 23060 21790 23112
rect 22465 23103 22523 23109
rect 22465 23069 22477 23103
rect 22511 23100 22523 23103
rect 23290 23100 23296 23112
rect 22511 23072 23296 23100
rect 22511 23069 22523 23072
rect 22465 23063 22523 23069
rect 23290 23060 23296 23072
rect 23348 23060 23354 23112
rect 23477 23103 23535 23109
rect 23477 23069 23489 23103
rect 23523 23100 23535 23103
rect 23750 23100 23756 23112
rect 23523 23072 23756 23100
rect 23523 23069 23535 23072
rect 23477 23063 23535 23069
rect 23750 23060 23756 23072
rect 23808 23060 23814 23112
rect 19794 22992 19800 23044
rect 19852 23032 19858 23044
rect 20358 23035 20416 23041
rect 20358 23032 20370 23035
rect 19852 23004 20370 23032
rect 19852 22992 19858 23004
rect 20358 23001 20370 23004
rect 20404 23001 20416 23035
rect 20732 23032 20760 23060
rect 22370 23032 22376 23044
rect 20732 23004 22376 23032
rect 20358 22995 20416 23001
rect 22370 22992 22376 23004
rect 22428 22992 22434 23044
rect 24044 23041 24072 23140
rect 24118 23060 24124 23112
rect 24176 23100 24182 23112
rect 24581 23103 24639 23109
rect 24581 23100 24593 23103
rect 24176 23072 24593 23100
rect 24176 23060 24182 23072
rect 24581 23069 24593 23072
rect 24627 23069 24639 23103
rect 24581 23063 24639 23069
rect 25406 23060 25412 23112
rect 25464 23060 25470 23112
rect 25866 23060 25872 23112
rect 25924 23060 25930 23112
rect 25976 23100 26004 23140
rect 26896 23140 28028 23168
rect 26896 23100 26924 23140
rect 27525 23103 27583 23109
rect 27525 23100 27537 23103
rect 25976 23072 26924 23100
rect 27264 23072 27537 23100
rect 24029 23035 24087 23041
rect 24029 23001 24041 23035
rect 24075 23032 24087 23035
rect 24854 23032 24860 23044
rect 24075 23004 24860 23032
rect 24075 23001 24087 23004
rect 24029 22995 24087 23001
rect 24854 22992 24860 23004
rect 24912 22992 24918 23044
rect 26136 23035 26194 23041
rect 26136 23001 26148 23035
rect 26182 23032 26194 23035
rect 26326 23032 26332 23044
rect 26182 23004 26332 23032
rect 26182 23001 26194 23004
rect 26136 22995 26194 23001
rect 26326 22992 26332 23004
rect 26384 22992 26390 23044
rect 27264 22976 27292 23072
rect 27525 23069 27537 23072
rect 27571 23069 27583 23103
rect 27525 23063 27583 23069
rect 27617 23103 27675 23109
rect 27617 23069 27629 23103
rect 27663 23069 27675 23103
rect 27617 23063 27675 23069
rect 27801 23103 27859 23109
rect 27801 23069 27813 23103
rect 27847 23100 27859 23103
rect 27890 23100 27896 23112
rect 27847 23072 27896 23100
rect 27847 23069 27859 23072
rect 27801 23063 27859 23069
rect 27632 23032 27660 23063
rect 27890 23060 27896 23072
rect 27948 23060 27954 23112
rect 28000 23100 28028 23140
rect 29270 23128 29276 23180
rect 29328 23128 29334 23180
rect 29549 23103 29607 23109
rect 28000 23072 29224 23100
rect 29196 23044 29224 23072
rect 29549 23069 29561 23103
rect 29595 23100 29607 23103
rect 30374 23100 30380 23112
rect 29595 23072 30380 23100
rect 29595 23069 29607 23072
rect 29549 23063 29607 23069
rect 30374 23060 30380 23072
rect 30432 23060 30438 23112
rect 31202 23060 31208 23112
rect 31260 23060 31266 23112
rect 27632 23004 27936 23032
rect 17402 22924 17408 22976
rect 17460 22924 17466 22976
rect 19058 22924 19064 22976
rect 19116 22964 19122 22976
rect 19245 22967 19303 22973
rect 19245 22964 19257 22967
rect 19116 22936 19257 22964
rect 19116 22924 19122 22936
rect 19245 22933 19257 22936
rect 19291 22933 19303 22967
rect 19245 22927 19303 22933
rect 19978 22924 19984 22976
rect 20036 22964 20042 22976
rect 21818 22964 21824 22976
rect 20036 22936 21824 22964
rect 20036 22924 20042 22936
rect 21818 22924 21824 22936
rect 21876 22924 21882 22976
rect 27246 22924 27252 22976
rect 27304 22924 27310 22976
rect 27338 22924 27344 22976
rect 27396 22924 27402 22976
rect 27908 22973 27936 23004
rect 28994 22992 29000 23044
rect 29052 23041 29058 23044
rect 29052 22995 29064 23041
rect 29052 22992 29058 22995
rect 29178 22992 29184 23044
rect 29236 22992 29242 23044
rect 29816 23035 29874 23041
rect 29816 23001 29828 23035
rect 29862 23032 29874 23035
rect 29914 23032 29920 23044
rect 29862 23004 29920 23032
rect 29862 23001 29874 23004
rect 29816 22995 29874 23001
rect 29914 22992 29920 23004
rect 29972 22992 29978 23044
rect 27893 22967 27951 22973
rect 27893 22933 27905 22967
rect 27939 22964 27951 22967
rect 27982 22964 27988 22976
rect 27939 22936 27988 22964
rect 27939 22933 27951 22936
rect 27893 22927 27951 22933
rect 27982 22924 27988 22936
rect 28040 22924 28046 22976
rect 31018 22924 31024 22976
rect 31076 22924 31082 22976
rect 1104 22874 35027 22896
rect 1104 22822 9390 22874
rect 9442 22822 9454 22874
rect 9506 22822 9518 22874
rect 9570 22822 9582 22874
rect 9634 22822 9646 22874
rect 9698 22822 17831 22874
rect 17883 22822 17895 22874
rect 17947 22822 17959 22874
rect 18011 22822 18023 22874
rect 18075 22822 18087 22874
rect 18139 22822 26272 22874
rect 26324 22822 26336 22874
rect 26388 22822 26400 22874
rect 26452 22822 26464 22874
rect 26516 22822 26528 22874
rect 26580 22822 34713 22874
rect 34765 22822 34777 22874
rect 34829 22822 34841 22874
rect 34893 22822 34905 22874
rect 34957 22822 34969 22874
rect 35021 22822 35027 22874
rect 1104 22800 35027 22822
rect 17402 22720 17408 22772
rect 17460 22720 17466 22772
rect 18322 22720 18328 22772
rect 18380 22720 18386 22772
rect 19146 22763 19204 22769
rect 19146 22729 19158 22763
rect 19192 22760 19204 22763
rect 19794 22760 19800 22772
rect 19192 22732 19800 22760
rect 19192 22729 19204 22732
rect 19146 22723 19204 22729
rect 19794 22720 19800 22732
rect 19852 22720 19858 22772
rect 21726 22720 21732 22772
rect 21784 22760 21790 22772
rect 23014 22760 23020 22772
rect 21784 22732 23020 22760
rect 21784 22720 21790 22732
rect 23014 22720 23020 22732
rect 23072 22760 23078 22772
rect 23072 22732 23336 22760
rect 23072 22720 23078 22732
rect 17212 22695 17270 22701
rect 17212 22661 17224 22695
rect 17258 22692 17270 22695
rect 17420 22692 17448 22720
rect 17258 22664 17448 22692
rect 18340 22692 18368 22720
rect 18877 22695 18935 22701
rect 18340 22664 18736 22692
rect 17258 22661 17270 22664
rect 17212 22655 17270 22661
rect 18708 22633 18736 22664
rect 18877 22661 18889 22695
rect 18923 22692 18935 22695
rect 19245 22695 19303 22701
rect 19245 22692 19257 22695
rect 18923 22664 19257 22692
rect 18923 22661 18935 22664
rect 18877 22655 18935 22661
rect 19245 22661 19257 22664
rect 19291 22661 19303 22695
rect 19245 22655 19303 22661
rect 21637 22695 21695 22701
rect 21637 22661 21649 22695
rect 21683 22692 21695 22695
rect 21683 22664 22324 22692
rect 21683 22661 21695 22664
rect 21637 22655 21695 22661
rect 18601 22627 18659 22633
rect 18601 22593 18613 22627
rect 18647 22593 18659 22627
rect 18601 22587 18659 22593
rect 18693 22627 18751 22633
rect 18693 22593 18705 22627
rect 18739 22624 18751 22627
rect 18782 22624 18788 22636
rect 18739 22596 18788 22624
rect 18739 22593 18751 22596
rect 18693 22587 18751 22593
rect 16942 22516 16948 22568
rect 17000 22516 17006 22568
rect 18616 22500 18644 22587
rect 18782 22584 18788 22596
rect 18840 22624 18846 22636
rect 18969 22627 19027 22633
rect 18969 22624 18981 22627
rect 18840 22596 18981 22624
rect 18840 22584 18846 22596
rect 18969 22593 18981 22596
rect 19015 22593 19027 22627
rect 18969 22587 19027 22593
rect 19058 22584 19064 22636
rect 19116 22584 19122 22636
rect 21358 22584 21364 22636
rect 21416 22584 21422 22636
rect 22094 22584 22100 22636
rect 22152 22584 22158 22636
rect 22296 22633 22324 22664
rect 22370 22652 22376 22704
rect 22428 22692 22434 22704
rect 23308 22692 23336 22732
rect 23382 22720 23388 22772
rect 23440 22720 23446 22772
rect 24946 22760 24952 22772
rect 24504 22732 24952 22760
rect 24504 22692 24532 22732
rect 24946 22720 24952 22732
rect 25004 22720 25010 22772
rect 25406 22720 25412 22772
rect 25464 22760 25470 22772
rect 25777 22763 25835 22769
rect 25777 22760 25789 22763
rect 25464 22732 25789 22760
rect 25464 22720 25470 22732
rect 25777 22729 25789 22732
rect 25823 22729 25835 22763
rect 26142 22760 26148 22772
rect 25777 22723 25835 22729
rect 25884 22732 26148 22760
rect 25884 22701 25912 22732
rect 26142 22720 26148 22732
rect 26200 22720 26206 22772
rect 26513 22763 26571 22769
rect 26513 22729 26525 22763
rect 26559 22760 26571 22763
rect 26602 22760 26608 22772
rect 26559 22732 26608 22760
rect 26559 22729 26571 22732
rect 26513 22723 26571 22729
rect 26602 22720 26608 22732
rect 26660 22720 26666 22772
rect 27525 22763 27583 22769
rect 27525 22729 27537 22763
rect 27571 22760 27583 22763
rect 27982 22760 27988 22772
rect 27571 22732 27988 22760
rect 27571 22729 27583 22732
rect 27525 22723 27583 22729
rect 27982 22720 27988 22732
rect 28040 22760 28046 22772
rect 28040 22732 28672 22760
rect 28040 22720 28046 22732
rect 22428 22664 22508 22692
rect 23308 22664 24532 22692
rect 22428 22652 22434 22664
rect 22480 22633 22508 22664
rect 22189 22627 22247 22633
rect 22189 22593 22201 22627
rect 22235 22593 22247 22627
rect 22189 22587 22247 22593
rect 22281 22627 22339 22633
rect 22281 22593 22293 22627
rect 22327 22593 22339 22627
rect 22281 22587 22339 22593
rect 22465 22627 22523 22633
rect 22465 22593 22477 22627
rect 22511 22593 22523 22627
rect 22465 22587 22523 22593
rect 18874 22516 18880 22568
rect 18932 22516 18938 22568
rect 18598 22448 18604 22500
rect 18656 22488 18662 22500
rect 19076 22488 19104 22584
rect 21637 22559 21695 22565
rect 21637 22556 21649 22559
rect 18656 22460 19104 22488
rect 20824 22528 21649 22556
rect 18656 22448 18662 22460
rect 20824 22432 20852 22528
rect 21637 22525 21649 22528
rect 21683 22556 21695 22559
rect 22204 22556 22232 22587
rect 21683 22528 22232 22556
rect 22480 22556 22508 22587
rect 22922 22584 22928 22636
rect 22980 22624 22986 22636
rect 23201 22627 23259 22633
rect 23201 22624 23213 22627
rect 22980 22596 23213 22624
rect 22980 22584 22986 22596
rect 23201 22593 23213 22596
rect 23247 22624 23259 22627
rect 23382 22624 23388 22636
rect 23247 22596 23388 22624
rect 23247 22593 23259 22596
rect 23201 22587 23259 22593
rect 23382 22584 23388 22596
rect 23440 22584 23446 22636
rect 24504 22633 24532 22664
rect 24581 22695 24639 22701
rect 24581 22661 24593 22695
rect 24627 22692 24639 22695
rect 25501 22695 25559 22701
rect 25501 22692 25513 22695
rect 24627 22664 25513 22692
rect 24627 22661 24639 22664
rect 24581 22655 24639 22661
rect 25501 22661 25513 22664
rect 25547 22692 25559 22695
rect 25869 22695 25927 22701
rect 25869 22692 25881 22695
rect 25547 22664 25881 22692
rect 25547 22661 25559 22664
rect 25501 22655 25559 22661
rect 25869 22661 25881 22664
rect 25915 22661 25927 22695
rect 27433 22695 27491 22701
rect 27433 22692 27445 22695
rect 25869 22655 25927 22661
rect 26160 22664 27445 22692
rect 23753 22627 23811 22633
rect 23753 22593 23765 22627
rect 23799 22593 23811 22627
rect 23753 22587 23811 22593
rect 23845 22627 23903 22633
rect 23845 22593 23857 22627
rect 23891 22593 23903 22627
rect 23845 22587 23903 22593
rect 24489 22627 24547 22633
rect 24489 22593 24501 22627
rect 24535 22593 24547 22627
rect 24949 22627 25007 22633
rect 24949 22624 24961 22627
rect 24489 22587 24547 22593
rect 24596 22596 24961 22624
rect 23658 22556 23664 22568
rect 22480 22528 23664 22556
rect 21683 22525 21695 22528
rect 21637 22519 21695 22525
rect 23658 22516 23664 22528
rect 23716 22516 23722 22568
rect 23768 22488 23796 22587
rect 23860 22556 23888 22587
rect 24596 22556 24624 22596
rect 24949 22593 24961 22596
rect 24995 22624 25007 22627
rect 25406 22624 25412 22636
rect 24995 22596 25412 22624
rect 24995 22593 25007 22596
rect 24949 22587 25007 22593
rect 25406 22584 25412 22596
rect 25464 22584 25470 22636
rect 26050 22584 26056 22636
rect 26108 22624 26114 22636
rect 26160 22633 26188 22664
rect 27433 22661 27445 22664
rect 27479 22661 27491 22695
rect 27433 22655 27491 22661
rect 26145 22627 26203 22633
rect 26145 22624 26157 22627
rect 26108 22596 26157 22624
rect 26108 22584 26114 22596
rect 26145 22593 26157 22596
rect 26191 22593 26203 22627
rect 26145 22587 26203 22593
rect 26329 22627 26387 22633
rect 26329 22593 26341 22627
rect 26375 22624 26387 22627
rect 26694 22624 26700 22636
rect 26375 22596 26700 22624
rect 26375 22593 26387 22596
rect 26329 22587 26387 22593
rect 26694 22584 26700 22596
rect 26752 22584 26758 22636
rect 27617 22627 27675 22633
rect 27617 22593 27629 22627
rect 27663 22624 27675 22627
rect 27890 22624 27896 22636
rect 27663 22596 27896 22624
rect 27663 22593 27675 22596
rect 27617 22587 27675 22593
rect 27890 22584 27896 22596
rect 27948 22584 27954 22636
rect 28644 22633 28672 22732
rect 28994 22720 29000 22772
rect 29052 22720 29058 22772
rect 31018 22720 31024 22772
rect 31076 22720 31082 22772
rect 32030 22720 32036 22772
rect 32088 22760 32094 22772
rect 32493 22763 32551 22769
rect 32493 22760 32505 22763
rect 32088 22732 32505 22760
rect 32088 22720 32094 22732
rect 32493 22729 32505 22732
rect 32539 22760 32551 22763
rect 32539 22732 32904 22760
rect 32539 22729 32551 22732
rect 32493 22723 32551 22729
rect 29546 22652 29552 22704
rect 29604 22652 29610 22704
rect 30736 22695 30794 22701
rect 30736 22661 30748 22695
rect 30782 22692 30794 22695
rect 31036 22692 31064 22720
rect 32876 22704 32904 22732
rect 30782 22664 31064 22692
rect 30782 22661 30794 22664
rect 30736 22655 30794 22661
rect 32858 22652 32864 22704
rect 32916 22652 32922 22704
rect 28077 22627 28135 22633
rect 28077 22593 28089 22627
rect 28123 22624 28135 22627
rect 28537 22627 28595 22633
rect 28537 22624 28549 22627
rect 28123 22596 28549 22624
rect 28123 22593 28135 22596
rect 28077 22587 28135 22593
rect 28537 22593 28549 22596
rect 28583 22593 28595 22627
rect 28537 22587 28595 22593
rect 28629 22627 28687 22633
rect 28629 22593 28641 22627
rect 28675 22593 28687 22627
rect 28629 22587 28687 22593
rect 28813 22627 28871 22633
rect 28813 22593 28825 22627
rect 28859 22593 28871 22627
rect 28813 22587 28871 22593
rect 32401 22627 32459 22633
rect 32401 22593 32413 22627
rect 32447 22624 32459 22627
rect 32766 22624 32772 22636
rect 32447 22596 32772 22624
rect 32447 22593 32459 22596
rect 32401 22587 32459 22593
rect 23860 22528 24624 22556
rect 24762 22516 24768 22568
rect 24820 22516 24826 22568
rect 25317 22559 25375 22565
rect 25317 22525 25329 22559
rect 25363 22556 25375 22559
rect 26234 22556 26240 22568
rect 25363 22528 26240 22556
rect 25363 22525 25375 22528
rect 25317 22519 25375 22525
rect 26234 22516 26240 22528
rect 26292 22556 26298 22568
rect 28092 22556 28120 22587
rect 26292 22528 28120 22556
rect 28261 22559 28319 22565
rect 26292 22516 26298 22528
rect 28261 22525 28273 22559
rect 28307 22556 28319 22559
rect 28828 22556 28856 22587
rect 32766 22584 32772 22596
rect 32824 22584 32830 22636
rect 28307 22528 28856 22556
rect 28307 22525 28319 22528
rect 28261 22519 28319 22525
rect 30374 22516 30380 22568
rect 30432 22556 30438 22568
rect 30469 22559 30527 22565
rect 30469 22556 30481 22559
rect 30432 22528 30481 22556
rect 30432 22516 30438 22528
rect 30469 22525 30481 22528
rect 30515 22525 30527 22559
rect 30469 22519 30527 22525
rect 25038 22488 25044 22500
rect 23768 22460 25044 22488
rect 25038 22448 25044 22460
rect 25096 22448 25102 22500
rect 27246 22448 27252 22500
rect 27304 22448 27310 22500
rect 32214 22448 32220 22500
rect 32272 22488 32278 22500
rect 32677 22491 32735 22497
rect 32677 22488 32689 22491
rect 32272 22460 32689 22488
rect 32272 22448 32278 22460
rect 32677 22457 32689 22460
rect 32723 22457 32735 22491
rect 32677 22451 32735 22457
rect 20806 22380 20812 22432
rect 20864 22380 20870 22432
rect 21450 22380 21456 22432
rect 21508 22380 21514 22432
rect 21818 22380 21824 22432
rect 21876 22380 21882 22432
rect 24029 22423 24087 22429
rect 24029 22389 24041 22423
rect 24075 22420 24087 22423
rect 24302 22420 24308 22432
rect 24075 22392 24308 22420
rect 24075 22389 24087 22392
rect 24029 22383 24087 22389
rect 24302 22380 24308 22392
rect 24360 22380 24366 22432
rect 25130 22380 25136 22432
rect 25188 22380 25194 22432
rect 27798 22380 27804 22432
rect 27856 22380 27862 22432
rect 28350 22380 28356 22432
rect 28408 22380 28414 22432
rect 28718 22380 28724 22432
rect 28776 22420 28782 22432
rect 29825 22423 29883 22429
rect 29825 22420 29837 22423
rect 28776 22392 29837 22420
rect 28776 22380 28782 22392
rect 29825 22389 29837 22392
rect 29871 22420 29883 22423
rect 31110 22420 31116 22432
rect 29871 22392 31116 22420
rect 29871 22389 29883 22392
rect 29825 22383 29883 22389
rect 31110 22380 31116 22392
rect 31168 22420 31174 22432
rect 31386 22420 31392 22432
rect 31168 22392 31392 22420
rect 31168 22380 31174 22392
rect 31386 22380 31392 22392
rect 31444 22380 31450 22432
rect 31754 22380 31760 22432
rect 31812 22420 31818 22432
rect 31849 22423 31907 22429
rect 31849 22420 31861 22423
rect 31812 22392 31861 22420
rect 31812 22380 31818 22392
rect 31849 22389 31861 22392
rect 31895 22389 31907 22423
rect 31849 22383 31907 22389
rect 1104 22330 34868 22352
rect 1104 22278 5170 22330
rect 5222 22278 5234 22330
rect 5286 22278 5298 22330
rect 5350 22278 5362 22330
rect 5414 22278 5426 22330
rect 5478 22278 13611 22330
rect 13663 22278 13675 22330
rect 13727 22278 13739 22330
rect 13791 22278 13803 22330
rect 13855 22278 13867 22330
rect 13919 22278 22052 22330
rect 22104 22278 22116 22330
rect 22168 22278 22180 22330
rect 22232 22278 22244 22330
rect 22296 22278 22308 22330
rect 22360 22278 30493 22330
rect 30545 22278 30557 22330
rect 30609 22278 30621 22330
rect 30673 22278 30685 22330
rect 30737 22278 30749 22330
rect 30801 22278 34868 22330
rect 1104 22256 34868 22278
rect 17218 22176 17224 22228
rect 17276 22216 17282 22228
rect 19978 22216 19984 22228
rect 17276 22188 19984 22216
rect 17276 22176 17282 22188
rect 19978 22176 19984 22188
rect 20036 22176 20042 22228
rect 20622 22176 20628 22228
rect 20680 22176 20686 22228
rect 21358 22176 21364 22228
rect 21416 22176 21422 22228
rect 23106 22216 23112 22228
rect 21744 22188 23112 22216
rect 20640 22148 20668 22176
rect 20640 22120 20760 22148
rect 19705 22083 19763 22089
rect 19705 22080 19717 22083
rect 18524 22052 19717 22080
rect 17037 22015 17095 22021
rect 17037 21981 17049 22015
rect 17083 22012 17095 22015
rect 17126 22012 17132 22024
rect 17083 21984 17132 22012
rect 17083 21981 17095 21984
rect 17037 21975 17095 21981
rect 17126 21972 17132 21984
rect 17184 22012 17190 22024
rect 18524 22012 18552 22052
rect 19705 22049 19717 22052
rect 19751 22049 19763 22083
rect 19705 22043 19763 22049
rect 20732 22080 20760 22120
rect 21744 22089 21772 22188
rect 23106 22176 23112 22188
rect 23164 22176 23170 22228
rect 25866 22176 25872 22228
rect 25924 22216 25930 22228
rect 26329 22219 26387 22225
rect 25924 22188 26096 22216
rect 25924 22176 25930 22188
rect 26068 22089 26096 22188
rect 26329 22185 26341 22219
rect 26375 22185 26387 22219
rect 26329 22179 26387 22185
rect 26344 22092 26372 22179
rect 26694 22176 26700 22228
rect 26752 22176 26758 22228
rect 30374 22176 30380 22228
rect 30432 22176 30438 22228
rect 30653 22219 30711 22225
rect 30653 22185 30665 22219
rect 30699 22216 30711 22219
rect 31202 22216 31208 22228
rect 30699 22188 31208 22216
rect 30699 22185 30711 22188
rect 30653 22179 30711 22185
rect 31202 22176 31208 22188
rect 31260 22176 31266 22228
rect 32766 22176 32772 22228
rect 32824 22216 32830 22228
rect 34333 22219 34391 22225
rect 34333 22216 34345 22219
rect 32824 22188 34345 22216
rect 32824 22176 32830 22188
rect 34333 22185 34345 22188
rect 34379 22185 34391 22219
rect 34333 22179 34391 22185
rect 21729 22083 21787 22089
rect 21729 22080 21741 22083
rect 20732 22052 21741 22080
rect 17184 21984 18552 22012
rect 17184 21972 17190 21984
rect 18598 21972 18604 22024
rect 18656 22012 18662 22024
rect 18656 21984 18701 22012
rect 18656 21972 18662 21984
rect 18782 21972 18788 22024
rect 18840 22012 18846 22024
rect 18877 22015 18935 22021
rect 18877 22012 18889 22015
rect 18840 21984 18889 22012
rect 18840 21972 18846 21984
rect 18877 21981 18889 21984
rect 18923 22012 18935 22015
rect 18966 22012 18972 22024
rect 18923 21984 18972 22012
rect 18923 21981 18935 21984
rect 18877 21975 18935 21981
rect 18966 21972 18972 21984
rect 19024 21972 19030 22024
rect 19720 22012 19748 22043
rect 20732 22012 20760 22052
rect 21729 22049 21741 22052
rect 21775 22049 21787 22083
rect 21729 22043 21787 22049
rect 26053 22083 26111 22089
rect 26053 22049 26065 22083
rect 26099 22049 26111 22083
rect 26053 22043 26111 22049
rect 26326 22040 26332 22092
rect 26384 22040 26390 22092
rect 19720 21984 20760 22012
rect 21637 22015 21695 22021
rect 21637 21981 21649 22015
rect 21683 21981 21695 22015
rect 21637 21975 21695 21981
rect 17304 21947 17362 21953
rect 17304 21913 17316 21947
rect 17350 21944 17362 21947
rect 17350 21916 17724 21944
rect 17350 21913 17362 21916
rect 17304 21907 17362 21913
rect 17696 21888 17724 21916
rect 18322 21904 18328 21956
rect 18380 21944 18386 21956
rect 18693 21947 18751 21953
rect 18380 21916 18644 21944
rect 18380 21904 18386 21916
rect 17678 21836 17684 21888
rect 17736 21836 17742 21888
rect 18417 21879 18475 21885
rect 18417 21845 18429 21879
rect 18463 21876 18475 21879
rect 18506 21876 18512 21888
rect 18463 21848 18512 21876
rect 18463 21845 18475 21848
rect 18417 21839 18475 21845
rect 18506 21836 18512 21848
rect 18564 21836 18570 21888
rect 18616 21876 18644 21916
rect 18693 21913 18705 21947
rect 18739 21944 18751 21947
rect 19426 21944 19432 21956
rect 18739 21916 19432 21944
rect 18739 21913 18751 21916
rect 18693 21907 18751 21913
rect 19426 21904 19432 21916
rect 19484 21904 19490 21956
rect 19972 21947 20030 21953
rect 19972 21913 19984 21947
rect 20018 21944 20030 21947
rect 20346 21944 20352 21956
rect 20018 21916 20352 21944
rect 20018 21913 20030 21916
rect 19972 21907 20030 21913
rect 20346 21904 20352 21916
rect 20404 21904 20410 21956
rect 21361 21947 21419 21953
rect 21361 21944 21373 21947
rect 21100 21916 21373 21944
rect 18782 21876 18788 21888
rect 18616 21848 18788 21876
rect 18782 21836 18788 21848
rect 18840 21836 18846 21888
rect 19061 21879 19119 21885
rect 19061 21845 19073 21879
rect 19107 21876 19119 21879
rect 19886 21876 19892 21888
rect 19107 21848 19892 21876
rect 19107 21845 19119 21848
rect 19061 21839 19119 21845
rect 19886 21836 19892 21848
rect 19944 21836 19950 21888
rect 20714 21836 20720 21888
rect 20772 21876 20778 21888
rect 21100 21885 21128 21916
rect 21361 21913 21373 21916
rect 21407 21913 21419 21947
rect 21652 21944 21680 21975
rect 21818 21972 21824 22024
rect 21876 22012 21882 22024
rect 21985 22015 22043 22021
rect 21985 22012 21997 22015
rect 21876 21984 21997 22012
rect 21876 21972 21882 21984
rect 21985 21981 21997 21984
rect 22031 21981 22043 22015
rect 21985 21975 22043 21981
rect 24302 21972 24308 22024
rect 24360 22012 24366 22024
rect 24581 22015 24639 22021
rect 24581 22012 24593 22015
rect 24360 21984 24593 22012
rect 24360 21972 24366 21984
rect 24581 21981 24593 21984
rect 24627 21981 24639 22015
rect 24581 21975 24639 21981
rect 26142 21972 26148 22024
rect 26200 22012 26206 22024
rect 26605 22015 26663 22021
rect 26605 22012 26617 22015
rect 26200 21984 26617 22012
rect 26200 21972 26206 21984
rect 26605 21981 26617 21984
rect 26651 21981 26663 22015
rect 26712 22012 26740 22176
rect 30392 22148 30420 22176
rect 29564 22120 29776 22148
rect 30392 22120 32168 22148
rect 26786 22040 26792 22092
rect 26844 22080 26850 22092
rect 26973 22083 27031 22089
rect 26973 22080 26985 22083
rect 26844 22052 26985 22080
rect 26844 22040 26850 22052
rect 26973 22049 26985 22052
rect 27019 22049 27031 22083
rect 26973 22043 27031 22049
rect 27246 22040 27252 22092
rect 27304 22080 27310 22092
rect 27341 22083 27399 22089
rect 27341 22080 27353 22083
rect 27304 22052 27353 22080
rect 27304 22040 27310 22052
rect 27341 22049 27353 22052
rect 27387 22049 27399 22083
rect 29564 22080 29592 22120
rect 27341 22043 27399 22049
rect 27816 22052 29592 22080
rect 29748 22080 29776 22120
rect 31665 22083 31723 22089
rect 29748 22052 31524 22080
rect 27157 22015 27215 22021
rect 27157 22012 27169 22015
rect 26712 21984 27169 22012
rect 26605 21975 26663 21981
rect 27157 21981 27169 21984
rect 27203 22012 27215 22015
rect 27816 22012 27844 22052
rect 30484 22024 30512 22052
rect 27203 21984 27844 22012
rect 27203 21981 27215 21984
rect 27157 21975 27215 21981
rect 28166 21972 28172 22024
rect 28224 21972 28230 22024
rect 29914 21972 29920 22024
rect 29972 21972 29978 22024
rect 30377 22015 30435 22021
rect 30377 21981 30389 22015
rect 30423 21981 30435 22015
rect 30377 21975 30435 21981
rect 24029 21947 24087 21953
rect 21652 21916 21956 21944
rect 21361 21907 21419 21913
rect 21928 21888 21956 21916
rect 24029 21913 24041 21947
rect 24075 21944 24087 21947
rect 24075 21916 25728 21944
rect 24075 21913 24087 21916
rect 24029 21907 24087 21913
rect 21085 21879 21143 21885
rect 21085 21876 21097 21879
rect 20772 21848 21097 21876
rect 20772 21836 20778 21848
rect 21085 21845 21097 21848
rect 21131 21845 21143 21879
rect 21085 21839 21143 21845
rect 21542 21836 21548 21888
rect 21600 21836 21606 21888
rect 21910 21836 21916 21888
rect 21968 21836 21974 21888
rect 22554 21836 22560 21888
rect 22612 21876 22618 21888
rect 23109 21879 23167 21885
rect 23109 21876 23121 21879
rect 22612 21848 23121 21876
rect 22612 21836 22618 21848
rect 23109 21845 23121 21848
rect 23155 21845 23167 21879
rect 23109 21839 23167 21845
rect 23382 21836 23388 21888
rect 23440 21876 23446 21888
rect 23937 21879 23995 21885
rect 23937 21876 23949 21879
rect 23440 21848 23949 21876
rect 23440 21836 23446 21848
rect 23937 21845 23949 21848
rect 23983 21845 23995 21879
rect 23937 21839 23995 21845
rect 24394 21836 24400 21888
rect 24452 21836 24458 21888
rect 24673 21879 24731 21885
rect 24673 21845 24685 21879
rect 24719 21876 24731 21879
rect 25314 21876 25320 21888
rect 24719 21848 25320 21876
rect 24719 21845 24731 21848
rect 24673 21839 24731 21845
rect 25314 21836 25320 21848
rect 25372 21836 25378 21888
rect 25700 21876 25728 21916
rect 25774 21904 25780 21956
rect 25832 21953 25838 21956
rect 25832 21907 25844 21953
rect 25832 21904 25838 21907
rect 26326 21904 26332 21956
rect 26384 21944 26390 21956
rect 27522 21944 27528 21956
rect 26384 21916 27528 21944
rect 26384 21904 26390 21916
rect 27522 21904 27528 21916
rect 27580 21944 27586 21956
rect 29638 21944 29644 21956
rect 27580 21916 29644 21944
rect 27580 21904 27586 21916
rect 29638 21904 29644 21916
rect 29696 21904 29702 21956
rect 30392 21944 30420 21975
rect 30466 21972 30472 22024
rect 30524 21972 30530 22024
rect 31021 22015 31079 22021
rect 31021 21981 31033 22015
rect 31067 21981 31079 22015
rect 31021 21975 31079 21981
rect 31036 21944 31064 21975
rect 31110 21972 31116 22024
rect 31168 21972 31174 22024
rect 31202 21972 31208 22024
rect 31260 21972 31266 22024
rect 31386 21972 31392 22024
rect 31444 21972 31450 22024
rect 31496 22012 31524 22052
rect 31665 22049 31677 22083
rect 31711 22080 31723 22083
rect 31754 22080 31760 22092
rect 31711 22052 31760 22080
rect 31711 22049 31723 22052
rect 31665 22043 31723 22049
rect 31754 22040 31760 22052
rect 31812 22040 31818 22092
rect 31849 22015 31907 22021
rect 31849 22012 31861 22015
rect 31496 21984 31861 22012
rect 31849 21981 31861 21984
rect 31895 22012 31907 22015
rect 31938 22012 31944 22024
rect 31895 21984 31944 22012
rect 31895 21981 31907 21984
rect 31849 21975 31907 21981
rect 31938 21972 31944 21984
rect 31996 21972 32002 22024
rect 32140 22021 32168 22120
rect 32125 22015 32183 22021
rect 32125 21981 32137 22015
rect 32171 22012 32183 22015
rect 32214 22012 32220 22024
rect 32171 21984 32220 22012
rect 32171 21981 32183 21984
rect 32125 21975 32183 21981
rect 32214 21972 32220 21984
rect 32272 21972 32278 22024
rect 33781 22015 33839 22021
rect 33781 22012 33793 22015
rect 32324 21984 33793 22012
rect 32033 21947 32091 21953
rect 30392 21916 31340 21944
rect 31312 21888 31340 21916
rect 32033 21913 32045 21947
rect 32079 21944 32091 21947
rect 32324 21944 32352 21984
rect 33781 21981 33793 21984
rect 33827 21981 33839 22015
rect 33781 21975 33839 21981
rect 34517 22015 34575 22021
rect 34517 21981 34529 22015
rect 34563 22012 34575 22015
rect 34882 22012 34888 22024
rect 34563 21984 34888 22012
rect 34563 21981 34575 21984
rect 34517 21975 34575 21981
rect 34882 21972 34888 21984
rect 34940 21972 34946 22024
rect 32079 21916 32352 21944
rect 32392 21947 32450 21953
rect 32079 21913 32091 21916
rect 32033 21907 32091 21913
rect 32392 21913 32404 21947
rect 32438 21944 32450 21947
rect 32438 21916 33640 21944
rect 32438 21913 32450 21916
rect 32392 21907 32450 21913
rect 26878 21876 26884 21888
rect 25700 21848 26884 21876
rect 26878 21836 26884 21848
rect 26936 21836 26942 21888
rect 28350 21836 28356 21888
rect 28408 21836 28414 21888
rect 30101 21879 30159 21885
rect 30101 21845 30113 21879
rect 30147 21876 30159 21879
rect 30190 21876 30196 21888
rect 30147 21848 30196 21876
rect 30147 21845 30159 21848
rect 30101 21839 30159 21845
rect 30190 21836 30196 21848
rect 30248 21836 30254 21888
rect 30745 21879 30803 21885
rect 30745 21845 30757 21879
rect 30791 21876 30803 21879
rect 30834 21876 30840 21888
rect 30791 21848 30840 21876
rect 30791 21845 30803 21848
rect 30745 21839 30803 21845
rect 30834 21836 30840 21848
rect 30892 21836 30898 21888
rect 31294 21836 31300 21888
rect 31352 21836 31358 21888
rect 33502 21836 33508 21888
rect 33560 21836 33566 21888
rect 33612 21885 33640 21916
rect 33597 21879 33655 21885
rect 33597 21845 33609 21879
rect 33643 21845 33655 21879
rect 33597 21839 33655 21845
rect 1104 21786 35027 21808
rect 1104 21734 9390 21786
rect 9442 21734 9454 21786
rect 9506 21734 9518 21786
rect 9570 21734 9582 21786
rect 9634 21734 9646 21786
rect 9698 21734 17831 21786
rect 17883 21734 17895 21786
rect 17947 21734 17959 21786
rect 18011 21734 18023 21786
rect 18075 21734 18087 21786
rect 18139 21734 26272 21786
rect 26324 21734 26336 21786
rect 26388 21734 26400 21786
rect 26452 21734 26464 21786
rect 26516 21734 26528 21786
rect 26580 21734 34713 21786
rect 34765 21734 34777 21786
rect 34829 21734 34841 21786
rect 34893 21734 34905 21786
rect 34957 21734 34969 21786
rect 35021 21734 35027 21786
rect 1104 21712 35027 21734
rect 17678 21632 17684 21684
rect 17736 21632 17742 21684
rect 18322 21681 18328 21684
rect 18309 21675 18328 21681
rect 18309 21641 18321 21675
rect 18309 21635 18328 21641
rect 18322 21632 18328 21635
rect 18380 21632 18386 21684
rect 19610 21672 19616 21684
rect 18616 21644 19616 21672
rect 17218 21564 17224 21616
rect 17276 21604 17282 21616
rect 17405 21607 17463 21613
rect 17405 21604 17417 21607
rect 17276 21576 17417 21604
rect 17276 21564 17282 21576
rect 17405 21573 17417 21576
rect 17451 21573 17463 21607
rect 17405 21567 17463 21573
rect 18506 21564 18512 21616
rect 18564 21604 18570 21616
rect 18616 21613 18644 21644
rect 19610 21632 19616 21644
rect 19668 21632 19674 21684
rect 20346 21632 20352 21684
rect 20404 21632 20410 21684
rect 21634 21632 21640 21684
rect 21692 21632 21698 21684
rect 22370 21632 22376 21684
rect 22428 21632 22434 21684
rect 24581 21675 24639 21681
rect 24581 21672 24593 21675
rect 24504 21644 24593 21672
rect 18601 21607 18659 21613
rect 18601 21604 18613 21607
rect 18564 21576 18613 21604
rect 18564 21564 18570 21576
rect 18601 21573 18613 21576
rect 18647 21573 18659 21607
rect 18601 21567 18659 21573
rect 18966 21564 18972 21616
rect 19024 21564 19030 21616
rect 19153 21607 19211 21613
rect 19153 21573 19165 21607
rect 19199 21604 19211 21607
rect 19199 21576 20116 21604
rect 19199 21573 19211 21576
rect 19153 21567 19211 21573
rect 17681 21539 17739 21545
rect 17681 21505 17693 21539
rect 17727 21505 17739 21539
rect 17681 21499 17739 21505
rect 17696 21468 17724 21499
rect 18690 21496 18696 21548
rect 18748 21536 18754 21548
rect 18785 21539 18843 21545
rect 18785 21536 18797 21539
rect 18748 21508 18797 21536
rect 18748 21496 18754 21508
rect 18785 21505 18797 21508
rect 18831 21505 18843 21539
rect 18785 21499 18843 21505
rect 18877 21539 18935 21545
rect 18877 21505 18889 21539
rect 18923 21536 18935 21539
rect 18984 21536 19012 21564
rect 18923 21508 19012 21536
rect 19337 21539 19395 21545
rect 18923 21505 18935 21508
rect 18877 21499 18935 21505
rect 19337 21505 19349 21539
rect 19383 21505 19395 21539
rect 19337 21499 19395 21505
rect 18708 21468 18736 21496
rect 19352 21468 19380 21499
rect 19426 21496 19432 21548
rect 19484 21496 19490 21548
rect 19702 21496 19708 21548
rect 19760 21496 19766 21548
rect 19886 21496 19892 21548
rect 19944 21496 19950 21548
rect 20088 21545 20116 21576
rect 20254 21564 20260 21616
rect 20312 21604 20318 21616
rect 21269 21607 21327 21613
rect 21269 21604 21281 21607
rect 20312 21576 20944 21604
rect 20312 21564 20318 21576
rect 20916 21545 20944 21576
rect 21100 21576 21281 21604
rect 20073 21539 20131 21545
rect 20073 21505 20085 21539
rect 20119 21505 20131 21539
rect 20073 21499 20131 21505
rect 20533 21539 20591 21545
rect 20533 21505 20545 21539
rect 20579 21505 20591 21539
rect 20533 21499 20591 21505
rect 20901 21539 20959 21545
rect 20901 21505 20913 21539
rect 20947 21536 20959 21539
rect 20990 21536 20996 21548
rect 20947 21508 20996 21536
rect 20947 21505 20959 21508
rect 20901 21499 20959 21505
rect 17696 21440 18644 21468
rect 18616 21409 18644 21440
rect 18708 21440 19380 21468
rect 17589 21403 17647 21409
rect 17589 21369 17601 21403
rect 17635 21400 17647 21403
rect 18601 21403 18659 21409
rect 17635 21372 18092 21400
rect 17635 21369 17647 21372
rect 17589 21363 17647 21369
rect 18064 21344 18092 21372
rect 18601 21369 18613 21403
rect 18647 21369 18659 21403
rect 18601 21363 18659 21369
rect 18046 21292 18052 21344
rect 18104 21332 18110 21344
rect 18141 21335 18199 21341
rect 18141 21332 18153 21335
rect 18104 21304 18153 21332
rect 18104 21292 18110 21304
rect 18141 21301 18153 21304
rect 18187 21301 18199 21335
rect 18141 21295 18199 21301
rect 18325 21335 18383 21341
rect 18325 21301 18337 21335
rect 18371 21332 18383 21335
rect 18708 21332 18736 21440
rect 19444 21400 19472 21496
rect 19794 21428 19800 21480
rect 19852 21428 19858 21480
rect 20548 21400 20576 21499
rect 20990 21496 20996 21508
rect 21048 21496 21054 21548
rect 21100 21545 21128 21576
rect 21269 21573 21281 21576
rect 21315 21573 21327 21607
rect 21269 21567 21327 21573
rect 21485 21607 21543 21613
rect 21485 21573 21497 21607
rect 21531 21604 21543 21607
rect 21910 21604 21916 21616
rect 21531 21576 21916 21604
rect 21531 21573 21543 21576
rect 21485 21567 21543 21573
rect 21085 21539 21143 21545
rect 21085 21505 21097 21539
rect 21131 21505 21143 21539
rect 21085 21499 21143 21505
rect 20714 21428 20720 21480
rect 20772 21468 20778 21480
rect 20809 21471 20867 21477
rect 20809 21468 20821 21471
rect 20772 21440 20821 21468
rect 20772 21428 20778 21440
rect 20809 21437 20821 21440
rect 20855 21468 20867 21471
rect 21100 21468 21128 21499
rect 21174 21496 21180 21548
rect 21232 21496 21238 21548
rect 21284 21536 21312 21567
rect 21910 21564 21916 21576
rect 21968 21564 21974 21616
rect 23376 21607 23434 21613
rect 23376 21573 23388 21607
rect 23422 21604 23434 21607
rect 24394 21604 24400 21616
rect 23422 21576 24400 21604
rect 23422 21573 23434 21576
rect 23376 21567 23434 21573
rect 24394 21564 24400 21576
rect 24452 21564 24458 21616
rect 22373 21539 22431 21545
rect 22373 21536 22385 21539
rect 21284 21508 22385 21536
rect 22373 21505 22385 21508
rect 22419 21505 22431 21539
rect 22373 21499 22431 21505
rect 22554 21496 22560 21548
rect 22612 21536 22618 21548
rect 22833 21539 22891 21545
rect 22833 21536 22845 21539
rect 22612 21508 22845 21536
rect 22612 21496 22618 21508
rect 22833 21505 22845 21508
rect 22879 21505 22891 21539
rect 22833 21499 22891 21505
rect 23014 21496 23020 21548
rect 23072 21496 23078 21548
rect 23934 21496 23940 21548
rect 23992 21536 23998 21548
rect 24504 21536 24532 21644
rect 24581 21641 24593 21644
rect 24627 21641 24639 21675
rect 24581 21635 24639 21641
rect 24762 21632 24768 21684
rect 24820 21672 24826 21684
rect 25590 21672 25596 21684
rect 24820 21644 25596 21672
rect 24820 21632 24826 21644
rect 25590 21632 25596 21644
rect 25648 21632 25654 21684
rect 25774 21632 25780 21684
rect 25832 21672 25838 21684
rect 25869 21675 25927 21681
rect 25869 21672 25881 21675
rect 25832 21644 25881 21672
rect 25832 21632 25838 21644
rect 25869 21641 25881 21644
rect 25915 21641 25927 21675
rect 25869 21635 25927 21641
rect 31110 21632 31116 21684
rect 31168 21672 31174 21684
rect 32125 21675 32183 21681
rect 32125 21672 32137 21675
rect 31168 21644 32137 21672
rect 31168 21632 31174 21644
rect 32125 21641 32137 21644
rect 32171 21641 32183 21675
rect 32125 21635 32183 21641
rect 33413 21675 33471 21681
rect 33413 21641 33425 21675
rect 33459 21672 33471 21675
rect 33502 21672 33508 21684
rect 33459 21644 33508 21672
rect 33459 21641 33471 21644
rect 33413 21635 33471 21641
rect 33502 21632 33508 21644
rect 33560 21632 33566 21684
rect 25038 21564 25044 21616
rect 25096 21564 25102 21616
rect 25314 21564 25320 21616
rect 25372 21604 25378 21616
rect 25372 21576 26004 21604
rect 25372 21564 25378 21576
rect 23992 21508 24532 21536
rect 23992 21496 23998 21508
rect 25130 21496 25136 21548
rect 25188 21536 25194 21548
rect 25976 21545 26004 21576
rect 28350 21564 28356 21616
rect 28408 21604 28414 21616
rect 30190 21613 30196 21616
rect 29558 21607 29616 21613
rect 29558 21604 29570 21607
rect 28408 21576 29570 21604
rect 28408 21564 28414 21576
rect 29558 21573 29570 21576
rect 29604 21573 29616 21607
rect 29558 21567 29616 21573
rect 30184 21567 30196 21613
rect 30190 21564 30196 21567
rect 30248 21564 30254 21616
rect 31202 21564 31208 21616
rect 31260 21564 31266 21616
rect 32416 21576 33180 21604
rect 25685 21539 25743 21545
rect 25685 21536 25697 21539
rect 25188 21508 25697 21536
rect 25188 21496 25194 21508
rect 25685 21505 25697 21508
rect 25731 21505 25743 21539
rect 25685 21499 25743 21505
rect 25961 21539 26019 21545
rect 25961 21505 25973 21539
rect 26007 21505 26019 21539
rect 25961 21499 26019 21505
rect 26145 21539 26203 21545
rect 26145 21505 26157 21539
rect 26191 21505 26203 21539
rect 26145 21499 26203 21505
rect 20855 21440 21128 21468
rect 20855 21437 20867 21440
rect 20809 21431 20867 21437
rect 21542 21428 21548 21480
rect 21600 21428 21606 21480
rect 21821 21471 21879 21477
rect 21821 21437 21833 21471
rect 21867 21468 21879 21471
rect 21910 21468 21916 21480
rect 21867 21440 21916 21468
rect 21867 21437 21879 21440
rect 21821 21431 21879 21437
rect 21910 21428 21916 21440
rect 21968 21428 21974 21480
rect 22465 21471 22523 21477
rect 22465 21468 22477 21471
rect 22066 21440 22477 21468
rect 20901 21403 20959 21409
rect 20901 21400 20913 21403
rect 19444 21372 20484 21400
rect 20548 21372 20913 21400
rect 20456 21344 20484 21372
rect 20901 21369 20913 21372
rect 20947 21369 20959 21403
rect 20901 21363 20959 21369
rect 21560 21400 21588 21428
rect 22066 21400 22094 21440
rect 22465 21437 22477 21440
rect 22511 21468 22523 21471
rect 22649 21471 22707 21477
rect 22649 21468 22661 21471
rect 22511 21440 22661 21468
rect 22511 21437 22523 21440
rect 22465 21431 22523 21437
rect 22649 21437 22661 21440
rect 22695 21437 22707 21471
rect 23106 21468 23112 21480
rect 22649 21431 22707 21437
rect 22848 21440 23112 21468
rect 21560 21372 22094 21400
rect 18371 21304 18736 21332
rect 18371 21301 18383 21304
rect 18325 21295 18383 21301
rect 19610 21292 19616 21344
rect 19668 21292 19674 21344
rect 20254 21292 20260 21344
rect 20312 21292 20318 21344
rect 20438 21292 20444 21344
rect 20496 21292 20502 21344
rect 20717 21335 20775 21341
rect 20717 21301 20729 21335
rect 20763 21332 20775 21335
rect 20806 21332 20812 21344
rect 20763 21304 20812 21332
rect 20763 21301 20775 21304
rect 20717 21295 20775 21301
rect 20806 21292 20812 21304
rect 20864 21292 20870 21344
rect 21453 21335 21511 21341
rect 21453 21301 21465 21335
rect 21499 21332 21511 21335
rect 21560 21332 21588 21372
rect 22848 21344 22876 21440
rect 23106 21428 23112 21440
rect 23164 21428 23170 21480
rect 24504 21440 25544 21468
rect 24504 21344 24532 21440
rect 24762 21360 24768 21412
rect 24820 21360 24826 21412
rect 25222 21360 25228 21412
rect 25280 21360 25286 21412
rect 25516 21400 25544 21440
rect 25590 21428 25596 21480
rect 25648 21428 25654 21480
rect 26050 21428 26056 21480
rect 26108 21428 26114 21480
rect 26160 21400 26188 21499
rect 27062 21496 27068 21548
rect 27120 21536 27126 21548
rect 28086 21539 28144 21545
rect 28086 21536 28098 21539
rect 27120 21508 28098 21536
rect 27120 21496 27126 21508
rect 28086 21505 28098 21508
rect 28132 21505 28144 21539
rect 29270 21536 29276 21548
rect 28086 21499 28144 21505
rect 28368 21508 29276 21536
rect 28368 21477 28396 21508
rect 29270 21496 29276 21508
rect 29328 21496 29334 21548
rect 29825 21539 29883 21545
rect 29825 21505 29837 21539
rect 29871 21536 29883 21539
rect 29917 21539 29975 21545
rect 29917 21536 29929 21539
rect 29871 21508 29929 21536
rect 29871 21505 29883 21508
rect 29825 21499 29883 21505
rect 29917 21505 29929 21508
rect 29963 21536 29975 21539
rect 30006 21536 30012 21548
rect 29963 21508 30012 21536
rect 29963 21505 29975 21508
rect 29917 21499 29975 21505
rect 30006 21496 30012 21508
rect 30064 21496 30070 21548
rect 28353 21471 28411 21477
rect 28353 21437 28365 21471
rect 28399 21437 28411 21471
rect 31220 21468 31248 21564
rect 32416 21548 32444 21576
rect 32398 21496 32404 21548
rect 32456 21496 32462 21548
rect 32766 21496 32772 21548
rect 32824 21536 32830 21548
rect 33152 21545 33180 21576
rect 32861 21539 32919 21545
rect 32861 21536 32873 21539
rect 32824 21508 32873 21536
rect 32824 21496 32830 21508
rect 32861 21505 32873 21508
rect 32907 21536 32919 21539
rect 33137 21539 33195 21545
rect 32907 21508 33088 21536
rect 32907 21505 32919 21508
rect 32861 21499 32919 21505
rect 32953 21471 33011 21477
rect 32953 21468 32965 21471
rect 31220 21440 32965 21468
rect 28353 21431 28411 21437
rect 32953 21437 32965 21440
rect 32999 21437 33011 21471
rect 33060 21468 33088 21508
rect 33137 21505 33149 21539
rect 33183 21505 33195 21539
rect 33137 21499 33195 21505
rect 33229 21471 33287 21477
rect 33229 21468 33241 21471
rect 33060 21440 33241 21468
rect 32953 21431 33011 21437
rect 33229 21437 33241 21440
rect 33275 21437 33287 21471
rect 33229 21431 33287 21437
rect 33505 21471 33563 21477
rect 33505 21437 33517 21471
rect 33551 21437 33563 21471
rect 33505 21431 33563 21437
rect 25516 21372 26188 21400
rect 31294 21360 31300 21412
rect 31352 21360 31358 21412
rect 31754 21360 31760 21412
rect 31812 21400 31818 21412
rect 32585 21403 32643 21409
rect 32585 21400 32597 21403
rect 31812 21372 32597 21400
rect 31812 21360 31818 21372
rect 32585 21369 32597 21372
rect 32631 21400 32643 21403
rect 33520 21400 33548 21431
rect 33594 21428 33600 21480
rect 33652 21428 33658 21480
rect 32631 21372 33548 21400
rect 32631 21369 32643 21372
rect 32585 21363 32643 21369
rect 21499 21304 21588 21332
rect 21499 21301 21511 21304
rect 21453 21295 21511 21301
rect 22830 21292 22836 21344
rect 22888 21292 22894 21344
rect 24486 21292 24492 21344
rect 24544 21292 24550 21344
rect 25130 21292 25136 21344
rect 25188 21292 25194 21344
rect 25240 21332 25268 21360
rect 26970 21332 26976 21344
rect 25240 21304 26976 21332
rect 26970 21292 26976 21304
rect 27028 21292 27034 21344
rect 27982 21292 27988 21344
rect 28040 21332 28046 21344
rect 28445 21335 28503 21341
rect 28445 21332 28457 21335
rect 28040 21304 28457 21332
rect 28040 21292 28046 21304
rect 28445 21301 28457 21304
rect 28491 21301 28503 21335
rect 28445 21295 28503 21301
rect 32490 21292 32496 21344
rect 32548 21292 32554 21344
rect 32677 21335 32735 21341
rect 32677 21301 32689 21335
rect 32723 21332 32735 21335
rect 33502 21332 33508 21344
rect 32723 21304 33508 21332
rect 32723 21301 32735 21304
rect 32677 21295 32735 21301
rect 33502 21292 33508 21304
rect 33560 21292 33566 21344
rect 1104 21242 34868 21264
rect 1104 21190 5170 21242
rect 5222 21190 5234 21242
rect 5286 21190 5298 21242
rect 5350 21190 5362 21242
rect 5414 21190 5426 21242
rect 5478 21190 13611 21242
rect 13663 21190 13675 21242
rect 13727 21190 13739 21242
rect 13791 21190 13803 21242
rect 13855 21190 13867 21242
rect 13919 21190 22052 21242
rect 22104 21190 22116 21242
rect 22168 21190 22180 21242
rect 22232 21190 22244 21242
rect 22296 21190 22308 21242
rect 22360 21190 30493 21242
rect 30545 21190 30557 21242
rect 30609 21190 30621 21242
rect 30673 21190 30685 21242
rect 30737 21190 30749 21242
rect 30801 21190 34868 21242
rect 1104 21168 34868 21190
rect 19794 21088 19800 21140
rect 19852 21128 19858 21140
rect 20165 21131 20223 21137
rect 20165 21128 20177 21131
rect 19852 21100 20177 21128
rect 19852 21088 19858 21100
rect 20165 21097 20177 21100
rect 20211 21097 20223 21131
rect 20165 21091 20223 21097
rect 20438 21088 20444 21140
rect 20496 21088 20502 21140
rect 21910 21088 21916 21140
rect 21968 21088 21974 21140
rect 23014 21088 23020 21140
rect 23072 21128 23078 21140
rect 23661 21131 23719 21137
rect 23661 21128 23673 21131
rect 23072 21100 23673 21128
rect 23072 21088 23078 21100
rect 23661 21097 23673 21100
rect 23707 21097 23719 21131
rect 24949 21131 25007 21137
rect 24949 21128 24961 21131
rect 23661 21091 23719 21097
rect 23952 21100 24961 21128
rect 18141 20995 18199 21001
rect 18141 20961 18153 20995
rect 18187 20992 18199 20995
rect 18874 20992 18880 21004
rect 18187 20964 18880 20992
rect 18187 20961 18199 20964
rect 18141 20955 18199 20961
rect 18874 20952 18880 20964
rect 18932 20952 18938 21004
rect 20714 20992 20720 21004
rect 20272 20964 20720 20992
rect 17678 20884 17684 20936
rect 17736 20924 17742 20936
rect 17865 20927 17923 20933
rect 17865 20924 17877 20927
rect 17736 20896 17877 20924
rect 17736 20884 17742 20896
rect 17865 20893 17877 20896
rect 17911 20893 17923 20927
rect 17865 20887 17923 20893
rect 17957 20927 18015 20933
rect 17957 20893 17969 20927
rect 18003 20924 18015 20927
rect 18046 20924 18052 20936
rect 18003 20896 18052 20924
rect 18003 20893 18015 20896
rect 17957 20887 18015 20893
rect 17586 20816 17592 20868
rect 17644 20856 17650 20868
rect 17972 20856 18000 20887
rect 18046 20884 18052 20896
rect 18104 20924 18110 20936
rect 20272 20933 20300 20964
rect 20714 20952 20720 20964
rect 20772 20952 20778 21004
rect 22554 20992 22560 21004
rect 21836 20964 22560 20992
rect 21836 20933 21864 20964
rect 22554 20952 22560 20964
rect 22612 20952 22618 21004
rect 20257 20927 20315 20933
rect 18104 20896 18552 20924
rect 18104 20884 18110 20896
rect 17644 20828 18000 20856
rect 17644 20816 17650 20828
rect 18524 20800 18552 20896
rect 20257 20893 20269 20927
rect 20303 20893 20315 20927
rect 20257 20887 20315 20893
rect 20533 20927 20591 20933
rect 20533 20893 20545 20927
rect 20579 20924 20591 20927
rect 21821 20927 21879 20933
rect 21821 20924 21833 20927
rect 20579 20896 21833 20924
rect 20579 20893 20591 20896
rect 20533 20887 20591 20893
rect 21821 20893 21833 20896
rect 21867 20893 21879 20927
rect 21821 20887 21879 20893
rect 22005 20927 22063 20933
rect 22005 20893 22017 20927
rect 22051 20924 22063 20927
rect 23032 20924 23060 21088
rect 23952 21072 23980 21100
rect 24949 21097 24961 21100
rect 24995 21097 25007 21131
rect 24949 21091 25007 21097
rect 27062 21088 27068 21140
rect 27120 21088 27126 21140
rect 27338 21088 27344 21140
rect 27396 21128 27402 21140
rect 27525 21131 27583 21137
rect 27525 21128 27537 21131
rect 27396 21100 27537 21128
rect 27396 21088 27402 21100
rect 27525 21097 27537 21100
rect 27571 21097 27583 21131
rect 27525 21091 27583 21097
rect 29914 21088 29920 21140
rect 29972 21128 29978 21140
rect 30009 21131 30067 21137
rect 30009 21128 30021 21131
rect 29972 21100 30021 21128
rect 29972 21088 29978 21100
rect 30009 21097 30021 21100
rect 30055 21097 30067 21131
rect 30009 21091 30067 21097
rect 30392 21100 31754 21128
rect 23934 21020 23940 21072
rect 23992 21020 23998 21072
rect 26050 21060 26056 21072
rect 24228 21032 25084 21060
rect 24026 20992 24032 21004
rect 23861 20964 24032 20992
rect 23861 20933 23889 20964
rect 24026 20952 24032 20964
rect 24084 20952 24090 21004
rect 24121 20995 24179 21001
rect 24121 20961 24133 20995
rect 24167 20961 24179 20995
rect 24121 20955 24179 20961
rect 22051 20896 23060 20924
rect 23845 20927 23903 20933
rect 22051 20893 22063 20896
rect 22005 20887 22063 20893
rect 23845 20893 23857 20927
rect 23891 20893 23903 20927
rect 23845 20887 23903 20893
rect 23934 20884 23940 20936
rect 23992 20884 23998 20936
rect 24136 20856 24164 20955
rect 24228 20933 24256 21032
rect 24302 20952 24308 21004
rect 24360 20992 24366 21004
rect 25056 21001 25084 21032
rect 25231 21032 26056 21060
rect 25041 20995 25099 21001
rect 24360 20964 24808 20992
rect 24360 20952 24366 20964
rect 24780 20933 24808 20964
rect 25041 20961 25053 20995
rect 25087 20992 25099 20995
rect 25130 20992 25136 21004
rect 25087 20964 25136 20992
rect 25087 20961 25099 20964
rect 25041 20955 25099 20961
rect 25130 20952 25136 20964
rect 25188 20952 25194 21004
rect 24213 20927 24271 20933
rect 24213 20893 24225 20927
rect 24259 20893 24271 20927
rect 24673 20927 24731 20933
rect 24673 20921 24685 20927
rect 24213 20887 24271 20893
rect 24670 20893 24685 20921
rect 24719 20893 24731 20927
rect 24670 20887 24731 20893
rect 24765 20927 24823 20933
rect 24765 20893 24777 20927
rect 24811 20924 24823 20927
rect 25231 20924 25259 21032
rect 26050 21020 26056 21032
rect 26108 21020 26114 21072
rect 27706 21020 27712 21072
rect 27764 21060 27770 21072
rect 27985 21063 28043 21069
rect 27985 21060 27997 21063
rect 27764 21032 27997 21060
rect 27764 21020 27770 21032
rect 27985 21029 27997 21032
rect 28031 21029 28043 21063
rect 27985 21023 28043 21029
rect 27157 20995 27215 21001
rect 27157 20992 27169 20995
rect 26068 20964 26556 20992
rect 24811 20896 25259 20924
rect 24811 20893 24823 20896
rect 24765 20887 24823 20893
rect 24670 20856 24698 20887
rect 25314 20884 25320 20936
rect 25372 20884 25378 20936
rect 25409 20927 25467 20933
rect 25409 20893 25421 20927
rect 25455 20893 25467 20927
rect 25409 20887 25467 20893
rect 25133 20859 25191 20865
rect 25133 20856 25145 20859
rect 22066 20828 24072 20856
rect 24136 20828 25145 20856
rect 18141 20791 18199 20797
rect 18141 20757 18153 20791
rect 18187 20788 18199 20791
rect 18230 20788 18236 20800
rect 18187 20760 18236 20788
rect 18187 20757 18199 20760
rect 18141 20751 18199 20757
rect 18230 20748 18236 20760
rect 18288 20748 18294 20800
rect 18506 20748 18512 20800
rect 18564 20748 18570 20800
rect 21174 20748 21180 20800
rect 21232 20788 21238 20800
rect 21542 20788 21548 20800
rect 21232 20760 21548 20788
rect 21232 20748 21238 20760
rect 21542 20748 21548 20760
rect 21600 20788 21606 20800
rect 22066 20788 22094 20828
rect 21600 20760 22094 20788
rect 24044 20788 24072 20828
rect 25133 20825 25145 20828
rect 25179 20825 25191 20859
rect 25133 20819 25191 20825
rect 24489 20791 24547 20797
rect 24489 20788 24501 20791
rect 24044 20760 24501 20788
rect 21600 20748 21606 20760
rect 24489 20757 24501 20760
rect 24535 20757 24547 20791
rect 24489 20751 24547 20757
rect 24578 20748 24584 20800
rect 24636 20788 24642 20800
rect 25424 20788 25452 20887
rect 25590 20884 25596 20936
rect 25648 20924 25654 20936
rect 26068 20924 26096 20964
rect 25648 20896 26096 20924
rect 26421 20927 26479 20933
rect 25648 20884 25654 20896
rect 26421 20893 26433 20927
rect 26467 20893 26479 20927
rect 26421 20887 26479 20893
rect 24636 20760 25452 20788
rect 26436 20788 26464 20887
rect 26528 20856 26556 20964
rect 26712 20964 27169 20992
rect 26602 20884 26608 20936
rect 26660 20884 26666 20936
rect 26712 20933 26740 20964
rect 27157 20961 27169 20964
rect 27203 20961 27215 20995
rect 27157 20955 27215 20961
rect 30006 20952 30012 21004
rect 30064 20992 30070 21004
rect 30392 21001 30420 21100
rect 31726 21060 31754 21100
rect 31938 21088 31944 21140
rect 31996 21128 32002 21140
rect 32398 21128 32404 21140
rect 31996 21100 32404 21128
rect 31996 21088 32002 21100
rect 32398 21088 32404 21100
rect 32456 21088 32462 21140
rect 32766 21128 32772 21140
rect 32508 21100 32772 21128
rect 32508 21060 32536 21100
rect 32766 21088 32772 21100
rect 32824 21128 32830 21140
rect 33873 21131 33931 21137
rect 33873 21128 33885 21131
rect 32824 21100 33885 21128
rect 32824 21088 32830 21100
rect 33873 21097 33885 21100
rect 33919 21097 33931 21131
rect 33873 21091 33931 21097
rect 31726 21032 32536 21060
rect 30377 20995 30435 21001
rect 30064 20964 30328 20992
rect 30064 20952 30070 20964
rect 26697 20927 26755 20933
rect 26697 20893 26709 20927
rect 26743 20893 26755 20927
rect 26697 20887 26755 20893
rect 26786 20884 26792 20936
rect 26844 20884 26850 20936
rect 26970 20884 26976 20936
rect 27028 20924 27034 20936
rect 27430 20924 27436 20936
rect 27028 20896 27436 20924
rect 27028 20884 27034 20896
rect 27430 20884 27436 20896
rect 27488 20884 27494 20936
rect 27617 20927 27675 20933
rect 27617 20893 27629 20927
rect 27663 20924 27675 20927
rect 27798 20924 27804 20936
rect 27663 20896 27804 20924
rect 27663 20893 27675 20896
rect 27617 20887 27675 20893
rect 27798 20884 27804 20896
rect 27856 20884 27862 20936
rect 27893 20927 27951 20933
rect 27893 20893 27905 20927
rect 27939 20924 27951 20927
rect 27982 20924 27988 20936
rect 27939 20896 27988 20924
rect 27939 20893 27951 20896
rect 27893 20887 27951 20893
rect 27982 20884 27988 20896
rect 28040 20884 28046 20936
rect 29270 20884 29276 20936
rect 29328 20924 29334 20936
rect 29365 20927 29423 20933
rect 29365 20924 29377 20927
rect 29328 20896 29377 20924
rect 29328 20884 29334 20896
rect 29365 20893 29377 20896
rect 29411 20893 29423 20927
rect 29365 20887 29423 20893
rect 30193 20927 30251 20933
rect 30193 20893 30205 20927
rect 30239 20893 30251 20927
rect 30300 20924 30328 20964
rect 30377 20961 30389 20995
rect 30423 20961 30435 20995
rect 30377 20955 30435 20961
rect 30834 20933 30840 20936
rect 30561 20927 30619 20933
rect 30561 20924 30573 20927
rect 30300 20896 30573 20924
rect 30193 20887 30251 20893
rect 30561 20893 30573 20896
rect 30607 20893 30619 20927
rect 30828 20924 30840 20933
rect 30795 20896 30840 20924
rect 30561 20887 30619 20893
rect 30828 20887 30840 20896
rect 26528 20828 28856 20856
rect 26694 20788 26700 20800
rect 26436 20760 26700 20788
rect 24636 20748 24642 20760
rect 26694 20748 26700 20760
rect 26752 20788 26758 20800
rect 28718 20788 28724 20800
rect 26752 20760 28724 20788
rect 26752 20748 26758 20760
rect 28718 20748 28724 20760
rect 28776 20748 28782 20800
rect 28828 20788 28856 20828
rect 28994 20816 29000 20868
rect 29052 20856 29058 20868
rect 29098 20859 29156 20865
rect 29098 20856 29110 20859
rect 29052 20828 29110 20856
rect 29052 20816 29058 20828
rect 29098 20825 29110 20828
rect 29144 20825 29156 20859
rect 30208 20856 30236 20887
rect 30374 20856 30380 20868
rect 30208 20828 30380 20856
rect 29098 20819 29156 20825
rect 30374 20816 30380 20828
rect 30432 20816 30438 20868
rect 30576 20856 30604 20887
rect 30834 20884 30840 20887
rect 30892 20884 30898 20936
rect 32493 20927 32551 20933
rect 32493 20924 32505 20927
rect 31726 20896 32505 20924
rect 30926 20856 30932 20868
rect 30576 20828 30932 20856
rect 30926 20816 30932 20828
rect 30984 20856 30990 20868
rect 31726 20856 31754 20896
rect 32493 20893 32505 20896
rect 32539 20893 32551 20927
rect 32493 20887 32551 20893
rect 30984 20828 31754 20856
rect 32760 20859 32818 20865
rect 30984 20816 30990 20828
rect 32760 20825 32772 20859
rect 32806 20856 32818 20859
rect 33318 20856 33324 20868
rect 32806 20828 33324 20856
rect 32806 20825 32818 20828
rect 32760 20819 32818 20825
rect 33318 20816 33324 20828
rect 33376 20816 33382 20868
rect 31938 20788 31944 20800
rect 28828 20760 31944 20788
rect 31938 20748 31944 20760
rect 31996 20748 32002 20800
rect 1104 20698 35027 20720
rect 1104 20646 9390 20698
rect 9442 20646 9454 20698
rect 9506 20646 9518 20698
rect 9570 20646 9582 20698
rect 9634 20646 9646 20698
rect 9698 20646 17831 20698
rect 17883 20646 17895 20698
rect 17947 20646 17959 20698
rect 18011 20646 18023 20698
rect 18075 20646 18087 20698
rect 18139 20646 26272 20698
rect 26324 20646 26336 20698
rect 26388 20646 26400 20698
rect 26452 20646 26464 20698
rect 26516 20646 26528 20698
rect 26580 20646 34713 20698
rect 34765 20646 34777 20698
rect 34829 20646 34841 20698
rect 34893 20646 34905 20698
rect 34957 20646 34969 20698
rect 35021 20646 35027 20698
rect 1104 20624 35027 20646
rect 17126 20544 17132 20596
rect 17184 20584 17190 20596
rect 17770 20584 17776 20596
rect 17184 20556 17776 20584
rect 17184 20544 17190 20556
rect 17770 20544 17776 20556
rect 17828 20544 17834 20596
rect 18230 20544 18236 20596
rect 18288 20544 18294 20596
rect 19610 20544 19616 20596
rect 19668 20544 19674 20596
rect 19702 20544 19708 20596
rect 19760 20584 19766 20596
rect 20257 20587 20315 20593
rect 20257 20584 20269 20587
rect 19760 20556 20269 20584
rect 19760 20544 19766 20556
rect 18248 20516 18276 20544
rect 17420 20488 18276 20516
rect 19628 20516 19656 20544
rect 19797 20519 19855 20525
rect 19797 20516 19809 20519
rect 19628 20488 19809 20516
rect 17420 20457 17448 20488
rect 19797 20485 19809 20488
rect 19843 20485 19855 20519
rect 19797 20479 19855 20485
rect 17221 20451 17279 20457
rect 17221 20417 17233 20451
rect 17267 20417 17279 20451
rect 17221 20411 17279 20417
rect 17405 20451 17463 20457
rect 17405 20417 17417 20451
rect 17451 20417 17463 20451
rect 17405 20411 17463 20417
rect 17236 20312 17264 20411
rect 17586 20408 17592 20460
rect 17644 20448 17650 20460
rect 17681 20451 17739 20457
rect 17681 20448 17693 20451
rect 17644 20420 17693 20448
rect 17644 20408 17650 20420
rect 17681 20417 17693 20420
rect 17727 20417 17739 20451
rect 18213 20451 18271 20457
rect 18213 20448 18225 20451
rect 17681 20411 17739 20417
rect 17788 20420 18225 20448
rect 17313 20383 17371 20389
rect 17313 20349 17325 20383
rect 17359 20380 17371 20383
rect 17788 20380 17816 20420
rect 18213 20417 18225 20420
rect 18259 20417 18271 20451
rect 19567 20451 19625 20457
rect 19567 20448 19579 20451
rect 18213 20411 18271 20417
rect 19352 20420 19579 20448
rect 17359 20352 17816 20380
rect 17865 20383 17923 20389
rect 17359 20349 17371 20352
rect 17313 20343 17371 20349
rect 17865 20349 17877 20383
rect 17911 20349 17923 20383
rect 17865 20343 17923 20349
rect 17236 20284 17540 20312
rect 17512 20253 17540 20284
rect 17678 20272 17684 20324
rect 17736 20312 17742 20324
rect 17880 20312 17908 20343
rect 17954 20340 17960 20392
rect 18012 20340 18018 20392
rect 17736 20284 17908 20312
rect 17736 20272 17742 20284
rect 19352 20256 19380 20420
rect 19567 20417 19579 20420
rect 19613 20417 19625 20451
rect 19567 20411 19625 20417
rect 19702 20408 19708 20460
rect 19760 20408 19766 20460
rect 19996 20457 20024 20556
rect 20257 20553 20269 20556
rect 20303 20553 20315 20587
rect 23014 20584 23020 20596
rect 20257 20547 20315 20553
rect 22388 20556 23020 20584
rect 22388 20525 22416 20556
rect 23014 20544 23020 20556
rect 23072 20544 23078 20596
rect 26602 20544 26608 20596
rect 26660 20584 26666 20596
rect 27249 20587 27307 20593
rect 27249 20584 27261 20587
rect 26660 20556 27261 20584
rect 26660 20544 26666 20556
rect 27249 20553 27261 20556
rect 27295 20553 27307 20587
rect 27249 20547 27307 20553
rect 27706 20544 27712 20596
rect 27764 20544 27770 20596
rect 27798 20544 27804 20596
rect 27856 20544 27862 20596
rect 28721 20587 28779 20593
rect 28721 20553 28733 20587
rect 28767 20584 28779 20587
rect 28994 20584 29000 20596
rect 28767 20556 29000 20584
rect 28767 20553 28779 20556
rect 28721 20547 28779 20553
rect 28994 20544 29000 20556
rect 29052 20544 29058 20596
rect 29104 20556 31754 20584
rect 22373 20519 22431 20525
rect 22373 20485 22385 20519
rect 22419 20485 22431 20519
rect 22373 20479 22431 20485
rect 22462 20476 22468 20528
rect 22520 20516 22526 20528
rect 22520 20488 23888 20516
rect 22520 20476 22526 20488
rect 19980 20451 20038 20457
rect 19980 20417 19992 20451
rect 20026 20417 20038 20451
rect 19980 20411 20038 20417
rect 20073 20451 20131 20457
rect 20073 20417 20085 20451
rect 20119 20448 20131 20451
rect 20254 20448 20260 20460
rect 20119 20420 20260 20448
rect 20119 20417 20131 20420
rect 20073 20411 20131 20417
rect 20254 20408 20260 20420
rect 20312 20408 20318 20460
rect 20349 20451 20407 20457
rect 20349 20417 20361 20451
rect 20395 20448 20407 20451
rect 22557 20451 22615 20457
rect 22557 20448 22569 20451
rect 20395 20420 22569 20448
rect 20395 20417 20407 20420
rect 20349 20411 20407 20417
rect 22557 20417 22569 20420
rect 22603 20448 22615 20451
rect 22646 20448 22652 20460
rect 22603 20420 22652 20448
rect 22603 20417 22615 20420
rect 22557 20411 22615 20417
rect 22646 20408 22652 20420
rect 22704 20448 22710 20460
rect 23198 20448 23204 20460
rect 22704 20420 23204 20448
rect 22704 20408 22710 20420
rect 23198 20408 23204 20420
rect 23256 20448 23262 20460
rect 23385 20451 23443 20457
rect 23385 20448 23397 20451
rect 23256 20420 23397 20448
rect 23256 20408 23262 20420
rect 23385 20417 23397 20420
rect 23431 20417 23443 20451
rect 23385 20411 23443 20417
rect 23474 20408 23480 20460
rect 23532 20408 23538 20460
rect 23569 20451 23627 20457
rect 23569 20417 23581 20451
rect 23615 20417 23627 20451
rect 23569 20411 23627 20417
rect 23492 20312 23520 20408
rect 23584 20380 23612 20411
rect 23658 20408 23664 20460
rect 23716 20448 23722 20460
rect 23860 20457 23888 20488
rect 26878 20476 26884 20528
rect 26936 20516 26942 20528
rect 27816 20516 27844 20544
rect 29104 20516 29132 20556
rect 26936 20488 27752 20516
rect 27816 20488 28028 20516
rect 26936 20476 26942 20488
rect 23753 20451 23811 20457
rect 23753 20448 23765 20451
rect 23716 20420 23765 20448
rect 23716 20408 23722 20420
rect 23753 20417 23765 20420
rect 23799 20417 23811 20451
rect 23753 20411 23811 20417
rect 23845 20451 23903 20457
rect 23845 20417 23857 20451
rect 23891 20417 23903 20451
rect 23845 20411 23903 20417
rect 24029 20451 24087 20457
rect 24029 20417 24041 20451
rect 24075 20417 24087 20451
rect 24029 20411 24087 20417
rect 23937 20383 23995 20389
rect 23937 20380 23949 20383
rect 23584 20352 23949 20380
rect 23937 20349 23949 20352
rect 23983 20349 23995 20383
rect 23937 20343 23995 20349
rect 24044 20312 24072 20411
rect 26142 20408 26148 20460
rect 26200 20408 26206 20460
rect 26329 20451 26387 20457
rect 26329 20417 26341 20451
rect 26375 20448 26387 20451
rect 26605 20451 26663 20457
rect 26605 20448 26617 20451
rect 26375 20420 26617 20448
rect 26375 20417 26387 20420
rect 26329 20411 26387 20417
rect 26605 20417 26617 20420
rect 26651 20417 26663 20451
rect 26605 20411 26663 20417
rect 27154 20408 27160 20460
rect 27212 20408 27218 20460
rect 27430 20408 27436 20460
rect 27488 20408 27494 20460
rect 25961 20383 26019 20389
rect 25961 20349 25973 20383
rect 26007 20349 26019 20383
rect 25961 20343 26019 20349
rect 27525 20383 27583 20389
rect 27525 20349 27537 20383
rect 27571 20349 27583 20383
rect 27724 20380 27752 20488
rect 27890 20408 27896 20460
rect 27948 20408 27954 20460
rect 28000 20457 28028 20488
rect 28092 20488 29132 20516
rect 27985 20451 28043 20457
rect 27985 20417 27997 20451
rect 28031 20417 28043 20451
rect 27985 20411 28043 20417
rect 28092 20380 28120 20488
rect 30558 20476 30564 20528
rect 30616 20516 30622 20528
rect 31726 20516 31754 20556
rect 32490 20544 32496 20596
rect 32548 20584 32554 20596
rect 32585 20587 32643 20593
rect 32585 20584 32597 20587
rect 32548 20556 32597 20584
rect 32548 20544 32554 20556
rect 32585 20553 32597 20556
rect 32631 20553 32643 20587
rect 32585 20547 32643 20553
rect 33318 20544 33324 20596
rect 33376 20544 33382 20596
rect 32858 20516 32864 20528
rect 30616 20488 31156 20516
rect 31726 20488 32864 20516
rect 30616 20476 30622 20488
rect 28166 20408 28172 20460
rect 28224 20408 28230 20460
rect 31128 20457 31156 20488
rect 32858 20476 32864 20488
rect 32916 20476 32922 20528
rect 28353 20451 28411 20457
rect 28353 20417 28365 20451
rect 28399 20448 28411 20451
rect 28537 20451 28595 20457
rect 28537 20448 28549 20451
rect 28399 20420 28549 20448
rect 28399 20417 28411 20420
rect 28353 20411 28411 20417
rect 28537 20417 28549 20420
rect 28583 20417 28595 20451
rect 28537 20411 28595 20417
rect 31021 20451 31079 20457
rect 31021 20417 31033 20451
rect 31067 20417 31079 20451
rect 31021 20411 31079 20417
rect 31113 20451 31171 20457
rect 31113 20417 31125 20451
rect 31159 20448 31171 20451
rect 31202 20448 31208 20460
rect 31159 20420 31208 20448
rect 31159 20417 31171 20420
rect 31113 20411 31171 20417
rect 27724 20352 28120 20380
rect 31036 20380 31064 20411
rect 31202 20408 31208 20420
rect 31260 20408 31266 20460
rect 31297 20451 31355 20457
rect 31297 20417 31309 20451
rect 31343 20448 31355 20451
rect 31573 20451 31631 20457
rect 31573 20448 31585 20451
rect 31343 20420 31585 20448
rect 31343 20417 31355 20420
rect 31297 20411 31355 20417
rect 31573 20417 31585 20420
rect 31619 20417 31631 20451
rect 31573 20411 31631 20417
rect 31938 20408 31944 20460
rect 31996 20448 32002 20460
rect 32125 20451 32183 20457
rect 32125 20448 32137 20451
rect 31996 20420 32137 20448
rect 31996 20408 32002 20420
rect 32125 20417 32137 20420
rect 32171 20417 32183 20451
rect 32125 20411 32183 20417
rect 32398 20408 32404 20460
rect 32456 20408 32462 20460
rect 33226 20408 33232 20460
rect 33284 20408 33290 20460
rect 33502 20408 33508 20460
rect 33560 20408 33566 20460
rect 31036 20352 31754 20380
rect 27525 20343 27583 20349
rect 23492 20284 24072 20312
rect 25976 20312 26004 20343
rect 27540 20312 27568 20343
rect 27982 20312 27988 20324
rect 25976 20284 27988 20312
rect 27982 20272 27988 20284
rect 28040 20272 28046 20324
rect 17497 20247 17555 20253
rect 17497 20213 17509 20247
rect 17543 20244 17555 20247
rect 18138 20244 18144 20256
rect 17543 20216 18144 20244
rect 17543 20213 17555 20216
rect 17497 20207 17555 20213
rect 18138 20204 18144 20216
rect 18196 20204 18202 20256
rect 19334 20204 19340 20256
rect 19392 20204 19398 20256
rect 19426 20204 19432 20256
rect 19484 20204 19490 20256
rect 22738 20204 22744 20256
rect 22796 20204 22802 20256
rect 23106 20204 23112 20256
rect 23164 20204 23170 20256
rect 26418 20204 26424 20256
rect 26476 20204 26482 20256
rect 26970 20204 26976 20256
rect 27028 20204 27034 20256
rect 31386 20204 31392 20256
rect 31444 20204 31450 20256
rect 31726 20244 31754 20352
rect 32214 20340 32220 20392
rect 32272 20340 32278 20392
rect 32306 20272 32312 20324
rect 32364 20312 32370 20324
rect 32677 20315 32735 20321
rect 32677 20312 32689 20315
rect 32364 20284 32689 20312
rect 32364 20272 32370 20284
rect 32677 20281 32689 20284
rect 32723 20281 32735 20315
rect 32677 20275 32735 20281
rect 32401 20247 32459 20253
rect 32401 20244 32413 20247
rect 31726 20216 32413 20244
rect 32401 20213 32413 20216
rect 32447 20244 32459 20247
rect 32582 20244 32588 20256
rect 32447 20216 32588 20244
rect 32447 20213 32459 20216
rect 32401 20207 32459 20213
rect 32582 20204 32588 20216
rect 32640 20204 32646 20256
rect 33042 20204 33048 20256
rect 33100 20204 33106 20256
rect 1104 20154 34868 20176
rect 1104 20102 5170 20154
rect 5222 20102 5234 20154
rect 5286 20102 5298 20154
rect 5350 20102 5362 20154
rect 5414 20102 5426 20154
rect 5478 20102 13611 20154
rect 13663 20102 13675 20154
rect 13727 20102 13739 20154
rect 13791 20102 13803 20154
rect 13855 20102 13867 20154
rect 13919 20102 22052 20154
rect 22104 20102 22116 20154
rect 22168 20102 22180 20154
rect 22232 20102 22244 20154
rect 22296 20102 22308 20154
rect 22360 20102 30493 20154
rect 30545 20102 30557 20154
rect 30609 20102 30621 20154
rect 30673 20102 30685 20154
rect 30737 20102 30749 20154
rect 30801 20102 34868 20154
rect 1104 20080 34868 20102
rect 17678 20000 17684 20052
rect 17736 20000 17742 20052
rect 18138 20000 18144 20052
rect 18196 20000 18202 20052
rect 18509 20043 18567 20049
rect 18509 20009 18521 20043
rect 18555 20040 18567 20043
rect 19334 20040 19340 20052
rect 18555 20012 19340 20040
rect 18555 20009 18567 20012
rect 18509 20003 18567 20009
rect 17696 19972 17724 20000
rect 18524 19972 18552 20003
rect 19334 20000 19340 20012
rect 19392 20000 19398 20052
rect 19702 20000 19708 20052
rect 19760 20040 19766 20052
rect 19981 20043 20039 20049
rect 19981 20040 19993 20043
rect 19760 20012 19993 20040
rect 19760 20000 19766 20012
rect 19981 20009 19993 20012
rect 20027 20009 20039 20043
rect 19981 20003 20039 20009
rect 22373 20043 22431 20049
rect 22373 20009 22385 20043
rect 22419 20040 22431 20043
rect 22462 20040 22468 20052
rect 22419 20012 22468 20040
rect 22419 20009 22431 20012
rect 22373 20003 22431 20009
rect 22462 20000 22468 20012
rect 22520 20000 22526 20052
rect 22738 20000 22744 20052
rect 22796 20000 22802 20052
rect 23198 20000 23204 20052
rect 23256 20040 23262 20052
rect 24213 20043 24271 20049
rect 24213 20040 24225 20043
rect 23256 20012 24225 20040
rect 23256 20000 23262 20012
rect 24213 20009 24225 20012
rect 24259 20009 24271 20043
rect 24213 20003 24271 20009
rect 26418 20000 26424 20052
rect 26476 20000 26482 20052
rect 26786 20000 26792 20052
rect 26844 20000 26850 20052
rect 27798 20000 27804 20052
rect 27856 20040 27862 20052
rect 28261 20043 28319 20049
rect 28261 20040 28273 20043
rect 27856 20012 28273 20040
rect 27856 20000 27862 20012
rect 28261 20009 28273 20012
rect 28307 20009 28319 20043
rect 28261 20003 28319 20009
rect 29178 20000 29184 20052
rect 29236 20040 29242 20052
rect 29546 20040 29552 20052
rect 29236 20012 29552 20040
rect 29236 20000 29242 20012
rect 29546 20000 29552 20012
rect 29604 20000 29610 20052
rect 31202 20000 31208 20052
rect 31260 20040 31266 20052
rect 31260 20012 33364 20040
rect 31260 20000 31266 20012
rect 17696 19944 18552 19972
rect 18233 19907 18291 19913
rect 18233 19904 18245 19907
rect 17880 19876 18245 19904
rect 934 19796 940 19848
rect 992 19836 998 19848
rect 1397 19839 1455 19845
rect 1397 19836 1409 19839
rect 992 19808 1409 19836
rect 992 19796 998 19808
rect 1397 19805 1409 19808
rect 1443 19805 1455 19839
rect 1397 19799 1455 19805
rect 17678 19796 17684 19848
rect 17736 19796 17742 19848
rect 17436 19771 17494 19777
rect 17436 19737 17448 19771
rect 17482 19768 17494 19771
rect 17773 19771 17831 19777
rect 17773 19768 17785 19771
rect 17482 19740 17785 19768
rect 17482 19737 17494 19740
rect 17436 19731 17494 19737
rect 17773 19737 17785 19740
rect 17819 19737 17831 19771
rect 17773 19731 17831 19737
rect 16301 19703 16359 19709
rect 16301 19669 16313 19703
rect 16347 19700 16359 19703
rect 17880 19700 17908 19876
rect 18233 19873 18245 19876
rect 18279 19873 18291 19907
rect 18233 19867 18291 19873
rect 17957 19839 18015 19845
rect 17957 19805 17969 19839
rect 18003 19805 18015 19839
rect 18248 19836 18276 19867
rect 18248 19808 18736 19836
rect 17957 19799 18015 19805
rect 17972 19768 18000 19799
rect 18708 19780 18736 19808
rect 18506 19777 18512 19780
rect 18493 19771 18512 19777
rect 17972 19740 18276 19768
rect 18248 19712 18276 19740
rect 18493 19737 18505 19771
rect 18493 19731 18512 19737
rect 18506 19728 18512 19731
rect 18564 19728 18570 19780
rect 18690 19728 18696 19780
rect 18748 19728 18754 19780
rect 19352 19768 19380 20000
rect 19429 19839 19487 19845
rect 19429 19805 19441 19839
rect 19475 19836 19487 19839
rect 19720 19836 19748 20000
rect 19794 19932 19800 19984
rect 19852 19972 19858 19984
rect 21910 19972 21916 19984
rect 19852 19944 21916 19972
rect 19852 19932 19858 19944
rect 21910 19932 21916 19944
rect 21968 19932 21974 19984
rect 21545 19907 21603 19913
rect 21545 19873 21557 19907
rect 21591 19873 21603 19907
rect 21545 19867 21603 19873
rect 21729 19907 21787 19913
rect 21729 19873 21741 19907
rect 21775 19904 21787 19907
rect 22186 19904 22192 19916
rect 21775 19876 22192 19904
rect 21775 19873 21787 19876
rect 21729 19867 21787 19873
rect 19475 19808 19748 19836
rect 19475 19805 19487 19808
rect 19429 19799 19487 19805
rect 20070 19796 20076 19848
rect 20128 19796 20134 19848
rect 21174 19796 21180 19848
rect 21232 19796 21238 19848
rect 21453 19839 21511 19845
rect 21453 19805 21465 19839
rect 21499 19805 21511 19839
rect 21453 19799 21511 19805
rect 19613 19771 19671 19777
rect 19613 19768 19625 19771
rect 19352 19740 19625 19768
rect 19613 19737 19625 19740
rect 19659 19737 19671 19771
rect 19613 19731 19671 19737
rect 16347 19672 17908 19700
rect 16347 19669 16359 19672
rect 16301 19663 16359 19669
rect 18230 19660 18236 19712
rect 18288 19660 18294 19712
rect 18322 19660 18328 19712
rect 18380 19660 18386 19712
rect 19242 19660 19248 19712
rect 19300 19660 19306 19712
rect 20714 19660 20720 19712
rect 20772 19700 20778 19712
rect 20993 19703 21051 19709
rect 20993 19700 21005 19703
rect 20772 19672 21005 19700
rect 20772 19660 20778 19672
rect 20993 19669 21005 19672
rect 21039 19669 21051 19703
rect 20993 19663 21051 19669
rect 21358 19660 21364 19712
rect 21416 19660 21422 19712
rect 21468 19700 21496 19799
rect 21560 19768 21588 19867
rect 22186 19864 22192 19876
rect 22244 19904 22250 19916
rect 22649 19907 22707 19913
rect 22649 19904 22661 19907
rect 22244 19876 22661 19904
rect 22244 19864 22250 19876
rect 22649 19873 22661 19876
rect 22695 19873 22707 19907
rect 22649 19867 22707 19873
rect 21821 19839 21879 19845
rect 21821 19805 21833 19839
rect 21867 19836 21879 19839
rect 22097 19839 22155 19845
rect 22097 19836 22109 19839
rect 21867 19808 22109 19836
rect 21867 19805 21879 19808
rect 21821 19799 21879 19805
rect 22097 19805 22109 19808
rect 22143 19836 22155 19839
rect 22370 19836 22376 19848
rect 22143 19808 22376 19836
rect 22143 19805 22155 19808
rect 22097 19799 22155 19805
rect 22370 19796 22376 19808
rect 22428 19796 22434 19848
rect 22756 19845 22784 20000
rect 22830 19864 22836 19916
rect 22888 19864 22894 19916
rect 23106 19845 23112 19848
rect 22557 19839 22615 19845
rect 22557 19805 22569 19839
rect 22603 19805 22615 19839
rect 22557 19799 22615 19805
rect 22741 19839 22799 19845
rect 22741 19805 22753 19839
rect 22787 19805 22799 19839
rect 23100 19836 23112 19845
rect 23067 19808 23112 19836
rect 22741 19799 22799 19805
rect 23100 19799 23112 19808
rect 22572 19768 22600 19799
rect 23106 19796 23112 19799
rect 23164 19796 23170 19848
rect 25409 19839 25467 19845
rect 25409 19805 25421 19839
rect 25455 19805 25467 19839
rect 25409 19799 25467 19805
rect 25676 19839 25734 19845
rect 25676 19805 25688 19839
rect 25722 19836 25734 19839
rect 26436 19836 26464 20000
rect 32398 19932 32404 19984
rect 32456 19972 32462 19984
rect 32456 19944 32481 19972
rect 32456 19932 32462 19944
rect 30926 19864 30932 19916
rect 30984 19904 30990 19916
rect 31021 19907 31079 19913
rect 31021 19904 31033 19907
rect 30984 19876 31033 19904
rect 30984 19864 30990 19876
rect 31021 19873 31033 19876
rect 31067 19873 31079 19907
rect 31021 19867 31079 19873
rect 32122 19864 32128 19916
rect 32180 19904 32186 19916
rect 32416 19904 32444 19932
rect 32493 19907 32551 19913
rect 32493 19904 32505 19907
rect 32180 19876 32505 19904
rect 32180 19864 32186 19876
rect 32493 19873 32505 19876
rect 32539 19873 32551 19907
rect 32493 19867 32551 19873
rect 25722 19808 26464 19836
rect 26881 19839 26939 19845
rect 25722 19805 25734 19808
rect 25676 19799 25734 19805
rect 26881 19805 26893 19839
rect 26927 19805 26939 19839
rect 26881 19799 26939 19805
rect 25424 19768 25452 19799
rect 25866 19768 25872 19780
rect 21560 19740 22968 19768
rect 25424 19740 25872 19768
rect 22940 19712 22968 19740
rect 25866 19728 25872 19740
rect 25924 19768 25930 19780
rect 26896 19768 26924 19799
rect 26970 19796 26976 19848
rect 27028 19836 27034 19848
rect 27137 19839 27195 19845
rect 27137 19836 27149 19839
rect 27028 19808 27149 19836
rect 27028 19796 27034 19808
rect 27137 19805 27149 19808
rect 27183 19805 27195 19839
rect 27137 19799 27195 19805
rect 32214 19796 32220 19848
rect 32272 19836 32278 19848
rect 32769 19839 32827 19845
rect 32769 19836 32781 19839
rect 32272 19808 32781 19836
rect 32272 19796 32278 19808
rect 32769 19805 32781 19808
rect 32815 19836 32827 19839
rect 33134 19836 33140 19848
rect 32815 19808 33140 19836
rect 32815 19805 32827 19808
rect 32769 19799 32827 19805
rect 33134 19796 33140 19808
rect 33192 19796 33198 19848
rect 33336 19845 33364 20012
rect 33502 20000 33508 20052
rect 33560 20000 33566 20052
rect 33321 19839 33379 19845
rect 33321 19805 33333 19839
rect 33367 19805 33379 19839
rect 33321 19799 33379 19805
rect 33594 19796 33600 19848
rect 33652 19796 33658 19848
rect 25924 19740 26924 19768
rect 25924 19728 25930 19740
rect 29362 19728 29368 19780
rect 29420 19768 29426 19780
rect 30662 19771 30720 19777
rect 30662 19768 30674 19771
rect 29420 19740 30674 19768
rect 29420 19728 29426 19740
rect 30662 19737 30674 19740
rect 30708 19737 30720 19771
rect 30662 19731 30720 19737
rect 31288 19771 31346 19777
rect 31288 19737 31300 19771
rect 31334 19768 31346 19771
rect 31386 19768 31392 19780
rect 31334 19740 31392 19768
rect 31334 19737 31346 19740
rect 31288 19731 31346 19737
rect 31386 19728 31392 19740
rect 31444 19728 31450 19780
rect 33045 19771 33103 19777
rect 33045 19737 33057 19771
rect 33091 19768 33103 19771
rect 33612 19768 33640 19796
rect 33091 19740 33640 19768
rect 33091 19737 33103 19740
rect 33045 19731 33103 19737
rect 21545 19703 21603 19709
rect 21545 19700 21557 19703
rect 21468 19672 21557 19700
rect 21545 19669 21557 19672
rect 21591 19700 21603 19703
rect 21726 19700 21732 19712
rect 21591 19672 21732 19700
rect 21591 19669 21603 19672
rect 21545 19663 21603 19669
rect 21726 19660 21732 19672
rect 21784 19660 21790 19712
rect 22922 19660 22928 19712
rect 22980 19660 22986 19712
rect 32582 19660 32588 19712
rect 32640 19700 32646 19712
rect 32677 19703 32735 19709
rect 32677 19700 32689 19703
rect 32640 19672 32689 19700
rect 32640 19660 32646 19672
rect 32677 19669 32689 19672
rect 32723 19669 32735 19703
rect 32677 19663 32735 19669
rect 32858 19660 32864 19712
rect 32916 19660 32922 19712
rect 1104 19610 35027 19632
rect 1104 19558 9390 19610
rect 9442 19558 9454 19610
rect 9506 19558 9518 19610
rect 9570 19558 9582 19610
rect 9634 19558 9646 19610
rect 9698 19558 17831 19610
rect 17883 19558 17895 19610
rect 17947 19558 17959 19610
rect 18011 19558 18023 19610
rect 18075 19558 18087 19610
rect 18139 19558 26272 19610
rect 26324 19558 26336 19610
rect 26388 19558 26400 19610
rect 26452 19558 26464 19610
rect 26516 19558 26528 19610
rect 26580 19558 34713 19610
rect 34765 19558 34777 19610
rect 34829 19558 34841 19610
rect 34893 19558 34905 19610
rect 34957 19558 34969 19610
rect 35021 19558 35027 19610
rect 1104 19536 35027 19558
rect 19242 19496 19248 19508
rect 19076 19468 19248 19496
rect 19076 19437 19104 19468
rect 19242 19456 19248 19468
rect 19300 19456 19306 19508
rect 19426 19456 19432 19508
rect 19484 19456 19490 19508
rect 20070 19456 20076 19508
rect 20128 19496 20134 19508
rect 20993 19499 21051 19505
rect 20993 19496 21005 19499
rect 20128 19468 21005 19496
rect 20128 19456 20134 19468
rect 20993 19465 21005 19468
rect 21039 19465 21051 19499
rect 20993 19459 21051 19465
rect 19061 19431 19119 19437
rect 19061 19397 19073 19431
rect 19107 19397 19119 19431
rect 19061 19391 19119 19397
rect 17221 19363 17279 19369
rect 17221 19329 17233 19363
rect 17267 19329 17279 19363
rect 17221 19323 17279 19329
rect 17405 19363 17463 19369
rect 17405 19329 17417 19363
rect 17451 19360 17463 19363
rect 18322 19360 18328 19372
rect 17451 19332 18328 19360
rect 17451 19329 17463 19332
rect 17405 19323 17463 19329
rect 17126 19184 17132 19236
rect 17184 19224 17190 19236
rect 17236 19224 17264 19323
rect 18322 19320 18328 19332
rect 18380 19320 18386 19372
rect 18690 19320 18696 19372
rect 18748 19360 18754 19372
rect 18877 19363 18935 19369
rect 18877 19360 18889 19363
rect 18748 19332 18889 19360
rect 18748 19320 18754 19332
rect 18877 19329 18889 19332
rect 18923 19329 18935 19363
rect 18877 19323 18935 19329
rect 17313 19295 17371 19301
rect 17313 19261 17325 19295
rect 17359 19292 17371 19295
rect 18230 19292 18236 19304
rect 17359 19264 18236 19292
rect 17359 19261 17371 19264
rect 17313 19255 17371 19261
rect 18230 19252 18236 19264
rect 18288 19252 18294 19304
rect 18892 19292 18920 19323
rect 18966 19320 18972 19372
rect 19024 19320 19030 19372
rect 19245 19363 19303 19369
rect 19245 19329 19257 19363
rect 19291 19360 19303 19363
rect 19444 19360 19472 19456
rect 20898 19428 20904 19440
rect 19291 19332 19472 19360
rect 19536 19400 20904 19428
rect 19291 19329 19303 19332
rect 19245 19323 19303 19329
rect 19334 19292 19340 19304
rect 18892 19264 19340 19292
rect 19334 19252 19340 19264
rect 19392 19252 19398 19304
rect 19536 19224 19564 19400
rect 20898 19388 20904 19400
rect 20956 19388 20962 19440
rect 19613 19363 19671 19369
rect 19613 19329 19625 19363
rect 19659 19360 19671 19363
rect 19702 19360 19708 19372
rect 19659 19332 19708 19360
rect 19659 19329 19671 19332
rect 19613 19323 19671 19329
rect 19702 19320 19708 19332
rect 19760 19320 19766 19372
rect 19880 19363 19938 19369
rect 19880 19329 19892 19363
rect 19926 19360 19938 19363
rect 20162 19360 20168 19372
rect 19926 19332 20168 19360
rect 19926 19329 19938 19332
rect 19880 19323 19938 19329
rect 20162 19320 20168 19332
rect 20220 19320 20226 19372
rect 21008 19360 21036 19459
rect 21358 19456 21364 19508
rect 21416 19496 21422 19508
rect 21637 19499 21695 19505
rect 21637 19496 21649 19499
rect 21416 19468 21649 19496
rect 21416 19456 21422 19468
rect 21637 19465 21649 19468
rect 21683 19465 21695 19499
rect 21637 19459 21695 19465
rect 21652 19428 21680 19459
rect 21910 19456 21916 19508
rect 21968 19496 21974 19508
rect 23201 19499 23259 19505
rect 23201 19496 23213 19499
rect 21968 19468 23213 19496
rect 21968 19456 21974 19468
rect 23201 19465 23213 19468
rect 23247 19465 23259 19499
rect 23201 19459 23259 19465
rect 21818 19428 21824 19440
rect 21652 19400 21824 19428
rect 21818 19388 21824 19400
rect 21876 19428 21882 19440
rect 22833 19431 22891 19437
rect 21876 19400 22048 19428
rect 21876 19388 21882 19400
rect 21082 19360 21088 19372
rect 21008 19332 21088 19360
rect 21082 19320 21088 19332
rect 21140 19360 21146 19372
rect 21269 19363 21327 19369
rect 21269 19360 21281 19363
rect 21140 19332 21281 19360
rect 21140 19320 21146 19332
rect 21269 19329 21281 19332
rect 21315 19329 21327 19363
rect 21269 19323 21327 19329
rect 21450 19320 21456 19372
rect 21508 19360 21514 19372
rect 22020 19369 22048 19400
rect 22833 19397 22845 19431
rect 22879 19428 22891 19431
rect 23014 19428 23020 19440
rect 22879 19400 23020 19428
rect 22879 19397 22891 19400
rect 22833 19391 22891 19397
rect 23014 19388 23020 19400
rect 23072 19388 23078 19440
rect 23216 19428 23244 19459
rect 24854 19456 24860 19508
rect 24912 19496 24918 19508
rect 25682 19496 25688 19508
rect 24912 19468 25688 19496
rect 24912 19456 24918 19468
rect 25682 19456 25688 19468
rect 25740 19496 25746 19508
rect 26329 19499 26387 19505
rect 26329 19496 26341 19499
rect 25740 19468 26341 19496
rect 25740 19456 25746 19468
rect 26329 19465 26341 19468
rect 26375 19465 26387 19499
rect 26329 19459 26387 19465
rect 27154 19456 27160 19508
rect 27212 19496 27218 19508
rect 27341 19499 27399 19505
rect 27341 19496 27353 19499
rect 27212 19468 27353 19496
rect 27212 19456 27218 19468
rect 27341 19465 27353 19468
rect 27387 19465 27399 19499
rect 27341 19459 27399 19465
rect 29362 19456 29368 19508
rect 29420 19456 29426 19508
rect 30469 19499 30527 19505
rect 30469 19465 30481 19499
rect 30515 19465 30527 19499
rect 30469 19459 30527 19465
rect 28166 19428 28172 19440
rect 23216 19400 24900 19428
rect 24872 19372 24900 19400
rect 27586 19400 28172 19428
rect 21913 19363 21971 19369
rect 21913 19360 21925 19363
rect 21508 19332 21925 19360
rect 21508 19320 21514 19332
rect 21913 19329 21925 19332
rect 21959 19329 21971 19363
rect 21913 19323 21971 19329
rect 22005 19363 22063 19369
rect 22005 19329 22017 19363
rect 22051 19329 22063 19363
rect 22005 19323 22063 19329
rect 22189 19363 22247 19369
rect 22189 19329 22201 19363
rect 22235 19360 22247 19363
rect 22370 19360 22376 19372
rect 22235 19332 22376 19360
rect 22235 19329 22247 19332
rect 22189 19323 22247 19329
rect 22370 19320 22376 19332
rect 22428 19320 22434 19372
rect 22738 19320 22744 19372
rect 22796 19360 22802 19372
rect 23382 19360 23388 19372
rect 22796 19332 23388 19360
rect 22796 19320 22802 19332
rect 23382 19320 23388 19332
rect 23440 19320 23446 19372
rect 23842 19320 23848 19372
rect 23900 19360 23906 19372
rect 24590 19363 24648 19369
rect 24590 19360 24602 19363
rect 23900 19332 24602 19360
rect 23900 19320 23906 19332
rect 24590 19329 24602 19332
rect 24636 19329 24648 19363
rect 24590 19323 24648 19329
rect 24854 19320 24860 19372
rect 24912 19320 24918 19372
rect 24949 19363 25007 19369
rect 24949 19329 24961 19363
rect 24995 19360 25007 19363
rect 25038 19360 25044 19372
rect 24995 19332 25044 19360
rect 24995 19329 25007 19332
rect 24949 19323 25007 19329
rect 25038 19320 25044 19332
rect 25096 19320 25102 19372
rect 25216 19363 25274 19369
rect 25216 19329 25228 19363
rect 25262 19360 25274 19363
rect 25498 19360 25504 19372
rect 25262 19332 25504 19360
rect 25262 19329 25274 19332
rect 25216 19323 25274 19329
rect 25498 19320 25504 19332
rect 25556 19320 25562 19372
rect 26786 19320 26792 19372
rect 26844 19360 26850 19372
rect 26973 19363 27031 19369
rect 26973 19360 26985 19363
rect 26844 19332 26985 19360
rect 26844 19320 26850 19332
rect 26973 19329 26985 19332
rect 27019 19329 27031 19363
rect 26973 19323 27031 19329
rect 27157 19363 27215 19369
rect 27157 19329 27169 19363
rect 27203 19360 27215 19363
rect 27586 19360 27614 19400
rect 28166 19388 28172 19400
rect 28224 19388 28230 19440
rect 29270 19428 29276 19440
rect 28920 19400 29276 19428
rect 27203 19332 27614 19360
rect 27203 19329 27215 19332
rect 27157 19323 27215 19329
rect 21358 19252 21364 19304
rect 21416 19252 21422 19304
rect 17184 19196 19564 19224
rect 22097 19227 22155 19233
rect 17184 19184 17190 19196
rect 18248 19168 18276 19196
rect 22097 19193 22109 19227
rect 22143 19224 22155 19227
rect 22186 19224 22192 19236
rect 22143 19196 22192 19224
rect 22143 19193 22155 19196
rect 22097 19187 22155 19193
rect 22186 19184 22192 19196
rect 22244 19184 22250 19236
rect 18230 19116 18236 19168
rect 18288 19116 18294 19168
rect 18693 19159 18751 19165
rect 18693 19125 18705 19159
rect 18739 19156 18751 19159
rect 19150 19156 19156 19168
rect 18739 19128 19156 19156
rect 18739 19125 18751 19128
rect 18693 19119 18751 19125
rect 19150 19116 19156 19128
rect 19208 19116 19214 19168
rect 22373 19159 22431 19165
rect 22373 19125 22385 19159
rect 22419 19156 22431 19159
rect 22462 19156 22468 19168
rect 22419 19128 22468 19156
rect 22419 19125 22431 19128
rect 22373 19119 22431 19125
rect 22462 19116 22468 19128
rect 22520 19116 22526 19168
rect 22554 19116 22560 19168
rect 22612 19116 22618 19168
rect 23477 19159 23535 19165
rect 23477 19125 23489 19159
rect 23523 19156 23535 19159
rect 23658 19156 23664 19168
rect 23523 19128 23664 19156
rect 23523 19125 23535 19128
rect 23477 19119 23535 19125
rect 23658 19116 23664 19128
rect 23716 19116 23722 19168
rect 25590 19116 25596 19168
rect 25648 19156 25654 19168
rect 26142 19156 26148 19168
rect 25648 19128 26148 19156
rect 25648 19116 25654 19128
rect 26142 19116 26148 19128
rect 26200 19156 26206 19168
rect 27172 19156 27200 19323
rect 28258 19320 28264 19372
rect 28316 19320 28322 19372
rect 28718 19320 28724 19372
rect 28776 19320 28782 19372
rect 28920 19369 28948 19400
rect 29270 19388 29276 19400
rect 29328 19388 29334 19440
rect 30484 19428 30512 19459
rect 31938 19456 31944 19508
rect 31996 19496 32002 19508
rect 32858 19496 32864 19508
rect 31996 19468 32864 19496
rect 31996 19456 32002 19468
rect 32858 19456 32864 19468
rect 32916 19456 32922 19508
rect 33134 19456 33140 19508
rect 33192 19496 33198 19508
rect 33689 19499 33747 19505
rect 33689 19496 33701 19499
rect 33192 19468 33701 19496
rect 33192 19456 33198 19468
rect 33689 19465 33701 19468
rect 33735 19465 33747 19499
rect 33689 19459 33747 19465
rect 30806 19431 30864 19437
rect 30806 19428 30818 19431
rect 30484 19400 30818 19428
rect 30806 19397 30818 19400
rect 30852 19397 30864 19431
rect 30806 19391 30864 19397
rect 32576 19431 32634 19437
rect 32576 19397 32588 19431
rect 32622 19428 32634 19431
rect 33042 19428 33048 19440
rect 32622 19400 33048 19428
rect 32622 19397 32634 19400
rect 32576 19391 32634 19397
rect 33042 19388 33048 19400
rect 33100 19388 33106 19440
rect 28905 19363 28963 19369
rect 28905 19329 28917 19363
rect 28951 19329 28963 19363
rect 28905 19323 28963 19329
rect 28994 19320 29000 19372
rect 29052 19320 29058 19372
rect 29086 19320 29092 19372
rect 29144 19320 29150 19372
rect 30285 19363 30343 19369
rect 30285 19329 30297 19363
rect 30331 19360 30343 19363
rect 31202 19360 31208 19372
rect 30331 19332 31208 19360
rect 30331 19329 30343 19332
rect 30285 19323 30343 19329
rect 31202 19320 31208 19332
rect 31260 19320 31266 19372
rect 30561 19295 30619 19301
rect 30561 19261 30573 19295
rect 30607 19261 30619 19295
rect 32306 19292 32312 19304
rect 30561 19255 30619 19261
rect 31726 19264 32312 19292
rect 26200 19128 27200 19156
rect 26200 19116 26206 19128
rect 28442 19116 28448 19168
rect 28500 19116 28506 19168
rect 30576 19156 30604 19255
rect 30834 19156 30840 19168
rect 30576 19128 30840 19156
rect 30834 19116 30840 19128
rect 30892 19156 30898 19168
rect 31726 19156 31754 19264
rect 32306 19252 32312 19264
rect 32364 19252 32370 19304
rect 30892 19128 31754 19156
rect 30892 19116 30898 19128
rect 1104 19066 34868 19088
rect 1104 19014 5170 19066
rect 5222 19014 5234 19066
rect 5286 19014 5298 19066
rect 5350 19014 5362 19066
rect 5414 19014 5426 19066
rect 5478 19014 13611 19066
rect 13663 19014 13675 19066
rect 13727 19014 13739 19066
rect 13791 19014 13803 19066
rect 13855 19014 13867 19066
rect 13919 19014 22052 19066
rect 22104 19014 22116 19066
rect 22168 19014 22180 19066
rect 22232 19014 22244 19066
rect 22296 19014 22308 19066
rect 22360 19014 30493 19066
rect 30545 19014 30557 19066
rect 30609 19014 30621 19066
rect 30673 19014 30685 19066
rect 30737 19014 30749 19066
rect 30801 19014 34868 19066
rect 1104 18992 34868 19014
rect 17957 18955 18015 18961
rect 17957 18921 17969 18955
rect 18003 18952 18015 18955
rect 18322 18952 18328 18964
rect 18003 18924 18328 18952
rect 18003 18921 18015 18924
rect 17957 18915 18015 18921
rect 18322 18912 18328 18924
rect 18380 18912 18386 18964
rect 18966 18912 18972 18964
rect 19024 18912 19030 18964
rect 19702 18952 19708 18964
rect 19076 18924 19708 18952
rect 19076 18884 19104 18924
rect 19702 18912 19708 18924
rect 19760 18912 19766 18964
rect 20162 18912 20168 18964
rect 20220 18912 20226 18964
rect 20530 18912 20536 18964
rect 20588 18952 20594 18964
rect 20806 18952 20812 18964
rect 20588 18924 20812 18952
rect 20588 18912 20594 18924
rect 20806 18912 20812 18924
rect 20864 18912 20870 18964
rect 21361 18955 21419 18961
rect 21361 18921 21373 18955
rect 21407 18952 21419 18955
rect 21450 18952 21456 18964
rect 21407 18924 21456 18952
rect 21407 18921 21419 18924
rect 21361 18915 21419 18921
rect 21450 18912 21456 18924
rect 21508 18912 21514 18964
rect 21726 18912 21732 18964
rect 21784 18912 21790 18964
rect 22922 18912 22928 18964
rect 22980 18912 22986 18964
rect 23566 18912 23572 18964
rect 23624 18912 23630 18964
rect 23842 18912 23848 18964
rect 23900 18912 23906 18964
rect 28258 18912 28264 18964
rect 28316 18952 28322 18964
rect 28813 18955 28871 18961
rect 28813 18952 28825 18955
rect 28316 18924 28825 18952
rect 28316 18912 28322 18924
rect 28813 18921 28825 18924
rect 28859 18921 28871 18955
rect 28813 18915 28871 18921
rect 28994 18912 29000 18964
rect 29052 18952 29058 18964
rect 29549 18955 29607 18961
rect 29549 18952 29561 18955
rect 29052 18924 29561 18952
rect 29052 18912 29058 18924
rect 29549 18921 29561 18924
rect 29595 18921 29607 18955
rect 29549 18915 29607 18921
rect 29638 18912 29644 18964
rect 29696 18952 29702 18964
rect 30009 18955 30067 18961
rect 30009 18952 30021 18955
rect 29696 18924 30021 18952
rect 29696 18912 29702 18924
rect 30009 18921 30021 18924
rect 30055 18952 30067 18955
rect 30055 18924 30788 18952
rect 30055 18921 30067 18924
rect 30009 18915 30067 18921
rect 17144 18856 19104 18884
rect 21284 18856 22094 18884
rect 16117 18751 16175 18757
rect 16117 18717 16129 18751
rect 16163 18748 16175 18751
rect 16206 18748 16212 18760
rect 16163 18720 16212 18748
rect 16163 18717 16175 18720
rect 16117 18711 16175 18717
rect 16206 18708 16212 18720
rect 16264 18748 16270 18760
rect 17144 18748 17172 18856
rect 18966 18776 18972 18828
rect 19024 18816 19030 18828
rect 19521 18819 19579 18825
rect 19521 18816 19533 18819
rect 19024 18788 19533 18816
rect 19024 18776 19030 18788
rect 19521 18785 19533 18788
rect 19567 18785 19579 18819
rect 21082 18816 21088 18828
rect 19521 18779 19579 18785
rect 20456 18788 21088 18816
rect 16264 18720 17172 18748
rect 16264 18708 16270 18720
rect 17218 18708 17224 18760
rect 17276 18748 17282 18760
rect 17773 18751 17831 18757
rect 17773 18748 17785 18751
rect 17276 18720 17785 18748
rect 17276 18708 17282 18720
rect 17773 18717 17785 18720
rect 17819 18717 17831 18751
rect 18049 18751 18107 18757
rect 18049 18748 18061 18751
rect 17773 18711 17831 18717
rect 17972 18720 18061 18748
rect 16384 18683 16442 18689
rect 16384 18649 16396 18683
rect 16430 18680 16442 18683
rect 17589 18683 17647 18689
rect 17589 18680 17601 18683
rect 16430 18652 17601 18680
rect 16430 18649 16442 18652
rect 16384 18643 16442 18649
rect 17589 18649 17601 18652
rect 17635 18649 17647 18683
rect 17972 18680 18000 18720
rect 18049 18717 18061 18720
rect 18095 18717 18107 18751
rect 18049 18711 18107 18717
rect 19061 18751 19119 18757
rect 19061 18717 19073 18751
rect 19107 18717 19119 18751
rect 19061 18711 19119 18717
rect 17589 18643 17647 18649
rect 17696 18652 18000 18680
rect 17696 18624 17724 18652
rect 17497 18615 17555 18621
rect 17497 18581 17509 18615
rect 17543 18612 17555 18615
rect 17678 18612 17684 18624
rect 17543 18584 17684 18612
rect 17543 18581 17555 18584
rect 17497 18575 17555 18581
rect 17678 18572 17684 18584
rect 17736 18572 17742 18624
rect 19076 18612 19104 18711
rect 19150 18708 19156 18760
rect 19208 18748 19214 18760
rect 19245 18751 19303 18757
rect 19245 18748 19257 18751
rect 19208 18720 19257 18748
rect 19208 18708 19214 18720
rect 19245 18717 19257 18720
rect 19291 18717 19303 18751
rect 19245 18711 19303 18717
rect 19334 18708 19340 18760
rect 19392 18748 19398 18760
rect 19429 18751 19487 18757
rect 19429 18748 19441 18751
rect 19392 18720 19441 18748
rect 19392 18708 19398 18720
rect 19429 18717 19441 18720
rect 19475 18717 19487 18751
rect 19429 18711 19487 18717
rect 19610 18708 19616 18760
rect 19668 18708 19674 18760
rect 19794 18708 19800 18760
rect 19852 18708 19858 18760
rect 20456 18757 20484 18788
rect 21082 18776 21088 18788
rect 21140 18776 21146 18828
rect 21284 18825 21312 18856
rect 21269 18819 21327 18825
rect 21269 18785 21281 18819
rect 21315 18785 21327 18819
rect 21269 18779 21327 18785
rect 21450 18776 21456 18828
rect 21508 18776 21514 18828
rect 21542 18776 21548 18828
rect 21600 18776 21606 18828
rect 20441 18751 20499 18757
rect 20441 18717 20453 18751
rect 20487 18717 20499 18751
rect 20441 18711 20499 18717
rect 20530 18708 20536 18760
rect 20588 18708 20594 18760
rect 20625 18751 20683 18757
rect 20625 18717 20637 18751
rect 20671 18748 20683 18751
rect 20714 18748 20720 18760
rect 20671 18720 20720 18748
rect 20671 18717 20683 18720
rect 20625 18711 20683 18717
rect 20714 18708 20720 18720
rect 20772 18708 20778 18760
rect 20809 18751 20867 18757
rect 20809 18717 20821 18751
rect 20855 18717 20867 18751
rect 21100 18748 21128 18776
rect 21177 18751 21235 18757
rect 21177 18748 21189 18751
rect 21100 18720 21189 18748
rect 20809 18711 20867 18717
rect 21177 18717 21189 18720
rect 21223 18717 21235 18751
rect 21177 18711 21235 18717
rect 20824 18680 20852 18711
rect 21818 18708 21824 18760
rect 21876 18708 21882 18760
rect 22066 18748 22094 18856
rect 22554 18776 22560 18828
rect 22612 18816 22618 18828
rect 23584 18816 23612 18912
rect 28721 18887 28779 18893
rect 28721 18853 28733 18887
rect 28767 18884 28779 18887
rect 28767 18856 29132 18884
rect 28767 18853 28779 18856
rect 28721 18847 28779 18853
rect 29104 18828 29132 18856
rect 22612 18788 23060 18816
rect 22612 18776 22618 18788
rect 22646 18748 22652 18760
rect 22066 18720 22652 18748
rect 22646 18708 22652 18720
rect 22704 18748 22710 18760
rect 23032 18757 23060 18788
rect 23216 18788 23612 18816
rect 23216 18757 23244 18788
rect 26602 18776 26608 18828
rect 26660 18816 26666 18828
rect 26660 18788 27476 18816
rect 26660 18776 26666 18788
rect 27448 18760 27476 18788
rect 29086 18776 29092 18828
rect 29144 18816 29150 18828
rect 30760 18825 30788 18924
rect 31202 18912 31208 18964
rect 31260 18912 31266 18964
rect 32585 18955 32643 18961
rect 32585 18921 32597 18955
rect 32631 18952 32643 18955
rect 33226 18952 33232 18964
rect 32631 18924 33232 18952
rect 32631 18921 32643 18924
rect 32585 18915 32643 18921
rect 33226 18912 33232 18924
rect 33284 18912 33290 18964
rect 29181 18819 29239 18825
rect 29181 18816 29193 18819
rect 29144 18788 29193 18816
rect 29144 18776 29150 18788
rect 29181 18785 29193 18788
rect 29227 18785 29239 18819
rect 30745 18819 30803 18825
rect 29181 18779 29239 18785
rect 29472 18788 30604 18816
rect 22833 18751 22891 18757
rect 22833 18748 22845 18751
rect 22704 18720 22845 18748
rect 22704 18708 22710 18720
rect 22833 18717 22845 18720
rect 22879 18717 22891 18751
rect 22833 18711 22891 18717
rect 23017 18751 23075 18757
rect 23017 18717 23029 18751
rect 23063 18717 23075 18751
rect 23017 18711 23075 18717
rect 23201 18751 23259 18757
rect 23201 18717 23213 18751
rect 23247 18717 23259 18751
rect 23201 18711 23259 18717
rect 23385 18751 23443 18757
rect 23385 18717 23397 18751
rect 23431 18717 23443 18751
rect 23385 18711 23443 18717
rect 23216 18680 23244 18711
rect 19904 18652 20760 18680
rect 20824 18652 23244 18680
rect 23400 18680 23428 18711
rect 23474 18708 23480 18760
rect 23532 18708 23538 18760
rect 23569 18751 23627 18757
rect 23569 18717 23581 18751
rect 23615 18748 23627 18751
rect 23658 18748 23664 18760
rect 23615 18720 23664 18748
rect 23615 18717 23627 18720
rect 23569 18711 23627 18717
rect 23658 18708 23664 18720
rect 23716 18708 23722 18760
rect 26878 18708 26884 18760
rect 26936 18748 26942 18760
rect 27249 18751 27307 18757
rect 27249 18748 27261 18751
rect 26936 18720 27261 18748
rect 26936 18708 26942 18720
rect 27249 18717 27261 18720
rect 27295 18717 27307 18751
rect 27249 18711 27307 18717
rect 27341 18751 27399 18757
rect 27341 18717 27353 18751
rect 27387 18717 27399 18751
rect 27341 18711 27399 18717
rect 23934 18680 23940 18692
rect 23400 18652 23940 18680
rect 19904 18612 19932 18652
rect 20732 18624 20760 18652
rect 23934 18640 23940 18652
rect 23992 18640 23998 18692
rect 19076 18584 19932 18612
rect 19978 18572 19984 18624
rect 20036 18572 20042 18624
rect 20714 18572 20720 18624
rect 20772 18572 20778 18624
rect 21174 18572 21180 18624
rect 21232 18612 21238 18624
rect 21545 18615 21603 18621
rect 21545 18612 21557 18615
rect 21232 18584 21557 18612
rect 21232 18572 21238 18584
rect 21545 18581 21557 18584
rect 21591 18581 21603 18615
rect 21545 18575 21603 18581
rect 21634 18572 21640 18624
rect 21692 18612 21698 18624
rect 21910 18612 21916 18624
rect 21692 18584 21916 18612
rect 21692 18572 21698 18584
rect 21910 18572 21916 18584
rect 21968 18612 21974 18624
rect 23658 18612 23664 18624
rect 21968 18584 23664 18612
rect 21968 18572 21974 18584
rect 23658 18572 23664 18584
rect 23716 18572 23722 18624
rect 27065 18615 27123 18621
rect 27065 18581 27077 18615
rect 27111 18612 27123 18615
rect 27356 18612 27384 18711
rect 27430 18708 27436 18760
rect 27488 18748 27494 18760
rect 28997 18751 29055 18757
rect 28997 18748 29009 18751
rect 27488 18720 29009 18748
rect 27488 18708 27494 18720
rect 28997 18717 29009 18720
rect 29043 18748 29055 18751
rect 29472 18748 29500 18788
rect 29043 18720 29500 18748
rect 29043 18717 29055 18720
rect 28997 18711 29055 18717
rect 29546 18708 29552 18760
rect 29604 18748 29610 18760
rect 29825 18751 29883 18757
rect 29825 18748 29837 18751
rect 29604 18720 29837 18748
rect 29604 18708 29610 18720
rect 29825 18717 29837 18720
rect 29871 18717 29883 18751
rect 29825 18711 29883 18717
rect 29917 18751 29975 18757
rect 29917 18717 29929 18751
rect 29963 18717 29975 18751
rect 29917 18711 29975 18717
rect 27614 18689 27620 18692
rect 27608 18643 27620 18689
rect 27614 18640 27620 18643
rect 27672 18640 27678 18692
rect 29178 18640 29184 18692
rect 29236 18680 29242 18692
rect 29932 18680 29960 18711
rect 30098 18708 30104 18760
rect 30156 18708 30162 18760
rect 30576 18757 30604 18788
rect 30745 18785 30757 18819
rect 30791 18785 30803 18819
rect 30745 18779 30803 18785
rect 31573 18819 31631 18825
rect 31573 18785 31585 18819
rect 31619 18816 31631 18819
rect 32122 18816 32128 18828
rect 31619 18788 32128 18816
rect 31619 18785 31631 18788
rect 31573 18779 31631 18785
rect 32122 18776 32128 18788
rect 32180 18776 32186 18828
rect 30285 18751 30343 18757
rect 30285 18717 30297 18751
rect 30331 18717 30343 18751
rect 30285 18711 30343 18717
rect 30561 18751 30619 18757
rect 30561 18717 30573 18751
rect 30607 18748 30619 18751
rect 30926 18748 30932 18760
rect 30607 18720 30932 18748
rect 30607 18717 30619 18720
rect 30561 18711 30619 18717
rect 29236 18652 29960 18680
rect 29236 18640 29242 18652
rect 28534 18612 28540 18624
rect 27111 18584 28540 18612
rect 27111 18581 27123 18584
rect 27065 18575 27123 18581
rect 28534 18572 28540 18584
rect 28592 18572 28598 18624
rect 29454 18572 29460 18624
rect 29512 18612 29518 18624
rect 30300 18612 30328 18711
rect 30926 18708 30932 18720
rect 30984 18708 30990 18760
rect 31294 18708 31300 18760
rect 31352 18748 31358 18760
rect 31389 18751 31447 18757
rect 31389 18748 31401 18751
rect 31352 18720 31401 18748
rect 31352 18708 31358 18720
rect 31389 18717 31401 18720
rect 31435 18748 31447 18751
rect 31435 18720 31754 18748
rect 31435 18717 31447 18720
rect 31389 18711 31447 18717
rect 31726 18680 31754 18720
rect 31938 18708 31944 18760
rect 31996 18748 32002 18760
rect 32217 18751 32275 18757
rect 32217 18748 32229 18751
rect 31996 18720 32229 18748
rect 31996 18708 32002 18720
rect 32217 18717 32229 18720
rect 32263 18717 32275 18751
rect 32217 18711 32275 18717
rect 32401 18751 32459 18757
rect 32401 18717 32413 18751
rect 32447 18717 32459 18751
rect 32401 18711 32459 18717
rect 32416 18680 32444 18711
rect 31726 18652 32444 18680
rect 29512 18584 30328 18612
rect 29512 18572 29518 18584
rect 30374 18572 30380 18624
rect 30432 18572 30438 18624
rect 1104 18522 35027 18544
rect 1104 18470 9390 18522
rect 9442 18470 9454 18522
rect 9506 18470 9518 18522
rect 9570 18470 9582 18522
rect 9634 18470 9646 18522
rect 9698 18470 17831 18522
rect 17883 18470 17895 18522
rect 17947 18470 17959 18522
rect 18011 18470 18023 18522
rect 18075 18470 18087 18522
rect 18139 18470 26272 18522
rect 26324 18470 26336 18522
rect 26388 18470 26400 18522
rect 26452 18470 26464 18522
rect 26516 18470 26528 18522
rect 26580 18470 34713 18522
rect 34765 18470 34777 18522
rect 34829 18470 34841 18522
rect 34893 18470 34905 18522
rect 34957 18470 34969 18522
rect 35021 18470 35027 18522
rect 1104 18448 35027 18470
rect 17129 18411 17187 18417
rect 17129 18377 17141 18411
rect 17175 18408 17187 18411
rect 17218 18408 17224 18420
rect 17175 18380 17224 18408
rect 17175 18377 17187 18380
rect 17129 18371 17187 18377
rect 17218 18368 17224 18380
rect 17276 18368 17282 18420
rect 17983 18411 18041 18417
rect 17983 18408 17995 18411
rect 17512 18380 17995 18408
rect 17037 18275 17095 18281
rect 17037 18241 17049 18275
rect 17083 18272 17095 18275
rect 17126 18272 17132 18284
rect 17083 18244 17132 18272
rect 17083 18241 17095 18244
rect 17037 18235 17095 18241
rect 17126 18232 17132 18244
rect 17184 18232 17190 18284
rect 17512 18281 17540 18380
rect 17983 18377 17995 18380
rect 18029 18408 18041 18411
rect 18322 18408 18328 18420
rect 18029 18380 18328 18408
rect 18029 18377 18041 18380
rect 17983 18371 18041 18377
rect 18322 18368 18328 18380
rect 18380 18368 18386 18420
rect 19610 18408 19616 18420
rect 18892 18380 19616 18408
rect 18892 18349 18920 18380
rect 19610 18368 19616 18380
rect 19668 18368 19674 18420
rect 19978 18368 19984 18420
rect 20036 18368 20042 18420
rect 20714 18368 20720 18420
rect 20772 18408 20778 18420
rect 21634 18408 21640 18420
rect 20772 18380 21640 18408
rect 20772 18368 20778 18380
rect 21634 18368 21640 18380
rect 21692 18368 21698 18420
rect 25498 18368 25504 18420
rect 25556 18368 25562 18420
rect 27525 18411 27583 18417
rect 27525 18377 27537 18411
rect 27571 18408 27583 18411
rect 27614 18408 27620 18420
rect 27571 18380 27620 18408
rect 27571 18377 27583 18380
rect 27525 18371 27583 18377
rect 27614 18368 27620 18380
rect 27672 18368 27678 18420
rect 29454 18408 29460 18420
rect 28184 18380 29460 18408
rect 17773 18343 17831 18349
rect 17773 18309 17785 18343
rect 17819 18340 17831 18343
rect 18877 18343 18935 18349
rect 17819 18312 18276 18340
rect 17819 18309 17831 18312
rect 17773 18303 17831 18309
rect 18248 18284 18276 18312
rect 18877 18309 18889 18343
rect 18923 18309 18935 18343
rect 19334 18340 19340 18352
rect 18877 18303 18935 18309
rect 19076 18312 19340 18340
rect 17221 18275 17279 18281
rect 17221 18241 17233 18275
rect 17267 18272 17279 18275
rect 17497 18275 17555 18281
rect 17267 18244 17356 18272
rect 17267 18241 17279 18244
rect 17221 18235 17279 18241
rect 17328 18077 17356 18244
rect 17497 18241 17509 18275
rect 17543 18241 17555 18275
rect 17497 18235 17555 18241
rect 18230 18232 18236 18284
rect 18288 18272 18294 18284
rect 18647 18275 18705 18281
rect 18647 18272 18659 18275
rect 18288 18244 18659 18272
rect 18288 18232 18294 18244
rect 18647 18241 18659 18244
rect 18693 18241 18705 18275
rect 18647 18235 18705 18241
rect 18782 18232 18788 18284
rect 18840 18232 18846 18284
rect 17678 18164 17684 18216
rect 17736 18164 17742 18216
rect 17696 18136 17724 18164
rect 18892 18136 18920 18303
rect 19076 18281 19104 18312
rect 19334 18300 19340 18312
rect 19392 18340 19398 18352
rect 19794 18340 19800 18352
rect 19392 18312 19800 18340
rect 19392 18300 19398 18312
rect 19794 18300 19800 18312
rect 19852 18300 19858 18352
rect 19060 18275 19118 18281
rect 19060 18241 19072 18275
rect 19106 18241 19118 18275
rect 19060 18235 19118 18241
rect 19153 18275 19211 18281
rect 19153 18241 19165 18275
rect 19199 18272 19211 18275
rect 19996 18272 20024 18368
rect 22388 18312 22784 18340
rect 22388 18284 22416 18312
rect 19199 18244 20024 18272
rect 19199 18241 19211 18244
rect 19153 18235 19211 18241
rect 20714 18232 20720 18284
rect 20772 18272 20778 18284
rect 20901 18275 20959 18281
rect 20901 18272 20913 18275
rect 20772 18244 20913 18272
rect 20772 18232 20778 18244
rect 20901 18241 20913 18244
rect 20947 18272 20959 18275
rect 21542 18272 21548 18284
rect 20947 18244 21548 18272
rect 20947 18241 20959 18244
rect 20901 18235 20959 18241
rect 21542 18232 21548 18244
rect 21600 18232 21606 18284
rect 22370 18232 22376 18284
rect 22428 18232 22434 18284
rect 22462 18232 22468 18284
rect 22520 18272 22526 18284
rect 22756 18281 22784 18312
rect 26160 18312 26740 18340
rect 22557 18275 22615 18281
rect 22557 18272 22569 18275
rect 22520 18244 22569 18272
rect 22520 18232 22526 18244
rect 22557 18241 22569 18244
rect 22603 18241 22615 18275
rect 22557 18235 22615 18241
rect 22741 18275 22799 18281
rect 22741 18241 22753 18275
rect 22787 18241 22799 18275
rect 22741 18235 22799 18241
rect 24946 18232 24952 18284
rect 25004 18232 25010 18284
rect 25777 18275 25835 18281
rect 25700 18247 25789 18275
rect 17696 18108 18920 18136
rect 17313 18071 17371 18077
rect 17313 18037 17325 18071
rect 17359 18068 17371 18071
rect 17494 18068 17500 18080
rect 17359 18040 17500 18068
rect 17359 18037 17371 18040
rect 17313 18031 17371 18037
rect 17494 18028 17500 18040
rect 17552 18028 17558 18080
rect 17972 18077 18000 18108
rect 20806 18096 20812 18148
rect 20864 18136 20870 18148
rect 21085 18139 21143 18145
rect 21085 18136 21097 18139
rect 20864 18108 21097 18136
rect 20864 18096 20870 18108
rect 21085 18105 21097 18108
rect 21131 18105 21143 18139
rect 25700 18136 25728 18247
rect 25777 18241 25789 18247
rect 25823 18241 25835 18275
rect 25777 18235 25835 18241
rect 25866 18232 25872 18284
rect 25924 18232 25930 18284
rect 25961 18275 26019 18281
rect 25961 18241 25973 18275
rect 26007 18272 26019 18275
rect 26050 18272 26056 18284
rect 26007 18244 26056 18272
rect 26007 18241 26019 18244
rect 25961 18235 26019 18241
rect 26050 18232 26056 18244
rect 26108 18232 26114 18284
rect 26160 18281 26188 18312
rect 26712 18284 26740 18312
rect 26145 18275 26203 18281
rect 26145 18241 26157 18275
rect 26191 18241 26203 18275
rect 26145 18235 26203 18241
rect 26421 18275 26479 18281
rect 26421 18241 26433 18275
rect 26467 18272 26479 18275
rect 26510 18272 26516 18284
rect 26467 18244 26516 18272
rect 26467 18241 26479 18244
rect 26421 18235 26479 18241
rect 26510 18232 26516 18244
rect 26568 18232 26574 18284
rect 26694 18232 26700 18284
rect 26752 18232 26758 18284
rect 26970 18232 26976 18284
rect 27028 18232 27034 18284
rect 27522 18232 27528 18284
rect 27580 18232 27586 18284
rect 28184 18281 28212 18380
rect 29454 18368 29460 18380
rect 29512 18368 29518 18420
rect 29638 18368 29644 18420
rect 29696 18368 29702 18420
rect 29730 18368 29736 18420
rect 29788 18408 29794 18420
rect 30098 18408 30104 18420
rect 29788 18380 30104 18408
rect 29788 18368 29794 18380
rect 30098 18368 30104 18380
rect 30156 18368 30162 18420
rect 28442 18300 28448 18352
rect 28500 18340 28506 18352
rect 28500 18312 28580 18340
rect 28500 18300 28506 18312
rect 28552 18281 28580 18312
rect 27709 18275 27767 18281
rect 27709 18241 27721 18275
rect 27755 18272 27767 18275
rect 27801 18275 27859 18281
rect 27801 18272 27813 18275
rect 27755 18244 27813 18272
rect 27755 18241 27767 18244
rect 27709 18235 27767 18241
rect 27801 18241 27813 18244
rect 27847 18241 27859 18275
rect 27801 18235 27859 18241
rect 27985 18275 28043 18281
rect 27985 18241 27997 18275
rect 28031 18241 28043 18275
rect 27985 18235 28043 18241
rect 28169 18275 28227 18281
rect 28169 18241 28181 18275
rect 28215 18241 28227 18275
rect 28169 18235 28227 18241
rect 28528 18275 28586 18281
rect 28528 18241 28540 18275
rect 28574 18241 28586 18275
rect 28528 18235 28586 18241
rect 26605 18207 26663 18213
rect 26605 18173 26617 18207
rect 26651 18173 26663 18207
rect 27540 18204 27568 18232
rect 28000 18204 28028 18235
rect 30374 18232 30380 18284
rect 30432 18272 30438 18284
rect 30846 18275 30904 18281
rect 30846 18272 30858 18275
rect 30432 18244 30858 18272
rect 30432 18232 30438 18244
rect 30846 18241 30858 18244
rect 30892 18241 30904 18275
rect 30846 18235 30904 18241
rect 27540 18176 28028 18204
rect 28261 18207 28319 18213
rect 26605 18167 26663 18173
rect 28261 18173 28273 18207
rect 28307 18173 28319 18207
rect 28261 18167 28319 18173
rect 31113 18207 31171 18213
rect 31113 18173 31125 18207
rect 31159 18173 31171 18207
rect 31113 18167 31171 18173
rect 25774 18136 25780 18148
rect 25700 18108 25780 18136
rect 21085 18099 21143 18105
rect 25774 18096 25780 18108
rect 25832 18136 25838 18148
rect 26620 18136 26648 18167
rect 25832 18108 26648 18136
rect 25832 18096 25838 18108
rect 17957 18071 18015 18077
rect 17957 18037 17969 18071
rect 18003 18037 18015 18071
rect 17957 18031 18015 18037
rect 18141 18071 18199 18077
rect 18141 18037 18153 18071
rect 18187 18068 18199 18071
rect 18414 18068 18420 18080
rect 18187 18040 18420 18068
rect 18187 18037 18199 18040
rect 18141 18031 18199 18037
rect 18414 18028 18420 18040
rect 18472 18028 18478 18080
rect 18506 18028 18512 18080
rect 18564 18028 18570 18080
rect 22738 18028 22744 18080
rect 22796 18028 22802 18080
rect 24670 18028 24676 18080
rect 24728 18068 24734 18080
rect 24765 18071 24823 18077
rect 24765 18068 24777 18071
rect 24728 18040 24777 18068
rect 24728 18028 24734 18040
rect 24765 18037 24777 18040
rect 24811 18037 24823 18071
rect 24765 18031 24823 18037
rect 26234 18028 26240 18080
rect 26292 18028 26298 18080
rect 27157 18071 27215 18077
rect 27157 18037 27169 18071
rect 27203 18068 27215 18071
rect 27890 18068 27896 18080
rect 27203 18040 27896 18068
rect 27203 18037 27215 18040
rect 27157 18031 27215 18037
rect 27890 18028 27896 18040
rect 27948 18028 27954 18080
rect 28276 18068 28304 18167
rect 30834 18068 30840 18080
rect 28276 18040 30840 18068
rect 30834 18028 30840 18040
rect 30892 18068 30898 18080
rect 31128 18068 31156 18167
rect 31386 18068 31392 18080
rect 30892 18040 31392 18068
rect 30892 18028 30898 18040
rect 31386 18028 31392 18040
rect 31444 18028 31450 18080
rect 1104 17978 34868 18000
rect 1104 17926 5170 17978
rect 5222 17926 5234 17978
rect 5286 17926 5298 17978
rect 5350 17926 5362 17978
rect 5414 17926 5426 17978
rect 5478 17926 13611 17978
rect 13663 17926 13675 17978
rect 13727 17926 13739 17978
rect 13791 17926 13803 17978
rect 13855 17926 13867 17978
rect 13919 17926 22052 17978
rect 22104 17926 22116 17978
rect 22168 17926 22180 17978
rect 22232 17926 22244 17978
rect 22296 17926 22308 17978
rect 22360 17926 30493 17978
rect 30545 17926 30557 17978
rect 30609 17926 30621 17978
rect 30673 17926 30685 17978
rect 30737 17926 30749 17978
rect 30801 17926 34868 17978
rect 1104 17904 34868 17926
rect 17494 17824 17500 17876
rect 17552 17824 17558 17876
rect 18049 17867 18107 17873
rect 18049 17833 18061 17867
rect 18095 17864 18107 17867
rect 18138 17864 18144 17876
rect 18095 17836 18144 17864
rect 18095 17833 18107 17836
rect 18049 17827 18107 17833
rect 18138 17824 18144 17836
rect 18196 17824 18202 17876
rect 19334 17824 19340 17876
rect 19392 17824 19398 17876
rect 22094 17864 22100 17876
rect 19444 17836 22100 17864
rect 18156 17796 18184 17824
rect 18156 17768 18460 17796
rect 15197 17731 15255 17737
rect 15197 17697 15209 17731
rect 15243 17728 15255 17731
rect 16114 17728 16120 17740
rect 15243 17700 16120 17728
rect 15243 17697 15255 17700
rect 15197 17691 15255 17697
rect 16114 17688 16120 17700
rect 16172 17688 16178 17740
rect 18325 17731 18383 17737
rect 18325 17728 18337 17731
rect 17328 17700 18337 17728
rect 15562 17620 15568 17672
rect 15620 17620 15626 17672
rect 17328 17669 17356 17700
rect 18325 17697 18337 17700
rect 18371 17697 18383 17731
rect 18325 17691 18383 17697
rect 18432 17669 18460 17768
rect 19444 17669 19472 17836
rect 22094 17824 22100 17836
rect 22152 17824 22158 17876
rect 22554 17864 22560 17876
rect 22204 17836 22560 17864
rect 20579 17799 20637 17805
rect 20579 17796 20591 17799
rect 19720 17768 20591 17796
rect 17313 17663 17371 17669
rect 17313 17629 17325 17663
rect 17359 17629 17371 17663
rect 17313 17623 17371 17629
rect 17589 17663 17647 17669
rect 17589 17629 17601 17663
rect 17635 17660 17647 17663
rect 18233 17663 18291 17669
rect 17635 17632 18184 17660
rect 17635 17629 17647 17632
rect 17589 17623 17647 17629
rect 16114 17552 16120 17604
rect 16172 17552 16178 17604
rect 16991 17595 17049 17601
rect 16991 17561 17003 17595
rect 17037 17592 17049 17595
rect 17773 17595 17831 17601
rect 17773 17592 17785 17595
rect 17037 17564 17785 17592
rect 17037 17561 17049 17564
rect 16991 17555 17049 17561
rect 17773 17561 17785 17564
rect 17819 17561 17831 17595
rect 17773 17555 17831 17561
rect 17126 17484 17132 17536
rect 17184 17484 17190 17536
rect 18156 17524 18184 17632
rect 18233 17629 18245 17663
rect 18279 17629 18291 17663
rect 18233 17623 18291 17629
rect 18417 17663 18475 17669
rect 18417 17629 18429 17663
rect 18463 17629 18475 17663
rect 18417 17623 18475 17629
rect 19429 17663 19487 17669
rect 19429 17629 19441 17663
rect 19475 17629 19487 17663
rect 19429 17623 19487 17629
rect 18248 17592 18276 17623
rect 18248 17564 18460 17592
rect 18432 17536 18460 17564
rect 19720 17536 19748 17768
rect 20579 17765 20591 17768
rect 20625 17796 20637 17799
rect 21177 17799 21235 17805
rect 21177 17796 21189 17799
rect 20625 17768 21189 17796
rect 20625 17765 20637 17768
rect 20579 17759 20637 17765
rect 21177 17765 21189 17768
rect 21223 17796 21235 17799
rect 21821 17799 21879 17805
rect 21821 17796 21833 17799
rect 21223 17768 21833 17796
rect 21223 17765 21235 17768
rect 21177 17759 21235 17765
rect 21821 17765 21833 17768
rect 21867 17765 21879 17799
rect 21821 17759 21879 17765
rect 20441 17731 20499 17737
rect 20441 17697 20453 17731
rect 20487 17728 20499 17731
rect 20487 17700 21036 17728
rect 20487 17697 20499 17700
rect 20441 17691 20499 17697
rect 21008 17672 21036 17700
rect 21450 17688 21456 17740
rect 21508 17728 21514 17740
rect 22204 17728 22232 17836
rect 22554 17824 22560 17836
rect 22612 17824 22618 17876
rect 22738 17824 22744 17876
rect 22796 17864 22802 17876
rect 23106 17864 23112 17876
rect 22796 17836 23112 17864
rect 22796 17824 22802 17836
rect 23106 17824 23112 17836
rect 23164 17864 23170 17876
rect 23845 17867 23903 17873
rect 23845 17864 23857 17867
rect 23164 17836 23857 17864
rect 23164 17824 23170 17836
rect 23845 17833 23857 17836
rect 23891 17833 23903 17867
rect 23845 17827 23903 17833
rect 23934 17824 23940 17876
rect 23992 17824 23998 17876
rect 25774 17824 25780 17876
rect 25832 17824 25838 17876
rect 29454 17824 29460 17876
rect 29512 17824 29518 17876
rect 29825 17867 29883 17873
rect 29825 17833 29837 17867
rect 29871 17864 29883 17867
rect 30374 17864 30380 17876
rect 29871 17836 30380 17864
rect 29871 17833 29883 17836
rect 29825 17827 29883 17833
rect 30374 17824 30380 17836
rect 30432 17824 30438 17876
rect 22462 17756 22468 17808
rect 22520 17796 22526 17808
rect 23290 17796 23296 17808
rect 22520 17768 23296 17796
rect 22520 17756 22526 17768
rect 23290 17756 23296 17768
rect 23348 17756 23354 17808
rect 29472 17796 29500 17824
rect 30101 17799 30159 17805
rect 30101 17796 30113 17799
rect 29472 17768 30113 17796
rect 30101 17765 30113 17768
rect 30147 17765 30159 17799
rect 30101 17759 30159 17765
rect 30282 17756 30288 17808
rect 30340 17756 30346 17808
rect 24029 17731 24087 17737
rect 24029 17728 24041 17731
rect 21508 17700 22232 17728
rect 21508 17688 21514 17700
rect 20165 17663 20223 17669
rect 20165 17629 20177 17663
rect 20211 17629 20223 17663
rect 20165 17623 20223 17629
rect 20180 17592 20208 17623
rect 20254 17620 20260 17672
rect 20312 17660 20318 17672
rect 20622 17660 20628 17672
rect 20312 17632 20628 17660
rect 20312 17620 20318 17632
rect 20622 17620 20628 17632
rect 20680 17620 20686 17672
rect 20717 17663 20775 17669
rect 20717 17629 20729 17663
rect 20763 17629 20775 17663
rect 20717 17623 20775 17629
rect 20732 17592 20760 17623
rect 20806 17620 20812 17672
rect 20864 17620 20870 17672
rect 20990 17620 20996 17672
rect 21048 17620 21054 17672
rect 21560 17669 21588 17700
rect 21269 17663 21327 17669
rect 21269 17629 21281 17663
rect 21315 17629 21327 17663
rect 21269 17623 21327 17629
rect 21361 17663 21419 17669
rect 21361 17629 21373 17663
rect 21407 17629 21419 17663
rect 21361 17623 21419 17629
rect 21545 17663 21603 17669
rect 21545 17629 21557 17663
rect 21591 17629 21603 17663
rect 21545 17623 21603 17629
rect 21637 17663 21695 17669
rect 21637 17629 21649 17663
rect 21683 17660 21695 17663
rect 21726 17660 21732 17672
rect 21683 17632 21732 17660
rect 21683 17629 21695 17632
rect 21637 17623 21695 17629
rect 20898 17592 20904 17604
rect 20180 17564 20668 17592
rect 20732 17564 20904 17592
rect 20180 17536 20208 17564
rect 18230 17524 18236 17536
rect 18156 17496 18236 17524
rect 18230 17484 18236 17496
rect 18288 17484 18294 17536
rect 18414 17484 18420 17536
rect 18472 17484 18478 17536
rect 19702 17484 19708 17536
rect 19760 17484 19766 17536
rect 20070 17484 20076 17536
rect 20128 17484 20134 17536
rect 20162 17484 20168 17536
rect 20220 17484 20226 17536
rect 20346 17484 20352 17536
rect 20404 17484 20410 17536
rect 20640 17524 20668 17564
rect 20898 17552 20904 17564
rect 20956 17592 20962 17604
rect 21284 17592 21312 17623
rect 20956 17564 21312 17592
rect 20956 17552 20962 17564
rect 21376 17524 21404 17623
rect 21726 17620 21732 17632
rect 21784 17620 21790 17672
rect 21821 17663 21879 17669
rect 21821 17629 21833 17663
rect 21867 17629 21879 17663
rect 21821 17623 21879 17629
rect 21836 17536 21864 17623
rect 21910 17620 21916 17672
rect 21968 17660 21974 17672
rect 22204 17669 22232 17700
rect 22388 17700 23520 17728
rect 22388 17672 22416 17700
rect 22005 17663 22063 17669
rect 22005 17660 22017 17663
rect 21968 17632 22017 17660
rect 21968 17620 21974 17632
rect 22005 17629 22017 17632
rect 22051 17629 22063 17663
rect 22005 17623 22063 17629
rect 22189 17663 22247 17669
rect 22189 17629 22201 17663
rect 22235 17629 22247 17663
rect 22189 17623 22247 17629
rect 22370 17620 22376 17672
rect 22428 17620 22434 17672
rect 22922 17620 22928 17672
rect 22980 17620 22986 17672
rect 23198 17620 23204 17672
rect 23256 17620 23262 17672
rect 23290 17620 23296 17672
rect 23348 17620 23354 17672
rect 23492 17669 23520 17700
rect 23584 17700 24041 17728
rect 23584 17672 23612 17700
rect 24029 17697 24041 17700
rect 24075 17697 24087 17731
rect 24029 17691 24087 17697
rect 23477 17663 23535 17669
rect 23477 17629 23489 17663
rect 23523 17629 23535 17663
rect 23477 17623 23535 17629
rect 23566 17620 23572 17672
rect 23624 17620 23630 17672
rect 23661 17663 23719 17669
rect 23661 17629 23673 17663
rect 23707 17660 23719 17663
rect 23753 17663 23811 17669
rect 23753 17660 23765 17663
rect 23707 17632 23765 17660
rect 23707 17629 23719 17632
rect 23661 17623 23719 17629
rect 23753 17629 23765 17632
rect 23799 17629 23811 17663
rect 23753 17623 23811 17629
rect 24302 17620 24308 17672
rect 24360 17660 24366 17672
rect 24670 17669 24676 17672
rect 24397 17663 24455 17669
rect 24397 17660 24409 17663
rect 24360 17632 24409 17660
rect 24360 17620 24366 17632
rect 24397 17629 24409 17632
rect 24443 17629 24455 17663
rect 24664 17660 24676 17669
rect 24631 17632 24676 17660
rect 24397 17623 24455 17629
rect 24664 17623 24676 17632
rect 22097 17595 22155 17601
rect 22097 17561 22109 17595
rect 22143 17592 22155 17595
rect 22465 17595 22523 17601
rect 22465 17592 22477 17595
rect 22143 17564 22477 17592
rect 22143 17561 22155 17564
rect 22097 17555 22155 17561
rect 22465 17561 22477 17564
rect 22511 17561 22523 17595
rect 22465 17555 22523 17561
rect 22649 17595 22707 17601
rect 22649 17561 22661 17595
rect 22695 17592 22707 17595
rect 23216 17592 23244 17620
rect 22695 17564 23244 17592
rect 24412 17592 24440 17623
rect 24670 17620 24676 17623
rect 24728 17620 24734 17672
rect 25869 17663 25927 17669
rect 25869 17629 25881 17663
rect 25915 17629 25927 17663
rect 25869 17623 25927 17629
rect 25038 17592 25044 17604
rect 24412 17564 25044 17592
rect 22695 17561 22707 17564
rect 22649 17555 22707 17561
rect 25038 17552 25044 17564
rect 25096 17592 25102 17604
rect 25884 17592 25912 17623
rect 27890 17620 27896 17672
rect 27948 17660 27954 17672
rect 28454 17663 28512 17669
rect 28454 17660 28466 17663
rect 27948 17632 28466 17660
rect 27948 17620 27954 17632
rect 28454 17629 28466 17632
rect 28500 17629 28512 17663
rect 28721 17663 28779 17669
rect 28721 17660 28733 17663
rect 28454 17623 28512 17629
rect 28552 17632 28733 17660
rect 25096 17564 25912 17592
rect 25096 17552 25102 17564
rect 25958 17552 25964 17604
rect 26016 17592 26022 17604
rect 26114 17595 26172 17601
rect 26114 17592 26126 17595
rect 26016 17564 26126 17592
rect 26016 17552 26022 17564
rect 26114 17561 26126 17564
rect 26160 17561 26172 17595
rect 26114 17555 26172 17561
rect 28552 17536 28580 17632
rect 28721 17629 28733 17632
rect 28767 17629 28779 17663
rect 28721 17623 28779 17629
rect 29641 17663 29699 17669
rect 29641 17629 29653 17663
rect 29687 17660 29699 17663
rect 30300 17660 30328 17756
rect 29687 17632 30328 17660
rect 29687 17629 29699 17632
rect 29641 17623 29699 17629
rect 31386 17620 31392 17672
rect 31444 17660 31450 17672
rect 31481 17663 31539 17669
rect 31481 17660 31493 17663
rect 31444 17632 31493 17660
rect 31444 17620 31450 17632
rect 31481 17629 31493 17632
rect 31527 17629 31539 17663
rect 31481 17623 31539 17629
rect 30834 17552 30840 17604
rect 30892 17592 30898 17604
rect 31214 17595 31272 17601
rect 31214 17592 31226 17595
rect 30892 17564 31226 17592
rect 30892 17552 30898 17564
rect 31214 17561 31226 17564
rect 31260 17561 31272 17595
rect 31214 17555 31272 17561
rect 20640 17496 21404 17524
rect 21450 17484 21456 17536
rect 21508 17484 21514 17536
rect 21818 17484 21824 17536
rect 21876 17484 21882 17536
rect 22278 17484 22284 17536
rect 22336 17484 22342 17536
rect 22738 17484 22744 17536
rect 22796 17484 22802 17536
rect 27246 17484 27252 17536
rect 27304 17484 27310 17536
rect 27338 17484 27344 17536
rect 27396 17484 27402 17536
rect 28534 17484 28540 17536
rect 28592 17484 28598 17536
rect 1104 17434 35027 17456
rect 1104 17382 9390 17434
rect 9442 17382 9454 17434
rect 9506 17382 9518 17434
rect 9570 17382 9582 17434
rect 9634 17382 9646 17434
rect 9698 17382 17831 17434
rect 17883 17382 17895 17434
rect 17947 17382 17959 17434
rect 18011 17382 18023 17434
rect 18075 17382 18087 17434
rect 18139 17382 26272 17434
rect 26324 17382 26336 17434
rect 26388 17382 26400 17434
rect 26452 17382 26464 17434
rect 26516 17382 26528 17434
rect 26580 17382 34713 17434
rect 34765 17382 34777 17434
rect 34829 17382 34841 17434
rect 34893 17382 34905 17434
rect 34957 17382 34969 17434
rect 35021 17382 35027 17434
rect 1104 17360 35027 17382
rect 15562 17280 15568 17332
rect 15620 17280 15626 17332
rect 16114 17280 16120 17332
rect 16172 17320 16178 17332
rect 16209 17323 16267 17329
rect 16209 17320 16221 17323
rect 16172 17292 16221 17320
rect 16172 17280 16178 17292
rect 16209 17289 16221 17292
rect 16255 17289 16267 17323
rect 16209 17283 16267 17289
rect 17126 17280 17132 17332
rect 17184 17280 17190 17332
rect 18049 17323 18107 17329
rect 18049 17289 18061 17323
rect 18095 17320 18107 17323
rect 18230 17320 18236 17332
rect 18095 17292 18236 17320
rect 18095 17289 18107 17292
rect 18049 17283 18107 17289
rect 18230 17280 18236 17292
rect 18288 17320 18294 17332
rect 18288 17292 18736 17320
rect 18288 17280 18294 17292
rect 15580 17193 15608 17280
rect 16022 17212 16028 17264
rect 16080 17252 16086 17264
rect 16936 17255 16994 17261
rect 16080 17224 16160 17252
rect 16080 17212 16086 17224
rect 16132 17193 16160 17224
rect 16936 17221 16948 17255
rect 16982 17252 16994 17255
rect 17144 17252 17172 17280
rect 16982 17224 17172 17252
rect 16982 17221 16994 17224
rect 16936 17215 16994 17221
rect 18506 17212 18512 17264
rect 18564 17252 18570 17264
rect 18564 17224 18644 17252
rect 18564 17212 18570 17224
rect 15565 17187 15623 17193
rect 15565 17153 15577 17187
rect 15611 17153 15623 17187
rect 15565 17147 15623 17153
rect 16117 17187 16175 17193
rect 16117 17153 16129 17187
rect 16163 17153 16175 17187
rect 16117 17147 16175 17153
rect 16206 17144 16212 17196
rect 16264 17184 16270 17196
rect 18414 17193 18420 17196
rect 16669 17187 16727 17193
rect 16669 17184 16681 17187
rect 16264 17156 16681 17184
rect 16264 17144 16270 17156
rect 16669 17153 16681 17156
rect 16715 17153 16727 17187
rect 16669 17147 16727 17153
rect 18141 17187 18199 17193
rect 18141 17153 18153 17187
rect 18187 17153 18199 17187
rect 18141 17147 18199 17153
rect 18325 17187 18383 17193
rect 18325 17153 18337 17187
rect 18371 17153 18383 17187
rect 18325 17147 18383 17153
rect 18413 17147 18420 17193
rect 18472 17184 18478 17196
rect 18616 17193 18644 17224
rect 18601 17187 18659 17193
rect 18472 17156 18513 17184
rect 18156 17048 18184 17147
rect 18340 17116 18368 17147
rect 18414 17144 18420 17147
rect 18472 17144 18478 17156
rect 18601 17153 18613 17187
rect 18647 17153 18659 17187
rect 18708 17184 18736 17292
rect 18782 17280 18788 17332
rect 18840 17280 18846 17332
rect 19978 17280 19984 17332
rect 20036 17320 20042 17332
rect 20165 17323 20223 17329
rect 20165 17320 20177 17323
rect 20036 17292 20177 17320
rect 20036 17280 20042 17292
rect 20165 17289 20177 17292
rect 20211 17289 20223 17323
rect 20165 17283 20223 17289
rect 20254 17280 20260 17332
rect 20312 17280 20318 17332
rect 20346 17280 20352 17332
rect 20404 17280 20410 17332
rect 20806 17280 20812 17332
rect 20864 17280 20870 17332
rect 20916 17292 22692 17320
rect 18800 17252 18828 17280
rect 18800 17224 20024 17252
rect 18892 17193 18920 17224
rect 18785 17187 18843 17193
rect 18785 17184 18797 17187
rect 18708 17156 18797 17184
rect 18601 17147 18659 17153
rect 18785 17153 18797 17156
rect 18831 17153 18843 17187
rect 18785 17147 18843 17153
rect 18877 17187 18935 17193
rect 18877 17153 18889 17187
rect 18923 17153 18935 17187
rect 18877 17147 18935 17153
rect 19153 17187 19211 17193
rect 19153 17153 19165 17187
rect 19199 17184 19211 17187
rect 19426 17184 19432 17196
rect 19199 17156 19432 17184
rect 19199 17153 19211 17156
rect 19153 17147 19211 17153
rect 19426 17144 19432 17156
rect 19484 17144 19490 17196
rect 19702 17144 19708 17196
rect 19760 17144 19766 17196
rect 19797 17187 19855 17193
rect 19797 17153 19809 17187
rect 19843 17184 19855 17187
rect 19996 17184 20024 17224
rect 20070 17184 20076 17196
rect 19843 17156 19932 17184
rect 19996 17156 20076 17184
rect 19843 17153 19855 17156
rect 19797 17147 19855 17153
rect 18966 17116 18972 17128
rect 18340 17088 18972 17116
rect 18966 17076 18972 17088
rect 19024 17076 19030 17128
rect 19904 17048 19932 17156
rect 20070 17144 20076 17156
rect 20128 17144 20134 17196
rect 19981 17119 20039 17125
rect 19981 17085 19993 17119
rect 20027 17116 20039 17119
rect 20272 17116 20300 17280
rect 20364 17252 20392 17280
rect 20364 17224 20668 17252
rect 20349 17187 20407 17193
rect 20349 17153 20361 17187
rect 20395 17184 20407 17187
rect 20438 17184 20444 17196
rect 20395 17156 20444 17184
rect 20395 17153 20407 17156
rect 20349 17147 20407 17153
rect 20438 17144 20444 17156
rect 20496 17144 20502 17196
rect 20530 17144 20536 17196
rect 20588 17144 20594 17196
rect 20640 17193 20668 17224
rect 20625 17187 20683 17193
rect 20625 17153 20637 17187
rect 20671 17153 20683 17187
rect 20625 17147 20683 17153
rect 20717 17187 20775 17193
rect 20717 17153 20729 17187
rect 20763 17184 20775 17187
rect 20824 17184 20852 17280
rect 20916 17193 20944 17292
rect 21008 17224 22140 17252
rect 20763 17156 20852 17184
rect 20901 17187 20959 17193
rect 20763 17153 20775 17156
rect 20717 17147 20775 17153
rect 20901 17153 20913 17187
rect 20947 17153 20959 17187
rect 20901 17147 20959 17153
rect 20027 17088 20300 17116
rect 20548 17116 20576 17144
rect 21008 17116 21036 17224
rect 21177 17187 21235 17193
rect 21177 17153 21189 17187
rect 21223 17184 21235 17187
rect 21818 17184 21824 17196
rect 21223 17156 21824 17184
rect 21223 17153 21235 17156
rect 21177 17147 21235 17153
rect 21818 17144 21824 17156
rect 21876 17184 21882 17196
rect 22005 17187 22063 17193
rect 22005 17184 22017 17187
rect 21876 17156 22017 17184
rect 21876 17144 21882 17156
rect 22005 17153 22017 17156
rect 22051 17153 22063 17187
rect 22005 17147 22063 17153
rect 20548 17088 21036 17116
rect 21269 17119 21327 17125
rect 20027 17085 20039 17088
rect 19981 17079 20039 17085
rect 21269 17085 21281 17119
rect 21315 17085 21327 17119
rect 21269 17079 21327 17085
rect 20993 17051 21051 17057
rect 20993 17048 21005 17051
rect 18156 17020 19840 17048
rect 19904 17020 21005 17048
rect 18141 16983 18199 16989
rect 18141 16949 18153 16983
rect 18187 16980 18199 16983
rect 18230 16980 18236 16992
rect 18187 16952 18236 16980
rect 18187 16949 18199 16952
rect 18141 16943 18199 16949
rect 18230 16940 18236 16952
rect 18288 16940 18294 16992
rect 19334 16940 19340 16992
rect 19392 16940 19398 16992
rect 19521 16983 19579 16989
rect 19521 16949 19533 16983
rect 19567 16980 19579 16983
rect 19702 16980 19708 16992
rect 19567 16952 19708 16980
rect 19567 16949 19579 16952
rect 19521 16943 19579 16949
rect 19702 16940 19708 16952
rect 19760 16940 19766 16992
rect 19812 16980 19840 17020
rect 20993 17017 21005 17020
rect 21039 17017 21051 17051
rect 21284 17048 21312 17079
rect 21634 17076 21640 17128
rect 21692 17116 21698 17128
rect 22112 17116 22140 17224
rect 22204 17224 22416 17252
rect 22204 17193 22232 17224
rect 22388 17196 22416 17224
rect 22189 17187 22247 17193
rect 22189 17153 22201 17187
rect 22235 17153 22247 17187
rect 22189 17147 22247 17153
rect 22278 17144 22284 17196
rect 22336 17144 22342 17196
rect 22370 17144 22376 17196
rect 22428 17144 22434 17196
rect 22462 17144 22468 17196
rect 22520 17144 22526 17196
rect 22664 17184 22692 17292
rect 22738 17280 22744 17332
rect 22796 17280 22802 17332
rect 22830 17280 22836 17332
rect 22888 17320 22894 17332
rect 24394 17320 24400 17332
rect 22888 17292 24400 17320
rect 22888 17280 22894 17292
rect 24394 17280 24400 17292
rect 24452 17280 24458 17332
rect 24946 17280 24952 17332
rect 25004 17320 25010 17332
rect 25041 17323 25099 17329
rect 25041 17320 25053 17323
rect 25004 17292 25053 17320
rect 25004 17280 25010 17292
rect 25041 17289 25053 17292
rect 25087 17289 25099 17323
rect 25041 17283 25099 17289
rect 25590 17280 25596 17332
rect 25648 17280 25654 17332
rect 25777 17323 25835 17329
rect 25777 17289 25789 17323
rect 25823 17289 25835 17323
rect 25777 17283 25835 17289
rect 22756 17252 22784 17280
rect 23566 17252 23572 17264
rect 22756 17224 22968 17252
rect 22741 17187 22799 17193
rect 22741 17184 22753 17187
rect 22664 17156 22753 17184
rect 22741 17153 22753 17156
rect 22787 17184 22799 17187
rect 22830 17184 22836 17196
rect 22787 17156 22836 17184
rect 22787 17153 22799 17156
rect 22741 17147 22799 17153
rect 22830 17144 22836 17156
rect 22888 17144 22894 17196
rect 22940 17193 22968 17224
rect 23124 17224 23572 17252
rect 22925 17187 22983 17193
rect 22925 17153 22937 17187
rect 22971 17153 22983 17187
rect 22925 17147 22983 17153
rect 23014 17144 23020 17196
rect 23072 17144 23078 17196
rect 23124 17125 23152 17224
rect 23566 17212 23572 17224
rect 23624 17212 23630 17264
rect 25608 17252 25636 17280
rect 25240 17224 25636 17252
rect 25792 17252 25820 17283
rect 25866 17280 25872 17332
rect 25924 17280 25930 17332
rect 25958 17280 25964 17332
rect 26016 17280 26022 17332
rect 26142 17280 26148 17332
rect 26200 17280 26206 17332
rect 26602 17280 26608 17332
rect 26660 17280 26666 17332
rect 26970 17280 26976 17332
rect 27028 17280 27034 17332
rect 27246 17280 27252 17332
rect 27304 17280 27310 17332
rect 29270 17280 29276 17332
rect 29328 17280 29334 17332
rect 29546 17280 29552 17332
rect 29604 17280 29610 17332
rect 29638 17280 29644 17332
rect 29696 17280 29702 17332
rect 29730 17280 29736 17332
rect 29788 17280 29794 17332
rect 30834 17280 30840 17332
rect 30892 17280 30898 17332
rect 25976 17252 26004 17280
rect 26160 17252 26188 17280
rect 25792 17224 26004 17252
rect 26068 17224 26188 17252
rect 26620 17252 26648 17280
rect 26620 17224 27200 17252
rect 25240 17196 25268 17224
rect 23293 17187 23351 17193
rect 23293 17153 23305 17187
rect 23339 17184 23351 17187
rect 23382 17184 23388 17196
rect 23339 17156 23388 17184
rect 23339 17153 23351 17156
rect 23293 17147 23351 17153
rect 23382 17144 23388 17156
rect 23440 17144 23446 17196
rect 23477 17187 23535 17193
rect 23477 17153 23489 17187
rect 23523 17184 23535 17187
rect 24682 17187 24740 17193
rect 24682 17184 24694 17187
rect 23523 17156 24694 17184
rect 23523 17153 23535 17156
rect 23477 17147 23535 17153
rect 24682 17153 24694 17156
rect 24728 17153 24740 17187
rect 24682 17147 24740 17153
rect 24854 17144 24860 17196
rect 24912 17184 24918 17196
rect 24949 17187 25007 17193
rect 24949 17184 24961 17187
rect 24912 17156 24961 17184
rect 24912 17144 24918 17156
rect 24949 17153 24961 17156
rect 24995 17153 25007 17187
rect 24949 17147 25007 17153
rect 25222 17144 25228 17196
rect 25280 17144 25286 17196
rect 25593 17187 25651 17193
rect 25593 17153 25605 17187
rect 25639 17184 25651 17187
rect 26068 17184 26096 17224
rect 25639 17156 26096 17184
rect 25639 17153 25651 17156
rect 25593 17147 25651 17153
rect 26142 17144 26148 17196
rect 26200 17144 26206 17196
rect 26234 17144 26240 17196
rect 26292 17184 26298 17196
rect 26605 17187 26663 17193
rect 26605 17184 26617 17187
rect 26292 17156 26617 17184
rect 26292 17144 26298 17156
rect 26605 17153 26617 17156
rect 26651 17184 26663 17187
rect 26970 17184 26976 17196
rect 26651 17156 26976 17184
rect 26651 17153 26663 17156
rect 26605 17147 26663 17153
rect 26970 17144 26976 17156
rect 27028 17144 27034 17196
rect 27172 17193 27200 17224
rect 27264 17193 27292 17280
rect 27157 17187 27215 17193
rect 27157 17153 27169 17187
rect 27203 17153 27215 17187
rect 27157 17147 27215 17153
rect 27249 17187 27307 17193
rect 27249 17153 27261 17187
rect 27295 17153 27307 17187
rect 27249 17147 27307 17153
rect 29457 17187 29515 17193
rect 29457 17153 29469 17187
rect 29503 17184 29515 17187
rect 29564 17184 29592 17280
rect 29656 17252 29684 17280
rect 29825 17255 29883 17261
rect 29825 17252 29837 17255
rect 29656 17224 29837 17252
rect 29825 17221 29837 17224
rect 29871 17221 29883 17255
rect 29825 17215 29883 17221
rect 29503 17156 29592 17184
rect 29503 17153 29515 17156
rect 29457 17147 29515 17153
rect 23109 17119 23167 17125
rect 23109 17116 23121 17119
rect 21692 17088 21864 17116
rect 22112 17088 23121 17116
rect 21692 17076 21698 17088
rect 21284 17020 21772 17048
rect 20993 17011 21051 17017
rect 21744 16992 21772 17020
rect 21082 16980 21088 16992
rect 19812 16952 21088 16980
rect 21082 16940 21088 16952
rect 21140 16940 21146 16992
rect 21726 16940 21732 16992
rect 21784 16940 21790 16992
rect 21836 16980 21864 17088
rect 23109 17085 23121 17088
rect 23155 17085 23167 17119
rect 23109 17079 23167 17085
rect 22370 17008 22376 17060
rect 22428 17048 22434 17060
rect 22922 17048 22928 17060
rect 22428 17020 22928 17048
rect 22428 17008 22434 17020
rect 22922 17008 22928 17020
rect 22980 17008 22986 17060
rect 23400 17048 23428 17144
rect 25409 17119 25467 17125
rect 25409 17085 25421 17119
rect 25455 17116 25467 17119
rect 26252 17116 26280 17144
rect 25455 17088 26280 17116
rect 26329 17119 26387 17125
rect 25455 17085 25467 17088
rect 25409 17079 25467 17085
rect 26329 17085 26341 17119
rect 26375 17116 26387 17119
rect 26418 17116 26424 17128
rect 26375 17088 26424 17116
rect 26375 17085 26387 17088
rect 26329 17079 26387 17085
rect 26418 17076 26424 17088
rect 26476 17116 26482 17128
rect 27264 17116 27292 17147
rect 30374 17144 30380 17196
rect 30432 17184 30438 17196
rect 30653 17187 30711 17193
rect 30653 17184 30665 17187
rect 30432 17156 30665 17184
rect 30432 17144 30438 17156
rect 30653 17153 30665 17156
rect 30699 17153 30711 17187
rect 30653 17147 30711 17153
rect 29549 17119 29607 17125
rect 29549 17116 29561 17119
rect 26476 17088 27292 17116
rect 29472 17088 29561 17116
rect 26476 17076 26482 17088
rect 29472 17060 29500 17088
rect 29549 17085 29561 17088
rect 29595 17085 29607 17119
rect 29549 17079 29607 17085
rect 29914 17076 29920 17128
rect 29972 17076 29978 17128
rect 23569 17051 23627 17057
rect 23569 17048 23581 17051
rect 23400 17020 23581 17048
rect 23569 17017 23581 17020
rect 23615 17017 23627 17051
rect 23569 17011 23627 17017
rect 25682 17008 25688 17060
rect 25740 17048 25746 17060
rect 26142 17048 26148 17060
rect 25740 17020 26148 17048
rect 25740 17008 25746 17020
rect 26142 17008 26148 17020
rect 26200 17008 26206 17060
rect 26237 17051 26295 17057
rect 26237 17017 26249 17051
rect 26283 17048 26295 17051
rect 26694 17048 26700 17060
rect 26283 17020 26700 17048
rect 26283 17017 26295 17020
rect 26237 17011 26295 17017
rect 26694 17008 26700 17020
rect 26752 17008 26758 17060
rect 29454 17008 29460 17060
rect 29512 17008 29518 17060
rect 22830 16980 22836 16992
rect 21836 16952 22836 16980
rect 22830 16940 22836 16952
rect 22888 16940 22894 16992
rect 26326 16940 26332 16992
rect 26384 16980 26390 16992
rect 26421 16983 26479 16989
rect 26421 16980 26433 16983
rect 26384 16952 26433 16980
rect 26384 16940 26390 16952
rect 26421 16949 26433 16952
rect 26467 16980 26479 16983
rect 27338 16980 27344 16992
rect 26467 16952 27344 16980
rect 26467 16949 26479 16952
rect 26421 16943 26479 16949
rect 27338 16940 27344 16952
rect 27396 16940 27402 16992
rect 1104 16890 34868 16912
rect 1104 16838 5170 16890
rect 5222 16838 5234 16890
rect 5286 16838 5298 16890
rect 5350 16838 5362 16890
rect 5414 16838 5426 16890
rect 5478 16838 13611 16890
rect 13663 16838 13675 16890
rect 13727 16838 13739 16890
rect 13791 16838 13803 16890
rect 13855 16838 13867 16890
rect 13919 16838 22052 16890
rect 22104 16838 22116 16890
rect 22168 16838 22180 16890
rect 22232 16838 22244 16890
rect 22296 16838 22308 16890
rect 22360 16838 30493 16890
rect 30545 16838 30557 16890
rect 30609 16838 30621 16890
rect 30673 16838 30685 16890
rect 30737 16838 30749 16890
rect 30801 16838 34868 16890
rect 1104 16816 34868 16838
rect 18877 16779 18935 16785
rect 18877 16745 18889 16779
rect 18923 16776 18935 16779
rect 18966 16776 18972 16788
rect 18923 16748 18972 16776
rect 18923 16745 18935 16748
rect 18877 16739 18935 16745
rect 18966 16736 18972 16748
rect 19024 16736 19030 16788
rect 19334 16736 19340 16788
rect 19392 16776 19398 16788
rect 19521 16779 19579 16785
rect 19521 16776 19533 16779
rect 19392 16748 19533 16776
rect 19392 16736 19398 16748
rect 19521 16745 19533 16748
rect 19567 16745 19579 16779
rect 19521 16739 19579 16745
rect 19886 16736 19892 16788
rect 19944 16736 19950 16788
rect 20717 16779 20775 16785
rect 20717 16745 20729 16779
rect 20763 16776 20775 16779
rect 20990 16776 20996 16788
rect 20763 16748 20996 16776
rect 20763 16745 20775 16748
rect 20717 16739 20775 16745
rect 20990 16736 20996 16748
rect 21048 16736 21054 16788
rect 21726 16736 21732 16788
rect 21784 16736 21790 16788
rect 21818 16736 21824 16788
rect 21876 16776 21882 16788
rect 22281 16779 22339 16785
rect 21876 16748 22094 16776
rect 21876 16736 21882 16748
rect 16206 16600 16212 16652
rect 16264 16640 16270 16652
rect 17497 16643 17555 16649
rect 17497 16640 17509 16643
rect 16264 16612 17509 16640
rect 16264 16600 16270 16612
rect 17497 16609 17509 16612
rect 17543 16640 17555 16643
rect 17543 16612 17632 16640
rect 17543 16609 17555 16612
rect 17497 16603 17555 16609
rect 17604 16572 17632 16612
rect 18506 16572 18512 16584
rect 17604 16544 18512 16572
rect 18506 16532 18512 16544
rect 18564 16532 18570 16584
rect 18984 16572 19012 16736
rect 19904 16708 19932 16736
rect 19628 16680 19932 16708
rect 19628 16649 19656 16680
rect 19613 16643 19671 16649
rect 19613 16609 19625 16643
rect 19659 16609 19671 16643
rect 19613 16603 19671 16609
rect 19702 16600 19708 16652
rect 19760 16640 19766 16652
rect 19904 16640 19932 16680
rect 20898 16668 20904 16720
rect 20956 16668 20962 16720
rect 22066 16708 22094 16748
rect 22281 16745 22293 16779
rect 22327 16776 22339 16779
rect 22370 16776 22376 16788
rect 22327 16748 22376 16776
rect 22327 16745 22339 16748
rect 22281 16739 22339 16745
rect 22370 16736 22376 16748
rect 22428 16736 22434 16788
rect 22462 16736 22468 16788
rect 22520 16776 22526 16788
rect 22557 16779 22615 16785
rect 22557 16776 22569 16779
rect 22520 16748 22569 16776
rect 22520 16736 22526 16748
rect 22557 16745 22569 16748
rect 22603 16745 22615 16779
rect 22557 16739 22615 16745
rect 22925 16779 22983 16785
rect 22925 16745 22937 16779
rect 22971 16776 22983 16779
rect 23014 16776 23020 16788
rect 22971 16748 23020 16776
rect 22971 16745 22983 16748
rect 22925 16739 22983 16745
rect 23014 16736 23020 16748
rect 23072 16736 23078 16788
rect 23198 16736 23204 16788
rect 23256 16776 23262 16788
rect 23385 16779 23443 16785
rect 23385 16776 23397 16779
rect 23256 16748 23397 16776
rect 23256 16736 23262 16748
rect 23385 16745 23397 16748
rect 23431 16745 23443 16779
rect 23385 16739 23443 16745
rect 25869 16779 25927 16785
rect 25869 16745 25881 16779
rect 25915 16776 25927 16779
rect 26050 16776 26056 16788
rect 25915 16748 26056 16776
rect 25915 16745 25927 16748
rect 25869 16739 25927 16745
rect 26050 16736 26056 16748
rect 26108 16736 26114 16788
rect 26142 16736 26148 16788
rect 26200 16736 26206 16788
rect 26418 16736 26424 16788
rect 26476 16736 26482 16788
rect 29362 16736 29368 16788
rect 29420 16776 29426 16788
rect 29420 16748 29776 16776
rect 29420 16736 29426 16748
rect 22649 16711 22707 16717
rect 22649 16708 22661 16711
rect 22066 16680 22661 16708
rect 22649 16677 22661 16680
rect 22695 16677 22707 16711
rect 26160 16708 26188 16736
rect 22649 16671 22707 16677
rect 22756 16680 23612 16708
rect 20533 16643 20591 16649
rect 19760 16612 19840 16640
rect 19904 16612 20024 16640
rect 19760 16600 19766 16612
rect 19812 16581 19840 16612
rect 19996 16581 20024 16612
rect 20533 16609 20545 16643
rect 20579 16640 20591 16643
rect 22097 16643 22155 16649
rect 22097 16640 22109 16643
rect 20579 16612 22109 16640
rect 20579 16609 20591 16612
rect 20533 16603 20591 16609
rect 19245 16575 19303 16581
rect 19245 16572 19257 16575
rect 18984 16544 19257 16572
rect 19245 16541 19257 16544
rect 19291 16541 19303 16575
rect 19245 16535 19303 16541
rect 19797 16575 19855 16581
rect 19797 16541 19809 16575
rect 19843 16541 19855 16575
rect 19797 16535 19855 16541
rect 19981 16575 20039 16581
rect 19981 16541 19993 16575
rect 20027 16541 20039 16575
rect 19981 16535 20039 16541
rect 20438 16532 20444 16584
rect 20496 16572 20502 16584
rect 20622 16572 20628 16584
rect 20496 16544 20628 16572
rect 20496 16532 20502 16544
rect 20622 16532 20628 16544
rect 20680 16532 20686 16584
rect 21100 16581 21128 16612
rect 22097 16609 22109 16612
rect 22143 16640 22155 16643
rect 22465 16643 22523 16649
rect 22465 16640 22477 16643
rect 22143 16612 22477 16640
rect 22143 16609 22155 16612
rect 22097 16603 22155 16609
rect 22465 16609 22477 16612
rect 22511 16640 22523 16643
rect 22554 16640 22560 16652
rect 22511 16612 22560 16640
rect 22511 16609 22523 16612
rect 22465 16603 22523 16609
rect 22554 16600 22560 16612
rect 22612 16640 22618 16652
rect 22756 16640 22784 16680
rect 22612 16612 22784 16640
rect 22612 16600 22618 16612
rect 21085 16575 21143 16581
rect 21085 16541 21097 16575
rect 21131 16541 21143 16575
rect 21085 16535 21143 16541
rect 21177 16575 21235 16581
rect 21177 16541 21189 16575
rect 21223 16541 21235 16575
rect 21177 16535 21235 16541
rect 21361 16575 21419 16581
rect 21361 16541 21373 16575
rect 21407 16541 21419 16575
rect 21361 16535 21419 16541
rect 17764 16507 17822 16513
rect 17764 16473 17776 16507
rect 17810 16473 17822 16507
rect 17764 16467 17822 16473
rect 17678 16396 17684 16448
rect 17736 16436 17742 16448
rect 17788 16436 17816 16467
rect 19702 16464 19708 16516
rect 19760 16464 19766 16516
rect 21192 16504 21220 16535
rect 21008 16476 21220 16504
rect 17736 16408 17816 16436
rect 19337 16439 19395 16445
rect 17736 16396 17742 16408
rect 19337 16405 19349 16439
rect 19383 16436 19395 16439
rect 19426 16436 19432 16448
rect 19383 16408 19432 16436
rect 19383 16405 19395 16408
rect 19337 16399 19395 16405
rect 19426 16396 19432 16408
rect 19484 16396 19490 16448
rect 19886 16396 19892 16448
rect 19944 16396 19950 16448
rect 20162 16396 20168 16448
rect 20220 16436 20226 16448
rect 21008 16436 21036 16476
rect 20220 16408 21036 16436
rect 20220 16396 20226 16408
rect 21082 16396 21088 16448
rect 21140 16436 21146 16448
rect 21376 16436 21404 16535
rect 21450 16532 21456 16584
rect 21508 16572 21514 16584
rect 21545 16575 21603 16581
rect 21545 16572 21557 16575
rect 21508 16544 21557 16572
rect 21508 16532 21514 16544
rect 21545 16541 21557 16544
rect 21591 16541 21603 16575
rect 21545 16535 21603 16541
rect 22005 16575 22063 16581
rect 22005 16541 22017 16575
rect 22051 16572 22063 16575
rect 22741 16575 22799 16581
rect 22051 16544 22085 16572
rect 22051 16541 22063 16544
rect 22005 16535 22063 16541
rect 22741 16541 22753 16575
rect 22787 16541 22799 16575
rect 22741 16535 22799 16541
rect 21910 16464 21916 16516
rect 21968 16504 21974 16516
rect 22020 16504 22048 16535
rect 22756 16504 22784 16535
rect 22830 16532 22836 16584
rect 22888 16532 22894 16584
rect 22922 16532 22928 16584
rect 22980 16572 22986 16584
rect 23017 16575 23075 16581
rect 23017 16572 23029 16575
rect 22980 16544 23029 16572
rect 22980 16532 22986 16544
rect 23017 16541 23029 16544
rect 23063 16541 23075 16575
rect 23017 16535 23075 16541
rect 23106 16532 23112 16584
rect 23164 16581 23170 16584
rect 23164 16575 23213 16581
rect 23164 16541 23167 16575
rect 23201 16541 23213 16575
rect 23164 16535 23213 16541
rect 23164 16532 23170 16535
rect 23290 16532 23296 16584
rect 23348 16532 23354 16584
rect 23584 16581 23612 16680
rect 26068 16680 26188 16708
rect 23658 16600 23664 16652
rect 23716 16640 23722 16652
rect 26068 16649 26096 16680
rect 26234 16668 26240 16720
rect 26292 16668 26298 16720
rect 23753 16643 23811 16649
rect 23753 16640 23765 16643
rect 23716 16612 23765 16640
rect 23716 16600 23722 16612
rect 23753 16609 23765 16612
rect 23799 16609 23811 16643
rect 23753 16603 23811 16609
rect 26053 16643 26111 16649
rect 26053 16609 26065 16643
rect 26099 16609 26111 16643
rect 26053 16603 26111 16609
rect 26145 16643 26203 16649
rect 26145 16609 26157 16643
rect 26191 16640 26203 16643
rect 26252 16640 26280 16668
rect 26436 16649 26464 16736
rect 26191 16612 26280 16640
rect 26421 16643 26479 16649
rect 26191 16609 26203 16612
rect 26145 16603 26203 16609
rect 26421 16609 26433 16643
rect 26467 16609 26479 16643
rect 29549 16643 29607 16649
rect 29549 16640 29561 16643
rect 26421 16603 26479 16609
rect 29104 16612 29561 16640
rect 29104 16584 29132 16612
rect 29549 16609 29561 16612
rect 29595 16609 29607 16643
rect 29549 16603 29607 16609
rect 23569 16575 23627 16581
rect 23569 16541 23581 16575
rect 23615 16541 23627 16575
rect 23569 16535 23627 16541
rect 26234 16532 26240 16584
rect 26292 16572 26298 16584
rect 26513 16575 26571 16581
rect 26513 16572 26525 16575
rect 26292 16544 26525 16572
rect 26292 16532 26298 16544
rect 26513 16541 26525 16544
rect 26559 16541 26571 16575
rect 26513 16535 26571 16541
rect 26602 16532 26608 16584
rect 26660 16532 26666 16584
rect 28258 16532 28264 16584
rect 28316 16532 28322 16584
rect 29086 16532 29092 16584
rect 29144 16532 29150 16584
rect 29748 16581 29776 16748
rect 29914 16736 29920 16788
rect 29972 16776 29978 16788
rect 30101 16779 30159 16785
rect 30101 16776 30113 16779
rect 29972 16748 30113 16776
rect 29972 16736 29978 16748
rect 30101 16745 30113 16748
rect 30147 16745 30159 16779
rect 30101 16739 30159 16745
rect 30374 16736 30380 16788
rect 30432 16736 30438 16788
rect 30926 16776 30932 16788
rect 30668 16748 30932 16776
rect 30392 16708 30420 16736
rect 30561 16711 30619 16717
rect 30561 16708 30573 16711
rect 30392 16680 30573 16708
rect 30561 16677 30573 16680
rect 30607 16677 30619 16711
rect 30561 16671 30619 16677
rect 30668 16640 30696 16748
rect 30926 16736 30932 16748
rect 30984 16736 30990 16788
rect 30392 16612 30696 16640
rect 30392 16584 30420 16612
rect 29181 16575 29239 16581
rect 29181 16541 29193 16575
rect 29227 16572 29239 16575
rect 29733 16575 29791 16581
rect 29227 16544 29684 16572
rect 29227 16541 29239 16544
rect 29181 16535 29239 16541
rect 23382 16504 23388 16516
rect 21968 16476 23388 16504
rect 21968 16464 21974 16476
rect 23382 16464 23388 16476
rect 23440 16464 23446 16516
rect 26326 16464 26332 16516
rect 26384 16464 26390 16516
rect 29365 16507 29423 16513
rect 29365 16473 29377 16507
rect 29411 16473 29423 16507
rect 29656 16504 29684 16544
rect 29733 16541 29745 16575
rect 29779 16541 29791 16575
rect 29733 16535 29791 16541
rect 29825 16575 29883 16581
rect 29825 16541 29837 16575
rect 29871 16572 29883 16575
rect 30193 16575 30251 16581
rect 30193 16572 30205 16575
rect 29871 16544 30205 16572
rect 29871 16541 29883 16544
rect 29825 16535 29883 16541
rect 30024 16504 30052 16544
rect 30193 16541 30205 16544
rect 30239 16541 30251 16575
rect 30193 16535 30251 16541
rect 30374 16532 30380 16584
rect 30432 16532 30438 16584
rect 30650 16532 30656 16584
rect 30708 16572 30714 16584
rect 30745 16575 30803 16581
rect 30745 16572 30757 16575
rect 30708 16544 30757 16572
rect 30708 16532 30714 16544
rect 30745 16541 30757 16544
rect 30791 16572 30803 16575
rect 31386 16572 31392 16584
rect 30791 16544 31392 16572
rect 30791 16541 30803 16544
rect 30745 16535 30803 16541
rect 31386 16532 31392 16544
rect 31444 16532 31450 16584
rect 29656 16476 30052 16504
rect 29365 16467 29423 16473
rect 21140 16408 21404 16436
rect 26237 16439 26295 16445
rect 21140 16396 21146 16408
rect 26237 16405 26249 16439
rect 26283 16436 26295 16439
rect 26344 16436 26372 16464
rect 26283 16408 26372 16436
rect 26283 16405 26295 16408
rect 26237 16399 26295 16405
rect 26786 16396 26792 16448
rect 26844 16396 26850 16448
rect 28442 16396 28448 16448
rect 28500 16396 28506 16448
rect 28905 16439 28963 16445
rect 28905 16405 28917 16439
rect 28951 16436 28963 16439
rect 29178 16436 29184 16448
rect 28951 16408 29184 16436
rect 28951 16405 28963 16408
rect 28905 16399 28963 16405
rect 29178 16396 29184 16408
rect 29236 16396 29242 16448
rect 29380 16436 29408 16467
rect 30024 16448 30052 16476
rect 31012 16507 31070 16513
rect 31012 16473 31024 16507
rect 31058 16504 31070 16507
rect 31478 16504 31484 16516
rect 31058 16476 31484 16504
rect 31058 16473 31070 16476
rect 31012 16467 31070 16473
rect 31478 16464 31484 16476
rect 31536 16464 31542 16516
rect 29914 16436 29920 16448
rect 29380 16408 29920 16436
rect 29914 16396 29920 16408
rect 29972 16396 29978 16448
rect 30006 16396 30012 16448
rect 30064 16396 30070 16448
rect 32125 16439 32183 16445
rect 32125 16405 32137 16439
rect 32171 16436 32183 16439
rect 32214 16436 32220 16448
rect 32171 16408 32220 16436
rect 32171 16405 32183 16408
rect 32125 16399 32183 16405
rect 32214 16396 32220 16408
rect 32272 16396 32278 16448
rect 1104 16346 35027 16368
rect 1104 16294 9390 16346
rect 9442 16294 9454 16346
rect 9506 16294 9518 16346
rect 9570 16294 9582 16346
rect 9634 16294 9646 16346
rect 9698 16294 17831 16346
rect 17883 16294 17895 16346
rect 17947 16294 17959 16346
rect 18011 16294 18023 16346
rect 18075 16294 18087 16346
rect 18139 16294 26272 16346
rect 26324 16294 26336 16346
rect 26388 16294 26400 16346
rect 26452 16294 26464 16346
rect 26516 16294 26528 16346
rect 26580 16294 34713 16346
rect 34765 16294 34777 16346
rect 34829 16294 34841 16346
rect 34893 16294 34905 16346
rect 34957 16294 34969 16346
rect 35021 16294 35027 16346
rect 1104 16272 35027 16294
rect 17678 16192 17684 16244
rect 17736 16192 17742 16244
rect 18966 16192 18972 16244
rect 19024 16192 19030 16244
rect 19426 16192 19432 16244
rect 19484 16232 19490 16244
rect 20349 16235 20407 16241
rect 20349 16232 20361 16235
rect 19484 16204 20361 16232
rect 19484 16192 19490 16204
rect 20349 16201 20361 16204
rect 20395 16201 20407 16235
rect 20349 16195 20407 16201
rect 25222 16192 25228 16244
rect 25280 16192 25286 16244
rect 25869 16235 25927 16241
rect 25869 16201 25881 16235
rect 25915 16232 25927 16235
rect 25915 16204 26096 16232
rect 25915 16201 25927 16204
rect 25869 16195 25927 16201
rect 17696 16164 17724 16192
rect 17865 16167 17923 16173
rect 17865 16164 17877 16167
rect 17696 16136 17877 16164
rect 17865 16133 17877 16136
rect 17911 16133 17923 16167
rect 17865 16127 17923 16133
rect 18049 16099 18107 16105
rect 18049 16065 18061 16099
rect 18095 16096 18107 16099
rect 18230 16096 18236 16108
rect 18095 16068 18236 16096
rect 18095 16065 18107 16068
rect 18049 16059 18107 16065
rect 18230 16056 18236 16068
rect 18288 16056 18294 16108
rect 18325 16099 18383 16105
rect 18325 16065 18337 16099
rect 18371 16096 18383 16099
rect 18984 16096 19012 16192
rect 19052 16167 19110 16173
rect 19052 16133 19064 16167
rect 19098 16164 19110 16167
rect 19886 16164 19892 16176
rect 19098 16136 19892 16164
rect 19098 16133 19110 16136
rect 19052 16127 19110 16133
rect 19886 16124 19892 16136
rect 19944 16124 19950 16176
rect 25240 16164 25268 16192
rect 25148 16136 25268 16164
rect 25148 16105 25176 16136
rect 18371 16068 19012 16096
rect 20441 16099 20499 16105
rect 18371 16065 18383 16068
rect 18325 16059 18383 16065
rect 20441 16065 20453 16099
rect 20487 16065 20499 16099
rect 20441 16059 20499 16065
rect 24673 16099 24731 16105
rect 24673 16065 24685 16099
rect 24719 16096 24731 16099
rect 25133 16099 25191 16105
rect 25133 16096 25145 16099
rect 24719 16068 25145 16096
rect 24719 16065 24731 16068
rect 24673 16059 24731 16065
rect 18506 15988 18512 16040
rect 18564 16028 18570 16040
rect 18785 16031 18843 16037
rect 18785 16028 18797 16031
rect 18564 16000 18797 16028
rect 18564 15988 18570 16000
rect 18785 15997 18797 16000
rect 18831 15997 18843 16031
rect 20456 16028 20484 16059
rect 20622 16028 20628 16040
rect 20456 16000 20628 16028
rect 18785 15991 18843 15997
rect 20622 15988 20628 16000
rect 20680 15988 20686 16040
rect 18233 15963 18291 15969
rect 18233 15929 18245 15963
rect 18279 15960 18291 15963
rect 18414 15960 18420 15972
rect 18279 15932 18420 15960
rect 18279 15929 18291 15932
rect 18233 15923 18291 15929
rect 18414 15920 18420 15932
rect 18472 15920 18478 15972
rect 20162 15920 20168 15972
rect 20220 15920 20226 15972
rect 24780 15960 24808 16068
rect 25133 16065 25145 16068
rect 25179 16065 25191 16099
rect 25774 16096 25780 16108
rect 25133 16059 25191 16065
rect 25240 16068 25780 16096
rect 24857 16031 24915 16037
rect 24857 15997 24869 16031
rect 24903 16028 24915 16031
rect 25240 16028 25268 16068
rect 25774 16056 25780 16068
rect 25832 16056 25838 16108
rect 25958 16056 25964 16108
rect 26016 16056 26022 16108
rect 26068 16040 26096 16204
rect 26142 16192 26148 16244
rect 26200 16192 26206 16244
rect 26602 16192 26608 16244
rect 26660 16192 26666 16244
rect 26786 16192 26792 16244
rect 26844 16192 26850 16244
rect 26970 16192 26976 16244
rect 27028 16192 27034 16244
rect 28442 16192 28448 16244
rect 28500 16192 28506 16244
rect 29086 16192 29092 16244
rect 29144 16232 29150 16244
rect 29825 16235 29883 16241
rect 29825 16232 29837 16235
rect 29144 16204 29837 16232
rect 29144 16192 29150 16204
rect 29825 16201 29837 16204
rect 29871 16201 29883 16235
rect 29825 16195 29883 16201
rect 29914 16192 29920 16244
rect 29972 16232 29978 16244
rect 31297 16235 31355 16241
rect 31297 16232 31309 16235
rect 29972 16204 31309 16232
rect 29972 16192 29978 16204
rect 31297 16201 31309 16204
rect 31343 16201 31355 16235
rect 31297 16195 31355 16201
rect 26620 16164 26648 16192
rect 26804 16164 26832 16192
rect 28086 16167 28144 16173
rect 28086 16164 28098 16167
rect 26620 16136 26740 16164
rect 26804 16136 28098 16164
rect 26605 16099 26663 16105
rect 26605 16065 26617 16099
rect 26651 16065 26663 16099
rect 26712 16096 26740 16136
rect 28086 16133 28098 16136
rect 28132 16133 28144 16167
rect 28460 16164 28488 16192
rect 28690 16167 28748 16173
rect 28690 16164 28702 16167
rect 28460 16136 28702 16164
rect 28086 16127 28144 16133
rect 28690 16133 28702 16136
rect 28736 16133 28748 16167
rect 28690 16127 28748 16133
rect 30374 16124 30380 16176
rect 30432 16124 30438 16176
rect 31312 16164 31340 16195
rect 31312 16136 31708 16164
rect 26789 16099 26847 16105
rect 26789 16096 26801 16099
rect 26712 16068 26801 16096
rect 26605 16059 26663 16065
rect 26789 16065 26801 16068
rect 26835 16065 26847 16099
rect 26789 16059 26847 16065
rect 24903 16000 25268 16028
rect 25317 16031 25375 16037
rect 24903 15997 24915 16000
rect 24857 15991 24915 15997
rect 25317 15997 25329 16031
rect 25363 16028 25375 16031
rect 25363 16000 25636 16028
rect 25363 15997 25375 16000
rect 25317 15991 25375 15997
rect 25608 15969 25636 16000
rect 26050 15988 26056 16040
rect 26108 16028 26114 16040
rect 26421 16031 26479 16037
rect 26421 16028 26433 16031
rect 26108 16000 26433 16028
rect 26108 15988 26114 16000
rect 26421 15997 26433 16000
rect 26467 15997 26479 16031
rect 26421 15991 26479 15997
rect 25593 15963 25651 15969
rect 24780 15932 25544 15960
rect 24486 15852 24492 15904
rect 24544 15852 24550 15904
rect 24578 15852 24584 15904
rect 24636 15892 24642 15904
rect 24949 15895 25007 15901
rect 24949 15892 24961 15895
rect 24636 15864 24961 15892
rect 24636 15852 24642 15864
rect 24949 15861 24961 15864
rect 24995 15861 25007 15895
rect 25516 15892 25544 15932
rect 25593 15929 25605 15963
rect 25639 15960 25651 15963
rect 26234 15960 26240 15972
rect 25639 15932 26240 15960
rect 25639 15929 25651 15932
rect 25593 15923 25651 15929
rect 26234 15920 26240 15932
rect 26292 15920 26298 15972
rect 25866 15892 25872 15904
rect 25516 15864 25872 15892
rect 24949 15855 25007 15861
rect 25866 15852 25872 15864
rect 25924 15892 25930 15904
rect 26620 15892 26648 16059
rect 27614 16056 27620 16108
rect 27672 16096 27678 16108
rect 28353 16099 28411 16105
rect 28353 16096 28365 16099
rect 27672 16068 28365 16096
rect 27672 16056 27678 16068
rect 28353 16065 28365 16068
rect 28399 16096 28411 16099
rect 28445 16099 28503 16105
rect 28445 16096 28457 16099
rect 28399 16068 28457 16096
rect 28399 16065 28411 16068
rect 28353 16059 28411 16065
rect 28445 16065 28457 16068
rect 28491 16096 28503 16099
rect 28534 16096 28540 16108
rect 28491 16068 28540 16096
rect 28491 16065 28503 16068
rect 28445 16059 28503 16065
rect 28534 16056 28540 16068
rect 28592 16056 28598 16108
rect 29730 16056 29736 16108
rect 29788 16096 29794 16108
rect 30173 16099 30231 16105
rect 30173 16096 30185 16099
rect 29788 16068 30185 16096
rect 29788 16056 29794 16068
rect 30173 16065 30185 16068
rect 30219 16065 30231 16099
rect 30392 16096 30420 16124
rect 31680 16105 31708 16136
rect 31573 16099 31631 16105
rect 31573 16096 31585 16099
rect 30392 16068 31585 16096
rect 30173 16059 30231 16065
rect 31573 16065 31585 16068
rect 31619 16065 31631 16099
rect 31573 16059 31631 16065
rect 31665 16099 31723 16105
rect 31665 16065 31677 16099
rect 31711 16065 31723 16099
rect 31665 16059 31723 16065
rect 29917 16031 29975 16037
rect 29917 15997 29929 16031
rect 29963 15997 29975 16031
rect 29917 15991 29975 15997
rect 25924 15864 26648 15892
rect 29932 15892 29960 15991
rect 30650 15892 30656 15904
rect 29932 15864 30656 15892
rect 25924 15852 25930 15864
rect 30650 15852 30656 15864
rect 30708 15852 30714 15904
rect 31386 15852 31392 15904
rect 31444 15852 31450 15904
rect 1104 15802 34868 15824
rect 1104 15750 5170 15802
rect 5222 15750 5234 15802
rect 5286 15750 5298 15802
rect 5350 15750 5362 15802
rect 5414 15750 5426 15802
rect 5478 15750 13611 15802
rect 13663 15750 13675 15802
rect 13727 15750 13739 15802
rect 13791 15750 13803 15802
rect 13855 15750 13867 15802
rect 13919 15750 22052 15802
rect 22104 15750 22116 15802
rect 22168 15750 22180 15802
rect 22232 15750 22244 15802
rect 22296 15750 22308 15802
rect 22360 15750 30493 15802
rect 30545 15750 30557 15802
rect 30609 15750 30621 15802
rect 30673 15750 30685 15802
rect 30737 15750 30749 15802
rect 30801 15750 34868 15802
rect 1104 15728 34868 15750
rect 24578 15688 24584 15700
rect 24044 15660 24584 15688
rect 24044 15493 24072 15660
rect 24578 15648 24584 15660
rect 24636 15648 24642 15700
rect 25869 15691 25927 15697
rect 25869 15657 25881 15691
rect 25915 15688 25927 15691
rect 26050 15688 26056 15700
rect 25915 15660 26056 15688
rect 25915 15657 25927 15660
rect 25869 15651 25927 15657
rect 26050 15648 26056 15660
rect 26108 15648 26114 15700
rect 28258 15648 28264 15700
rect 28316 15688 28322 15700
rect 28353 15691 28411 15697
rect 28353 15688 28365 15691
rect 28316 15660 28365 15688
rect 28316 15648 28322 15660
rect 28353 15657 28365 15660
rect 28399 15657 28411 15691
rect 28353 15651 28411 15657
rect 29730 15648 29736 15700
rect 29788 15648 29794 15700
rect 30006 15648 30012 15700
rect 30064 15648 30070 15700
rect 30374 15648 30380 15700
rect 30432 15648 30438 15700
rect 31478 15648 31484 15700
rect 31536 15648 31542 15700
rect 28902 15620 28908 15632
rect 28552 15592 28908 15620
rect 24029 15487 24087 15493
rect 24029 15453 24041 15487
rect 24075 15453 24087 15487
rect 24029 15447 24087 15453
rect 24394 15444 24400 15496
rect 24452 15484 24458 15496
rect 27249 15487 27307 15493
rect 27249 15484 27261 15487
rect 24452 15456 24900 15484
rect 24452 15444 24458 15456
rect 24872 15428 24900 15456
rect 25608 15456 27261 15484
rect 24302 15376 24308 15428
rect 24360 15376 24366 15428
rect 24670 15425 24676 15428
rect 24664 15379 24676 15425
rect 24670 15376 24676 15379
rect 24728 15376 24734 15428
rect 24854 15376 24860 15428
rect 24912 15376 24918 15428
rect 24210 15308 24216 15360
rect 24268 15308 24274 15360
rect 24320 15348 24348 15376
rect 25608 15348 25636 15456
rect 27249 15453 27261 15456
rect 27295 15484 27307 15487
rect 27614 15484 27620 15496
rect 27295 15456 27620 15484
rect 27295 15453 27307 15456
rect 27249 15447 27307 15453
rect 27614 15444 27620 15456
rect 27672 15444 27678 15496
rect 28166 15444 28172 15496
rect 28224 15444 28230 15496
rect 28552 15493 28580 15592
rect 28902 15580 28908 15592
rect 28960 15620 28966 15632
rect 30392 15620 30420 15648
rect 28960 15592 30420 15620
rect 28960 15580 28966 15592
rect 28813 15555 28871 15561
rect 28813 15521 28825 15555
rect 28859 15552 28871 15555
rect 29086 15552 29092 15564
rect 28859 15524 29092 15552
rect 28859 15521 28871 15524
rect 28813 15515 28871 15521
rect 29086 15512 29092 15524
rect 29144 15512 29150 15564
rect 28537 15487 28595 15493
rect 28537 15453 28549 15487
rect 28583 15453 28595 15487
rect 28537 15447 28595 15453
rect 28721 15487 28779 15493
rect 28721 15453 28733 15487
rect 28767 15453 28779 15487
rect 28721 15447 28779 15453
rect 26234 15416 26240 15428
rect 25792 15388 26240 15416
rect 25792 15357 25820 15388
rect 26160 15360 26188 15388
rect 26234 15376 26240 15388
rect 26292 15376 26298 15428
rect 26694 15376 26700 15428
rect 26752 15416 26758 15428
rect 26982 15419 27040 15425
rect 26982 15416 26994 15419
rect 26752 15388 26994 15416
rect 26752 15376 26758 15388
rect 26982 15385 26994 15388
rect 27028 15385 27040 15419
rect 28736 15416 28764 15447
rect 28902 15444 28908 15496
rect 28960 15484 28966 15496
rect 28997 15487 29055 15493
rect 28997 15484 29009 15487
rect 28960 15456 29009 15484
rect 28960 15444 28966 15456
rect 28997 15453 29009 15456
rect 29043 15453 29055 15487
rect 28997 15447 29055 15453
rect 29181 15487 29239 15493
rect 29181 15453 29193 15487
rect 29227 15484 29239 15487
rect 29549 15487 29607 15493
rect 29549 15484 29561 15487
rect 29227 15456 29561 15484
rect 29227 15453 29239 15456
rect 29181 15447 29239 15453
rect 29549 15453 29561 15456
rect 29595 15453 29607 15487
rect 29549 15447 29607 15453
rect 31294 15444 31300 15496
rect 31352 15484 31358 15496
rect 31389 15487 31447 15493
rect 31389 15484 31401 15487
rect 31352 15456 31401 15484
rect 31352 15444 31358 15456
rect 31389 15453 31401 15456
rect 31435 15453 31447 15487
rect 31389 15447 31447 15453
rect 31662 15444 31668 15496
rect 31720 15444 31726 15496
rect 29362 15416 29368 15428
rect 28736 15388 29368 15416
rect 26982 15379 27040 15385
rect 29362 15376 29368 15388
rect 29420 15376 29426 15428
rect 30558 15376 30564 15428
rect 30616 15416 30622 15428
rect 31122 15419 31180 15425
rect 31122 15416 31134 15419
rect 30616 15388 31134 15416
rect 30616 15376 30622 15388
rect 31122 15385 31134 15388
rect 31168 15385 31180 15419
rect 31122 15379 31180 15385
rect 24320 15320 25636 15348
rect 25777 15351 25835 15357
rect 25777 15317 25789 15351
rect 25823 15317 25835 15351
rect 25777 15311 25835 15317
rect 26142 15308 26148 15360
rect 26200 15308 26206 15360
rect 27982 15308 27988 15360
rect 28040 15308 28046 15360
rect 1104 15258 35027 15280
rect 1104 15206 9390 15258
rect 9442 15206 9454 15258
rect 9506 15206 9518 15258
rect 9570 15206 9582 15258
rect 9634 15206 9646 15258
rect 9698 15206 17831 15258
rect 17883 15206 17895 15258
rect 17947 15206 17959 15258
rect 18011 15206 18023 15258
rect 18075 15206 18087 15258
rect 18139 15206 26272 15258
rect 26324 15206 26336 15258
rect 26388 15206 26400 15258
rect 26452 15206 26464 15258
rect 26516 15206 26528 15258
rect 26580 15206 34713 15258
rect 34765 15206 34777 15258
rect 34829 15206 34841 15258
rect 34893 15206 34905 15258
rect 34957 15206 34969 15258
rect 35021 15206 35027 15258
rect 1104 15184 35027 15206
rect 20622 15104 20628 15156
rect 20680 15144 20686 15156
rect 21177 15147 21235 15153
rect 21177 15144 21189 15147
rect 20680 15116 21189 15144
rect 20680 15104 20686 15116
rect 21177 15113 21189 15116
rect 21223 15113 21235 15147
rect 21177 15107 21235 15113
rect 25869 15147 25927 15153
rect 25869 15113 25881 15147
rect 25915 15144 25927 15147
rect 26421 15147 26479 15153
rect 25915 15116 26004 15144
rect 25915 15113 25927 15116
rect 25869 15107 25927 15113
rect 25976 15088 26004 15116
rect 26421 15113 26433 15147
rect 26467 15144 26479 15147
rect 26602 15144 26608 15156
rect 26467 15116 26608 15144
rect 26467 15113 26479 15116
rect 26421 15107 26479 15113
rect 26602 15104 26608 15116
rect 26660 15104 26666 15156
rect 26694 15104 26700 15156
rect 26752 15104 26758 15156
rect 28997 15147 29055 15153
rect 28997 15113 29009 15147
rect 29043 15144 29055 15147
rect 29362 15144 29368 15156
rect 29043 15116 29368 15144
rect 29043 15113 29055 15116
rect 28997 15107 29055 15113
rect 29362 15104 29368 15116
rect 29420 15104 29426 15156
rect 30009 15147 30067 15153
rect 30009 15113 30021 15147
rect 30055 15144 30067 15147
rect 30558 15144 30564 15156
rect 30055 15116 30564 15144
rect 30055 15113 30067 15116
rect 30009 15107 30067 15113
rect 30558 15104 30564 15116
rect 30616 15104 30622 15156
rect 31386 15104 31392 15156
rect 31444 15104 31450 15156
rect 31662 15104 31668 15156
rect 31720 15104 31726 15156
rect 22646 15076 22652 15088
rect 19812 15048 22652 15076
rect 19812 15017 19840 15048
rect 22646 15036 22652 15048
rect 22704 15036 22710 15088
rect 23032 15048 23428 15076
rect 20070 15017 20076 15020
rect 19797 15011 19855 15017
rect 19797 14977 19809 15011
rect 19843 14977 19855 15011
rect 20064 15008 20076 15017
rect 20031 14980 20076 15008
rect 19797 14971 19855 14977
rect 20064 14971 20076 14980
rect 20070 14968 20076 14971
rect 20128 14968 20134 15020
rect 23032 15017 23060 15048
rect 23290 15017 23296 15020
rect 23017 15011 23075 15017
rect 23017 14977 23029 15011
rect 23063 14977 23075 15011
rect 23017 14971 23075 14977
rect 23284 14971 23296 15017
rect 23290 14968 23296 14971
rect 23348 14968 23354 15020
rect 23400 15008 23428 15048
rect 24210 15036 24216 15088
rect 24268 15076 24274 15088
rect 24734 15079 24792 15085
rect 24734 15076 24746 15079
rect 24268 15048 24746 15076
rect 24268 15036 24274 15048
rect 24734 15045 24746 15048
rect 24780 15045 24792 15079
rect 24734 15039 24792 15045
rect 25958 15036 25964 15088
rect 26016 15036 26022 15088
rect 27884 15079 27942 15085
rect 27884 15045 27896 15079
rect 27930 15076 27942 15079
rect 27982 15076 27988 15088
rect 27930 15048 27988 15076
rect 27930 15045 27942 15048
rect 27884 15039 27942 15045
rect 27982 15036 27988 15048
rect 28040 15036 28046 15088
rect 24394 15008 24400 15020
rect 23400 14980 24400 15008
rect 24394 14968 24400 14980
rect 24452 14968 24458 15020
rect 26050 14968 26056 15020
rect 26108 15008 26114 15020
rect 26145 15011 26203 15017
rect 26145 15008 26157 15011
rect 26108 14980 26157 15008
rect 26108 14968 26114 14980
rect 26145 14977 26157 14980
rect 26191 14977 26203 15011
rect 26145 14971 26203 14977
rect 26234 14968 26240 15020
rect 26292 14968 26298 15020
rect 26510 14968 26516 15020
rect 26568 14968 26574 15020
rect 27614 14968 27620 15020
rect 27672 14968 27678 15020
rect 29825 15011 29883 15017
rect 29825 14977 29837 15011
rect 29871 15008 29883 15011
rect 31404 15008 31432 15104
rect 29871 14980 31432 15008
rect 29871 14977 29883 14980
rect 29825 14971 29883 14977
rect 31478 14968 31484 15020
rect 31536 14968 31542 15020
rect 24302 14900 24308 14952
rect 24360 14940 24366 14952
rect 24489 14943 24547 14949
rect 24489 14940 24501 14943
rect 24360 14912 24501 14940
rect 24360 14900 24366 14912
rect 24489 14909 24501 14912
rect 24535 14909 24547 14943
rect 31297 14943 31355 14949
rect 31297 14940 31309 14943
rect 24489 14903 24547 14909
rect 28644 14912 31309 14940
rect 24397 14807 24455 14813
rect 24397 14773 24409 14807
rect 24443 14804 24455 14807
rect 25774 14804 25780 14816
rect 24443 14776 25780 14804
rect 24443 14773 24455 14776
rect 24397 14767 24455 14773
rect 25774 14764 25780 14776
rect 25832 14804 25838 14816
rect 25961 14807 26019 14813
rect 25961 14804 25973 14807
rect 25832 14776 25973 14804
rect 25832 14764 25838 14776
rect 25961 14773 25973 14776
rect 26007 14773 26019 14807
rect 25961 14767 26019 14773
rect 27890 14764 27896 14816
rect 27948 14804 27954 14816
rect 28644 14804 28672 14912
rect 31297 14909 31309 14912
rect 31343 14909 31355 14943
rect 31297 14903 31355 14909
rect 27948 14776 28672 14804
rect 27948 14764 27954 14776
rect 1104 14714 34868 14736
rect 1104 14662 5170 14714
rect 5222 14662 5234 14714
rect 5286 14662 5298 14714
rect 5350 14662 5362 14714
rect 5414 14662 5426 14714
rect 5478 14662 13611 14714
rect 13663 14662 13675 14714
rect 13727 14662 13739 14714
rect 13791 14662 13803 14714
rect 13855 14662 13867 14714
rect 13919 14662 22052 14714
rect 22104 14662 22116 14714
rect 22168 14662 22180 14714
rect 22232 14662 22244 14714
rect 22296 14662 22308 14714
rect 22360 14662 30493 14714
rect 30545 14662 30557 14714
rect 30609 14662 30621 14714
rect 30673 14662 30685 14714
rect 30737 14662 30749 14714
rect 30801 14662 34868 14714
rect 1104 14640 34868 14662
rect 23290 14560 23296 14612
rect 23348 14600 23354 14612
rect 23385 14603 23443 14609
rect 23385 14600 23397 14603
rect 23348 14572 23397 14600
rect 23348 14560 23354 14572
rect 23385 14569 23397 14572
rect 23431 14569 23443 14603
rect 23385 14563 23443 14569
rect 24581 14603 24639 14609
rect 24581 14569 24593 14603
rect 24627 14600 24639 14603
rect 24670 14600 24676 14612
rect 24627 14572 24676 14600
rect 24627 14569 24639 14572
rect 24581 14563 24639 14569
rect 24670 14560 24676 14572
rect 24728 14560 24734 14612
rect 25958 14560 25964 14612
rect 26016 14560 26022 14612
rect 26145 14603 26203 14609
rect 26145 14569 26157 14603
rect 26191 14600 26203 14603
rect 26510 14600 26516 14612
rect 26191 14572 26516 14600
rect 26191 14569 26203 14572
rect 26145 14563 26203 14569
rect 26510 14560 26516 14572
rect 26568 14560 26574 14612
rect 28166 14560 28172 14612
rect 28224 14600 28230 14612
rect 28261 14603 28319 14609
rect 28261 14600 28273 14603
rect 28224 14572 28273 14600
rect 28224 14560 28230 14572
rect 28261 14569 28273 14572
rect 28307 14569 28319 14603
rect 28261 14563 28319 14569
rect 22465 14467 22523 14473
rect 22465 14433 22477 14467
rect 22511 14464 22523 14467
rect 25406 14464 25412 14476
rect 22511 14436 25412 14464
rect 22511 14433 22523 14436
rect 22465 14427 22523 14433
rect 25406 14424 25412 14436
rect 25464 14424 25470 14476
rect 25777 14467 25835 14473
rect 25777 14433 25789 14467
rect 25823 14464 25835 14467
rect 25976 14464 26004 14560
rect 25823 14436 26004 14464
rect 25823 14433 25835 14436
rect 25777 14427 25835 14433
rect 22649 14399 22707 14405
rect 22649 14365 22661 14399
rect 22695 14365 22707 14399
rect 22649 14359 22707 14365
rect 22833 14399 22891 14405
rect 22833 14365 22845 14399
rect 22879 14396 22891 14399
rect 23201 14399 23259 14405
rect 23201 14396 23213 14399
rect 22879 14368 23213 14396
rect 22879 14365 22891 14368
rect 22833 14359 22891 14365
rect 23201 14365 23213 14368
rect 23247 14365 23259 14399
rect 23201 14359 23259 14365
rect 24397 14399 24455 14405
rect 24397 14365 24409 14399
rect 24443 14396 24455 14399
rect 24486 14396 24492 14408
rect 24443 14368 24492 14396
rect 24443 14365 24455 14368
rect 24397 14359 24455 14365
rect 1670 14288 1676 14340
rect 1728 14328 1734 14340
rect 22664 14328 22692 14359
rect 24486 14356 24492 14368
rect 24544 14356 24550 14408
rect 1728 14300 22692 14328
rect 25424 14328 25452 14424
rect 25866 14356 25872 14408
rect 25924 14396 25930 14408
rect 25961 14399 26019 14405
rect 25961 14396 25973 14399
rect 25924 14368 25973 14396
rect 25924 14356 25930 14368
rect 25961 14365 25973 14368
rect 26007 14365 26019 14399
rect 25961 14359 26019 14365
rect 27890 14356 27896 14408
rect 27948 14356 27954 14408
rect 28077 14399 28135 14405
rect 28077 14365 28089 14399
rect 28123 14396 28135 14399
rect 28442 14396 28448 14408
rect 28123 14368 28448 14396
rect 28123 14365 28135 14368
rect 28077 14359 28135 14365
rect 28442 14356 28448 14368
rect 28500 14356 28506 14408
rect 27908 14328 27936 14356
rect 25424 14300 27936 14328
rect 1728 14288 1734 14300
rect 1104 14170 35027 14192
rect 1104 14118 9390 14170
rect 9442 14118 9454 14170
rect 9506 14118 9518 14170
rect 9570 14118 9582 14170
rect 9634 14118 9646 14170
rect 9698 14118 17831 14170
rect 17883 14118 17895 14170
rect 17947 14118 17959 14170
rect 18011 14118 18023 14170
rect 18075 14118 18087 14170
rect 18139 14118 26272 14170
rect 26324 14118 26336 14170
rect 26388 14118 26400 14170
rect 26452 14118 26464 14170
rect 26516 14118 26528 14170
rect 26580 14118 34713 14170
rect 34765 14118 34777 14170
rect 34829 14118 34841 14170
rect 34893 14118 34905 14170
rect 34957 14118 34969 14170
rect 35021 14118 35027 14170
rect 1104 14096 35027 14118
rect 1104 13626 34868 13648
rect 1104 13574 5170 13626
rect 5222 13574 5234 13626
rect 5286 13574 5298 13626
rect 5350 13574 5362 13626
rect 5414 13574 5426 13626
rect 5478 13574 13611 13626
rect 13663 13574 13675 13626
rect 13727 13574 13739 13626
rect 13791 13574 13803 13626
rect 13855 13574 13867 13626
rect 13919 13574 22052 13626
rect 22104 13574 22116 13626
rect 22168 13574 22180 13626
rect 22232 13574 22244 13626
rect 22296 13574 22308 13626
rect 22360 13574 30493 13626
rect 30545 13574 30557 13626
rect 30609 13574 30621 13626
rect 30673 13574 30685 13626
rect 30737 13574 30749 13626
rect 30801 13574 34868 13626
rect 1104 13552 34868 13574
rect 1104 13082 35027 13104
rect 1104 13030 9390 13082
rect 9442 13030 9454 13082
rect 9506 13030 9518 13082
rect 9570 13030 9582 13082
rect 9634 13030 9646 13082
rect 9698 13030 17831 13082
rect 17883 13030 17895 13082
rect 17947 13030 17959 13082
rect 18011 13030 18023 13082
rect 18075 13030 18087 13082
rect 18139 13030 26272 13082
rect 26324 13030 26336 13082
rect 26388 13030 26400 13082
rect 26452 13030 26464 13082
rect 26516 13030 26528 13082
rect 26580 13030 34713 13082
rect 34765 13030 34777 13082
rect 34829 13030 34841 13082
rect 34893 13030 34905 13082
rect 34957 13030 34969 13082
rect 35021 13030 35027 13082
rect 1104 13008 35027 13030
rect 1104 12538 34868 12560
rect 1104 12486 5170 12538
rect 5222 12486 5234 12538
rect 5286 12486 5298 12538
rect 5350 12486 5362 12538
rect 5414 12486 5426 12538
rect 5478 12486 13611 12538
rect 13663 12486 13675 12538
rect 13727 12486 13739 12538
rect 13791 12486 13803 12538
rect 13855 12486 13867 12538
rect 13919 12486 22052 12538
rect 22104 12486 22116 12538
rect 22168 12486 22180 12538
rect 22232 12486 22244 12538
rect 22296 12486 22308 12538
rect 22360 12486 30493 12538
rect 30545 12486 30557 12538
rect 30609 12486 30621 12538
rect 30673 12486 30685 12538
rect 30737 12486 30749 12538
rect 30801 12486 34868 12538
rect 1104 12464 34868 12486
rect 16022 12180 16028 12232
rect 16080 12220 16086 12232
rect 33965 12223 34023 12229
rect 33965 12220 33977 12223
rect 16080 12192 33977 12220
rect 16080 12180 16086 12192
rect 33965 12189 33977 12192
rect 34011 12189 34023 12223
rect 33965 12183 34023 12189
rect 34146 12044 34152 12096
rect 34204 12044 34210 12096
rect 1104 11994 35027 12016
rect 1104 11942 9390 11994
rect 9442 11942 9454 11994
rect 9506 11942 9518 11994
rect 9570 11942 9582 11994
rect 9634 11942 9646 11994
rect 9698 11942 17831 11994
rect 17883 11942 17895 11994
rect 17947 11942 17959 11994
rect 18011 11942 18023 11994
rect 18075 11942 18087 11994
rect 18139 11942 26272 11994
rect 26324 11942 26336 11994
rect 26388 11942 26400 11994
rect 26452 11942 26464 11994
rect 26516 11942 26528 11994
rect 26580 11942 34713 11994
rect 34765 11942 34777 11994
rect 34829 11942 34841 11994
rect 34893 11942 34905 11994
rect 34957 11942 34969 11994
rect 35021 11942 35027 11994
rect 1104 11920 35027 11942
rect 34146 11840 34152 11892
rect 34204 11840 34210 11892
rect 34164 11753 34192 11840
rect 34149 11747 34207 11753
rect 34149 11713 34161 11747
rect 34195 11713 34207 11747
rect 34149 11707 34207 11713
rect 34425 11611 34483 11617
rect 34425 11577 34437 11611
rect 34471 11608 34483 11611
rect 34514 11608 34520 11620
rect 34471 11580 34520 11608
rect 34471 11577 34483 11580
rect 34425 11571 34483 11577
rect 34514 11568 34520 11580
rect 34572 11568 34578 11620
rect 1104 11450 34868 11472
rect 1104 11398 5170 11450
rect 5222 11398 5234 11450
rect 5286 11398 5298 11450
rect 5350 11398 5362 11450
rect 5414 11398 5426 11450
rect 5478 11398 13611 11450
rect 13663 11398 13675 11450
rect 13727 11398 13739 11450
rect 13791 11398 13803 11450
rect 13855 11398 13867 11450
rect 13919 11398 22052 11450
rect 22104 11398 22116 11450
rect 22168 11398 22180 11450
rect 22232 11398 22244 11450
rect 22296 11398 22308 11450
rect 22360 11398 30493 11450
rect 30545 11398 30557 11450
rect 30609 11398 30621 11450
rect 30673 11398 30685 11450
rect 30737 11398 30749 11450
rect 30801 11398 34868 11450
rect 1104 11376 34868 11398
rect 1104 10906 35027 10928
rect 1104 10854 9390 10906
rect 9442 10854 9454 10906
rect 9506 10854 9518 10906
rect 9570 10854 9582 10906
rect 9634 10854 9646 10906
rect 9698 10854 17831 10906
rect 17883 10854 17895 10906
rect 17947 10854 17959 10906
rect 18011 10854 18023 10906
rect 18075 10854 18087 10906
rect 18139 10854 26272 10906
rect 26324 10854 26336 10906
rect 26388 10854 26400 10906
rect 26452 10854 26464 10906
rect 26516 10854 26528 10906
rect 26580 10854 34713 10906
rect 34765 10854 34777 10906
rect 34829 10854 34841 10906
rect 34893 10854 34905 10906
rect 34957 10854 34969 10906
rect 35021 10854 35027 10906
rect 1104 10832 35027 10854
rect 1104 10362 34868 10384
rect 1104 10310 5170 10362
rect 5222 10310 5234 10362
rect 5286 10310 5298 10362
rect 5350 10310 5362 10362
rect 5414 10310 5426 10362
rect 5478 10310 13611 10362
rect 13663 10310 13675 10362
rect 13727 10310 13739 10362
rect 13791 10310 13803 10362
rect 13855 10310 13867 10362
rect 13919 10310 22052 10362
rect 22104 10310 22116 10362
rect 22168 10310 22180 10362
rect 22232 10310 22244 10362
rect 22296 10310 22308 10362
rect 22360 10310 30493 10362
rect 30545 10310 30557 10362
rect 30609 10310 30621 10362
rect 30673 10310 30685 10362
rect 30737 10310 30749 10362
rect 30801 10310 34868 10362
rect 1104 10288 34868 10310
rect 1394 10004 1400 10056
rect 1452 10004 1458 10056
rect 1104 9818 35027 9840
rect 1104 9766 9390 9818
rect 9442 9766 9454 9818
rect 9506 9766 9518 9818
rect 9570 9766 9582 9818
rect 9634 9766 9646 9818
rect 9698 9766 17831 9818
rect 17883 9766 17895 9818
rect 17947 9766 17959 9818
rect 18011 9766 18023 9818
rect 18075 9766 18087 9818
rect 18139 9766 26272 9818
rect 26324 9766 26336 9818
rect 26388 9766 26400 9818
rect 26452 9766 26464 9818
rect 26516 9766 26528 9818
rect 26580 9766 34713 9818
rect 34765 9766 34777 9818
rect 34829 9766 34841 9818
rect 34893 9766 34905 9818
rect 34957 9766 34969 9818
rect 35021 9766 35027 9818
rect 1104 9744 35027 9766
rect 1104 9274 34868 9296
rect 1104 9222 5170 9274
rect 5222 9222 5234 9274
rect 5286 9222 5298 9274
rect 5350 9222 5362 9274
rect 5414 9222 5426 9274
rect 5478 9222 13611 9274
rect 13663 9222 13675 9274
rect 13727 9222 13739 9274
rect 13791 9222 13803 9274
rect 13855 9222 13867 9274
rect 13919 9222 22052 9274
rect 22104 9222 22116 9274
rect 22168 9222 22180 9274
rect 22232 9222 22244 9274
rect 22296 9222 22308 9274
rect 22360 9222 30493 9274
rect 30545 9222 30557 9274
rect 30609 9222 30621 9274
rect 30673 9222 30685 9274
rect 30737 9222 30749 9274
rect 30801 9222 34868 9274
rect 1104 9200 34868 9222
rect 1104 8730 35027 8752
rect 1104 8678 9390 8730
rect 9442 8678 9454 8730
rect 9506 8678 9518 8730
rect 9570 8678 9582 8730
rect 9634 8678 9646 8730
rect 9698 8678 17831 8730
rect 17883 8678 17895 8730
rect 17947 8678 17959 8730
rect 18011 8678 18023 8730
rect 18075 8678 18087 8730
rect 18139 8678 26272 8730
rect 26324 8678 26336 8730
rect 26388 8678 26400 8730
rect 26452 8678 26464 8730
rect 26516 8678 26528 8730
rect 26580 8678 34713 8730
rect 34765 8678 34777 8730
rect 34829 8678 34841 8730
rect 34893 8678 34905 8730
rect 34957 8678 34969 8730
rect 35021 8678 35027 8730
rect 1104 8656 35027 8678
rect 1104 8186 34868 8208
rect 1104 8134 5170 8186
rect 5222 8134 5234 8186
rect 5286 8134 5298 8186
rect 5350 8134 5362 8186
rect 5414 8134 5426 8186
rect 5478 8134 13611 8186
rect 13663 8134 13675 8186
rect 13727 8134 13739 8186
rect 13791 8134 13803 8186
rect 13855 8134 13867 8186
rect 13919 8134 22052 8186
rect 22104 8134 22116 8186
rect 22168 8134 22180 8186
rect 22232 8134 22244 8186
rect 22296 8134 22308 8186
rect 22360 8134 30493 8186
rect 30545 8134 30557 8186
rect 30609 8134 30621 8186
rect 30673 8134 30685 8186
rect 30737 8134 30749 8186
rect 30801 8134 34868 8186
rect 1104 8112 34868 8134
rect 1104 7642 35027 7664
rect 1104 7590 9390 7642
rect 9442 7590 9454 7642
rect 9506 7590 9518 7642
rect 9570 7590 9582 7642
rect 9634 7590 9646 7642
rect 9698 7590 17831 7642
rect 17883 7590 17895 7642
rect 17947 7590 17959 7642
rect 18011 7590 18023 7642
rect 18075 7590 18087 7642
rect 18139 7590 26272 7642
rect 26324 7590 26336 7642
rect 26388 7590 26400 7642
rect 26452 7590 26464 7642
rect 26516 7590 26528 7642
rect 26580 7590 34713 7642
rect 34765 7590 34777 7642
rect 34829 7590 34841 7642
rect 34893 7590 34905 7642
rect 34957 7590 34969 7642
rect 35021 7590 35027 7642
rect 1104 7568 35027 7590
rect 1104 7098 34868 7120
rect 1104 7046 5170 7098
rect 5222 7046 5234 7098
rect 5286 7046 5298 7098
rect 5350 7046 5362 7098
rect 5414 7046 5426 7098
rect 5478 7046 13611 7098
rect 13663 7046 13675 7098
rect 13727 7046 13739 7098
rect 13791 7046 13803 7098
rect 13855 7046 13867 7098
rect 13919 7046 22052 7098
rect 22104 7046 22116 7098
rect 22168 7046 22180 7098
rect 22232 7046 22244 7098
rect 22296 7046 22308 7098
rect 22360 7046 30493 7098
rect 30545 7046 30557 7098
rect 30609 7046 30621 7098
rect 30673 7046 30685 7098
rect 30737 7046 30749 7098
rect 30801 7046 34868 7098
rect 1104 7024 34868 7046
rect 1104 6554 35027 6576
rect 1104 6502 9390 6554
rect 9442 6502 9454 6554
rect 9506 6502 9518 6554
rect 9570 6502 9582 6554
rect 9634 6502 9646 6554
rect 9698 6502 17831 6554
rect 17883 6502 17895 6554
rect 17947 6502 17959 6554
rect 18011 6502 18023 6554
rect 18075 6502 18087 6554
rect 18139 6502 26272 6554
rect 26324 6502 26336 6554
rect 26388 6502 26400 6554
rect 26452 6502 26464 6554
rect 26516 6502 26528 6554
rect 26580 6502 34713 6554
rect 34765 6502 34777 6554
rect 34829 6502 34841 6554
rect 34893 6502 34905 6554
rect 34957 6502 34969 6554
rect 35021 6502 35027 6554
rect 1104 6480 35027 6502
rect 1104 6010 34868 6032
rect 1104 5958 5170 6010
rect 5222 5958 5234 6010
rect 5286 5958 5298 6010
rect 5350 5958 5362 6010
rect 5414 5958 5426 6010
rect 5478 5958 13611 6010
rect 13663 5958 13675 6010
rect 13727 5958 13739 6010
rect 13791 5958 13803 6010
rect 13855 5958 13867 6010
rect 13919 5958 22052 6010
rect 22104 5958 22116 6010
rect 22168 5958 22180 6010
rect 22232 5958 22244 6010
rect 22296 5958 22308 6010
rect 22360 5958 30493 6010
rect 30545 5958 30557 6010
rect 30609 5958 30621 6010
rect 30673 5958 30685 6010
rect 30737 5958 30749 6010
rect 30801 5958 34868 6010
rect 1104 5936 34868 5958
rect 1104 5466 35027 5488
rect 1104 5414 9390 5466
rect 9442 5414 9454 5466
rect 9506 5414 9518 5466
rect 9570 5414 9582 5466
rect 9634 5414 9646 5466
rect 9698 5414 17831 5466
rect 17883 5414 17895 5466
rect 17947 5414 17959 5466
rect 18011 5414 18023 5466
rect 18075 5414 18087 5466
rect 18139 5414 26272 5466
rect 26324 5414 26336 5466
rect 26388 5414 26400 5466
rect 26452 5414 26464 5466
rect 26516 5414 26528 5466
rect 26580 5414 34713 5466
rect 34765 5414 34777 5466
rect 34829 5414 34841 5466
rect 34893 5414 34905 5466
rect 34957 5414 34969 5466
rect 35021 5414 35027 5466
rect 1104 5392 35027 5414
rect 1104 4922 34868 4944
rect 1104 4870 5170 4922
rect 5222 4870 5234 4922
rect 5286 4870 5298 4922
rect 5350 4870 5362 4922
rect 5414 4870 5426 4922
rect 5478 4870 13611 4922
rect 13663 4870 13675 4922
rect 13727 4870 13739 4922
rect 13791 4870 13803 4922
rect 13855 4870 13867 4922
rect 13919 4870 22052 4922
rect 22104 4870 22116 4922
rect 22168 4870 22180 4922
rect 22232 4870 22244 4922
rect 22296 4870 22308 4922
rect 22360 4870 30493 4922
rect 30545 4870 30557 4922
rect 30609 4870 30621 4922
rect 30673 4870 30685 4922
rect 30737 4870 30749 4922
rect 30801 4870 34868 4922
rect 1104 4848 34868 4870
rect 1104 4378 35027 4400
rect 1104 4326 9390 4378
rect 9442 4326 9454 4378
rect 9506 4326 9518 4378
rect 9570 4326 9582 4378
rect 9634 4326 9646 4378
rect 9698 4326 17831 4378
rect 17883 4326 17895 4378
rect 17947 4326 17959 4378
rect 18011 4326 18023 4378
rect 18075 4326 18087 4378
rect 18139 4326 26272 4378
rect 26324 4326 26336 4378
rect 26388 4326 26400 4378
rect 26452 4326 26464 4378
rect 26516 4326 26528 4378
rect 26580 4326 34713 4378
rect 34765 4326 34777 4378
rect 34829 4326 34841 4378
rect 34893 4326 34905 4378
rect 34957 4326 34969 4378
rect 35021 4326 35027 4378
rect 1104 4304 35027 4326
rect 1104 3834 34868 3856
rect 1104 3782 5170 3834
rect 5222 3782 5234 3834
rect 5286 3782 5298 3834
rect 5350 3782 5362 3834
rect 5414 3782 5426 3834
rect 5478 3782 13611 3834
rect 13663 3782 13675 3834
rect 13727 3782 13739 3834
rect 13791 3782 13803 3834
rect 13855 3782 13867 3834
rect 13919 3782 22052 3834
rect 22104 3782 22116 3834
rect 22168 3782 22180 3834
rect 22232 3782 22244 3834
rect 22296 3782 22308 3834
rect 22360 3782 30493 3834
rect 30545 3782 30557 3834
rect 30609 3782 30621 3834
rect 30673 3782 30685 3834
rect 30737 3782 30749 3834
rect 30801 3782 34868 3834
rect 1104 3760 34868 3782
rect 1104 3290 35027 3312
rect 1104 3238 9390 3290
rect 9442 3238 9454 3290
rect 9506 3238 9518 3290
rect 9570 3238 9582 3290
rect 9634 3238 9646 3290
rect 9698 3238 17831 3290
rect 17883 3238 17895 3290
rect 17947 3238 17959 3290
rect 18011 3238 18023 3290
rect 18075 3238 18087 3290
rect 18139 3238 26272 3290
rect 26324 3238 26336 3290
rect 26388 3238 26400 3290
rect 26452 3238 26464 3290
rect 26516 3238 26528 3290
rect 26580 3238 34713 3290
rect 34765 3238 34777 3290
rect 34829 3238 34841 3290
rect 34893 3238 34905 3290
rect 34957 3238 34969 3290
rect 35021 3238 35027 3290
rect 1104 3216 35027 3238
rect 1104 2746 34868 2768
rect 1104 2694 5170 2746
rect 5222 2694 5234 2746
rect 5286 2694 5298 2746
rect 5350 2694 5362 2746
rect 5414 2694 5426 2746
rect 5478 2694 13611 2746
rect 13663 2694 13675 2746
rect 13727 2694 13739 2746
rect 13791 2694 13803 2746
rect 13855 2694 13867 2746
rect 13919 2694 22052 2746
rect 22104 2694 22116 2746
rect 22168 2694 22180 2746
rect 22232 2694 22244 2746
rect 22296 2694 22308 2746
rect 22360 2694 30493 2746
rect 30545 2694 30557 2746
rect 30609 2694 30621 2746
rect 30673 2694 30685 2746
rect 30737 2694 30749 2746
rect 30801 2694 34868 2746
rect 1104 2672 34868 2694
rect 28442 2592 28448 2644
rect 28500 2592 28506 2644
rect 31478 2592 31484 2644
rect 31536 2632 31542 2644
rect 34333 2635 34391 2641
rect 34333 2632 34345 2635
rect 31536 2604 34345 2632
rect 31536 2592 31542 2604
rect 34333 2601 34345 2604
rect 34379 2601 34391 2635
rect 34333 2595 34391 2601
rect 1670 2456 1676 2508
rect 1728 2456 1734 2508
rect 14 2388 20 2440
rect 72 2428 78 2440
rect 1397 2431 1455 2437
rect 1397 2428 1409 2431
rect 72 2400 1409 2428
rect 72 2388 78 2400
rect 1397 2397 1409 2400
rect 1443 2397 1455 2431
rect 1397 2391 1455 2397
rect 9122 2388 9128 2440
rect 9180 2388 9186 2440
rect 19610 2388 19616 2440
rect 19668 2388 19674 2440
rect 28350 2388 28356 2440
rect 28408 2428 28414 2440
rect 28629 2431 28687 2437
rect 28629 2428 28641 2431
rect 28408 2400 28641 2428
rect 28408 2388 28414 2400
rect 28629 2397 28641 2400
rect 28675 2397 28687 2431
rect 28629 2391 28687 2397
rect 34517 2431 34575 2437
rect 34517 2397 34529 2431
rect 34563 2428 34575 2431
rect 34563 2400 35204 2428
rect 34563 2397 34575 2400
rect 34517 2391 34575 2397
rect 35176 2304 35204 2400
rect 18782 2252 18788 2304
rect 18840 2292 18846 2304
rect 19337 2295 19395 2301
rect 19337 2292 19349 2295
rect 18840 2264 19349 2292
rect 18840 2252 18846 2264
rect 19337 2261 19349 2264
rect 19383 2261 19395 2295
rect 19337 2255 19395 2261
rect 35158 2252 35164 2304
rect 35216 2252 35222 2304
rect 1104 2202 35027 2224
rect 1104 2150 9390 2202
rect 9442 2150 9454 2202
rect 9506 2150 9518 2202
rect 9570 2150 9582 2202
rect 9634 2150 9646 2202
rect 9698 2150 17831 2202
rect 17883 2150 17895 2202
rect 17947 2150 17959 2202
rect 18011 2150 18023 2202
rect 18075 2150 18087 2202
rect 18139 2150 26272 2202
rect 26324 2150 26336 2202
rect 26388 2150 26400 2202
rect 26452 2150 26464 2202
rect 26516 2150 26528 2202
rect 26580 2150 34713 2202
rect 34765 2150 34777 2202
rect 34829 2150 34841 2202
rect 34893 2150 34905 2202
rect 34957 2150 34969 2202
rect 35021 2150 35027 2202
rect 1104 2128 35027 2150
<< via1 >>
rect 5170 39686 5222 39738
rect 5234 39686 5286 39738
rect 5298 39686 5350 39738
rect 5362 39686 5414 39738
rect 5426 39686 5478 39738
rect 13611 39686 13663 39738
rect 13675 39686 13727 39738
rect 13739 39686 13791 39738
rect 13803 39686 13855 39738
rect 13867 39686 13919 39738
rect 22052 39686 22104 39738
rect 22116 39686 22168 39738
rect 22180 39686 22232 39738
rect 22244 39686 22296 39738
rect 22308 39686 22360 39738
rect 30493 39686 30545 39738
rect 30557 39686 30609 39738
rect 30621 39686 30673 39738
rect 30685 39686 30737 39738
rect 30749 39686 30801 39738
rect 26424 39584 26476 39636
rect 35440 39584 35492 39636
rect 940 39380 992 39432
rect 7104 39380 7156 39432
rect 16764 39380 16816 39432
rect 34152 39355 34204 39364
rect 34152 39321 34161 39355
rect 34161 39321 34195 39355
rect 34195 39321 34204 39355
rect 34152 39312 34204 39321
rect 1584 39287 1636 39296
rect 1584 39253 1593 39287
rect 1593 39253 1627 39287
rect 1627 39253 1636 39287
rect 1584 39244 1636 39253
rect 16120 39244 16172 39296
rect 17592 39244 17644 39296
rect 9390 39142 9442 39194
rect 9454 39142 9506 39194
rect 9518 39142 9570 39194
rect 9582 39142 9634 39194
rect 9646 39142 9698 39194
rect 17831 39142 17883 39194
rect 17895 39142 17947 39194
rect 17959 39142 18011 39194
rect 18023 39142 18075 39194
rect 18087 39142 18139 39194
rect 26272 39142 26324 39194
rect 26336 39142 26388 39194
rect 26400 39142 26452 39194
rect 26464 39142 26516 39194
rect 26528 39142 26580 39194
rect 34713 39142 34765 39194
rect 34777 39142 34829 39194
rect 34841 39142 34893 39194
rect 34905 39142 34957 39194
rect 34969 39142 35021 39194
rect 5170 38598 5222 38650
rect 5234 38598 5286 38650
rect 5298 38598 5350 38650
rect 5362 38598 5414 38650
rect 5426 38598 5478 38650
rect 13611 38598 13663 38650
rect 13675 38598 13727 38650
rect 13739 38598 13791 38650
rect 13803 38598 13855 38650
rect 13867 38598 13919 38650
rect 22052 38598 22104 38650
rect 22116 38598 22168 38650
rect 22180 38598 22232 38650
rect 22244 38598 22296 38650
rect 22308 38598 22360 38650
rect 30493 38598 30545 38650
rect 30557 38598 30609 38650
rect 30621 38598 30673 38650
rect 30685 38598 30737 38650
rect 30749 38598 30801 38650
rect 9390 38054 9442 38106
rect 9454 38054 9506 38106
rect 9518 38054 9570 38106
rect 9582 38054 9634 38106
rect 9646 38054 9698 38106
rect 17831 38054 17883 38106
rect 17895 38054 17947 38106
rect 17959 38054 18011 38106
rect 18023 38054 18075 38106
rect 18087 38054 18139 38106
rect 26272 38054 26324 38106
rect 26336 38054 26388 38106
rect 26400 38054 26452 38106
rect 26464 38054 26516 38106
rect 26528 38054 26580 38106
rect 34713 38054 34765 38106
rect 34777 38054 34829 38106
rect 34841 38054 34893 38106
rect 34905 38054 34957 38106
rect 34969 38054 35021 38106
rect 5170 37510 5222 37562
rect 5234 37510 5286 37562
rect 5298 37510 5350 37562
rect 5362 37510 5414 37562
rect 5426 37510 5478 37562
rect 13611 37510 13663 37562
rect 13675 37510 13727 37562
rect 13739 37510 13791 37562
rect 13803 37510 13855 37562
rect 13867 37510 13919 37562
rect 22052 37510 22104 37562
rect 22116 37510 22168 37562
rect 22180 37510 22232 37562
rect 22244 37510 22296 37562
rect 22308 37510 22360 37562
rect 30493 37510 30545 37562
rect 30557 37510 30609 37562
rect 30621 37510 30673 37562
rect 30685 37510 30737 37562
rect 30749 37510 30801 37562
rect 9390 36966 9442 37018
rect 9454 36966 9506 37018
rect 9518 36966 9570 37018
rect 9582 36966 9634 37018
rect 9646 36966 9698 37018
rect 17831 36966 17883 37018
rect 17895 36966 17947 37018
rect 17959 36966 18011 37018
rect 18023 36966 18075 37018
rect 18087 36966 18139 37018
rect 26272 36966 26324 37018
rect 26336 36966 26388 37018
rect 26400 36966 26452 37018
rect 26464 36966 26516 37018
rect 26528 36966 26580 37018
rect 34713 36966 34765 37018
rect 34777 36966 34829 37018
rect 34841 36966 34893 37018
rect 34905 36966 34957 37018
rect 34969 36966 35021 37018
rect 5170 36422 5222 36474
rect 5234 36422 5286 36474
rect 5298 36422 5350 36474
rect 5362 36422 5414 36474
rect 5426 36422 5478 36474
rect 13611 36422 13663 36474
rect 13675 36422 13727 36474
rect 13739 36422 13791 36474
rect 13803 36422 13855 36474
rect 13867 36422 13919 36474
rect 22052 36422 22104 36474
rect 22116 36422 22168 36474
rect 22180 36422 22232 36474
rect 22244 36422 22296 36474
rect 22308 36422 22360 36474
rect 30493 36422 30545 36474
rect 30557 36422 30609 36474
rect 30621 36422 30673 36474
rect 30685 36422 30737 36474
rect 30749 36422 30801 36474
rect 9390 35878 9442 35930
rect 9454 35878 9506 35930
rect 9518 35878 9570 35930
rect 9582 35878 9634 35930
rect 9646 35878 9698 35930
rect 17831 35878 17883 35930
rect 17895 35878 17947 35930
rect 17959 35878 18011 35930
rect 18023 35878 18075 35930
rect 18087 35878 18139 35930
rect 26272 35878 26324 35930
rect 26336 35878 26388 35930
rect 26400 35878 26452 35930
rect 26464 35878 26516 35930
rect 26528 35878 26580 35930
rect 34713 35878 34765 35930
rect 34777 35878 34829 35930
rect 34841 35878 34893 35930
rect 34905 35878 34957 35930
rect 34969 35878 35021 35930
rect 5170 35334 5222 35386
rect 5234 35334 5286 35386
rect 5298 35334 5350 35386
rect 5362 35334 5414 35386
rect 5426 35334 5478 35386
rect 13611 35334 13663 35386
rect 13675 35334 13727 35386
rect 13739 35334 13791 35386
rect 13803 35334 13855 35386
rect 13867 35334 13919 35386
rect 22052 35334 22104 35386
rect 22116 35334 22168 35386
rect 22180 35334 22232 35386
rect 22244 35334 22296 35386
rect 22308 35334 22360 35386
rect 30493 35334 30545 35386
rect 30557 35334 30609 35386
rect 30621 35334 30673 35386
rect 30685 35334 30737 35386
rect 30749 35334 30801 35386
rect 9390 34790 9442 34842
rect 9454 34790 9506 34842
rect 9518 34790 9570 34842
rect 9582 34790 9634 34842
rect 9646 34790 9698 34842
rect 17831 34790 17883 34842
rect 17895 34790 17947 34842
rect 17959 34790 18011 34842
rect 18023 34790 18075 34842
rect 18087 34790 18139 34842
rect 26272 34790 26324 34842
rect 26336 34790 26388 34842
rect 26400 34790 26452 34842
rect 26464 34790 26516 34842
rect 26528 34790 26580 34842
rect 34713 34790 34765 34842
rect 34777 34790 34829 34842
rect 34841 34790 34893 34842
rect 34905 34790 34957 34842
rect 34969 34790 35021 34842
rect 5170 34246 5222 34298
rect 5234 34246 5286 34298
rect 5298 34246 5350 34298
rect 5362 34246 5414 34298
rect 5426 34246 5478 34298
rect 13611 34246 13663 34298
rect 13675 34246 13727 34298
rect 13739 34246 13791 34298
rect 13803 34246 13855 34298
rect 13867 34246 13919 34298
rect 22052 34246 22104 34298
rect 22116 34246 22168 34298
rect 22180 34246 22232 34298
rect 22244 34246 22296 34298
rect 22308 34246 22360 34298
rect 30493 34246 30545 34298
rect 30557 34246 30609 34298
rect 30621 34246 30673 34298
rect 30685 34246 30737 34298
rect 30749 34246 30801 34298
rect 25964 33940 26016 33992
rect 26884 33872 26936 33924
rect 26148 33804 26200 33856
rect 26792 33804 26844 33856
rect 9390 33702 9442 33754
rect 9454 33702 9506 33754
rect 9518 33702 9570 33754
rect 9582 33702 9634 33754
rect 9646 33702 9698 33754
rect 17831 33702 17883 33754
rect 17895 33702 17947 33754
rect 17959 33702 18011 33754
rect 18023 33702 18075 33754
rect 18087 33702 18139 33754
rect 26272 33702 26324 33754
rect 26336 33702 26388 33754
rect 26400 33702 26452 33754
rect 26464 33702 26516 33754
rect 26528 33702 26580 33754
rect 34713 33702 34765 33754
rect 34777 33702 34829 33754
rect 34841 33702 34893 33754
rect 34905 33702 34957 33754
rect 34969 33702 35021 33754
rect 26792 33600 26844 33652
rect 1584 33464 1636 33516
rect 23940 33507 23992 33516
rect 23940 33473 23949 33507
rect 23949 33473 23983 33507
rect 23983 33473 23992 33507
rect 23940 33464 23992 33473
rect 25504 33464 25556 33516
rect 23848 33396 23900 33448
rect 26148 33396 26200 33448
rect 26608 33396 26660 33448
rect 26976 33507 27028 33516
rect 26976 33473 26985 33507
rect 26985 33473 27019 33507
rect 27019 33473 27028 33507
rect 26976 33464 27028 33473
rect 29552 33464 29604 33516
rect 27068 33396 27120 33448
rect 27252 33396 27304 33448
rect 28356 33439 28408 33448
rect 28356 33405 28365 33439
rect 28365 33405 28399 33439
rect 28399 33405 28408 33439
rect 28356 33396 28408 33405
rect 26240 33371 26292 33380
rect 26240 33337 26249 33371
rect 26249 33337 26283 33371
rect 26283 33337 26292 33371
rect 26240 33328 26292 33337
rect 23480 33260 23532 33312
rect 24492 33260 24544 33312
rect 26332 33260 26384 33312
rect 27436 33328 27488 33380
rect 30196 33464 30248 33516
rect 30288 33464 30340 33516
rect 31024 33507 31076 33516
rect 31024 33473 31033 33507
rect 31033 33473 31067 33507
rect 31067 33473 31076 33507
rect 31024 33464 31076 33473
rect 32220 33464 32272 33516
rect 30012 33439 30064 33448
rect 30012 33405 30021 33439
rect 30021 33405 30055 33439
rect 30055 33405 30064 33439
rect 30012 33396 30064 33405
rect 31300 33328 31352 33380
rect 27160 33260 27212 33312
rect 29920 33303 29972 33312
rect 29920 33269 29929 33303
rect 29929 33269 29963 33303
rect 29963 33269 29972 33303
rect 29920 33260 29972 33269
rect 30104 33260 30156 33312
rect 30380 33260 30432 33312
rect 30840 33303 30892 33312
rect 30840 33269 30849 33303
rect 30849 33269 30883 33303
rect 30883 33269 30892 33303
rect 30840 33260 30892 33269
rect 5170 33158 5222 33210
rect 5234 33158 5286 33210
rect 5298 33158 5350 33210
rect 5362 33158 5414 33210
rect 5426 33158 5478 33210
rect 13611 33158 13663 33210
rect 13675 33158 13727 33210
rect 13739 33158 13791 33210
rect 13803 33158 13855 33210
rect 13867 33158 13919 33210
rect 22052 33158 22104 33210
rect 22116 33158 22168 33210
rect 22180 33158 22232 33210
rect 22244 33158 22296 33210
rect 22308 33158 22360 33210
rect 30493 33158 30545 33210
rect 30557 33158 30609 33210
rect 30621 33158 30673 33210
rect 30685 33158 30737 33210
rect 30749 33158 30801 33210
rect 23940 33056 23992 33108
rect 25596 33056 25648 33108
rect 27252 33056 27304 33108
rect 29552 33099 29604 33108
rect 29552 33065 29561 33099
rect 29561 33065 29595 33099
rect 29595 33065 29604 33099
rect 29552 33056 29604 33065
rect 26148 32988 26200 33040
rect 23388 32920 23440 32972
rect 23480 32852 23532 32904
rect 23940 32895 23992 32904
rect 23940 32861 23949 32895
rect 23949 32861 23983 32895
rect 23983 32861 23992 32895
rect 23940 32852 23992 32861
rect 24308 32852 24360 32904
rect 24492 32852 24544 32904
rect 26976 32988 27028 33040
rect 27160 32920 27212 32972
rect 26240 32895 26292 32904
rect 26240 32861 26249 32895
rect 26249 32861 26283 32895
rect 26283 32861 26292 32895
rect 26240 32852 26292 32861
rect 27344 32852 27396 32904
rect 29736 32895 29788 32904
rect 29736 32861 29745 32895
rect 29745 32861 29779 32895
rect 29779 32861 29788 32895
rect 29736 32852 29788 32861
rect 29920 32852 29972 32904
rect 31208 32895 31260 32904
rect 31208 32861 31217 32895
rect 31217 32861 31251 32895
rect 31251 32861 31260 32895
rect 31208 32852 31260 32861
rect 31300 32852 31352 32904
rect 30288 32784 30340 32836
rect 25688 32716 25740 32768
rect 25872 32759 25924 32768
rect 25872 32725 25881 32759
rect 25881 32725 25915 32759
rect 25915 32725 25924 32759
rect 25872 32716 25924 32725
rect 26148 32716 26200 32768
rect 27068 32759 27120 32768
rect 27068 32725 27077 32759
rect 27077 32725 27111 32759
rect 27111 32725 27120 32759
rect 27068 32716 27120 32725
rect 28908 32716 28960 32768
rect 29092 32716 29144 32768
rect 30012 32716 30064 32768
rect 9390 32614 9442 32666
rect 9454 32614 9506 32666
rect 9518 32614 9570 32666
rect 9582 32614 9634 32666
rect 9646 32614 9698 32666
rect 17831 32614 17883 32666
rect 17895 32614 17947 32666
rect 17959 32614 18011 32666
rect 18023 32614 18075 32666
rect 18087 32614 18139 32666
rect 26272 32614 26324 32666
rect 26336 32614 26388 32666
rect 26400 32614 26452 32666
rect 26464 32614 26516 32666
rect 26528 32614 26580 32666
rect 34713 32614 34765 32666
rect 34777 32614 34829 32666
rect 34841 32614 34893 32666
rect 34905 32614 34957 32666
rect 34969 32614 35021 32666
rect 18328 32376 18380 32428
rect 18696 32419 18748 32428
rect 18696 32385 18730 32419
rect 18730 32385 18748 32419
rect 18696 32376 18748 32385
rect 20536 32376 20588 32428
rect 18144 32308 18196 32360
rect 17132 32240 17184 32292
rect 19800 32283 19852 32292
rect 19800 32249 19809 32283
rect 19809 32249 19843 32283
rect 19843 32249 19852 32283
rect 20720 32351 20772 32360
rect 20720 32317 20729 32351
rect 20729 32317 20763 32351
rect 20763 32317 20772 32351
rect 20996 32419 21048 32428
rect 20996 32385 21005 32419
rect 21005 32385 21039 32419
rect 21039 32385 21048 32419
rect 20996 32376 21048 32385
rect 21732 32376 21784 32428
rect 23388 32376 23440 32428
rect 25780 32512 25832 32564
rect 25872 32512 25924 32564
rect 25964 32512 26016 32564
rect 25596 32444 25648 32496
rect 26608 32444 26660 32496
rect 26976 32555 27028 32564
rect 26976 32521 26985 32555
rect 26985 32521 27019 32555
rect 27019 32521 27028 32555
rect 26976 32512 27028 32521
rect 27160 32512 27212 32564
rect 26884 32444 26936 32496
rect 27436 32512 27488 32564
rect 28356 32512 28408 32564
rect 20720 32308 20772 32317
rect 19800 32240 19852 32249
rect 20444 32283 20496 32292
rect 20444 32249 20453 32283
rect 20453 32249 20487 32283
rect 20487 32249 20496 32283
rect 20444 32240 20496 32249
rect 25872 32308 25924 32360
rect 26240 32308 26292 32360
rect 25780 32240 25832 32292
rect 27436 32419 27488 32428
rect 27436 32385 27445 32419
rect 27445 32385 27479 32419
rect 27479 32385 27488 32419
rect 27436 32376 27488 32385
rect 29092 32419 29144 32428
rect 29092 32385 29121 32419
rect 29121 32385 29144 32419
rect 29920 32555 29972 32564
rect 29920 32521 29929 32555
rect 29929 32521 29963 32555
rect 29963 32521 29972 32555
rect 29920 32512 29972 32521
rect 30104 32555 30156 32564
rect 30104 32521 30113 32555
rect 30113 32521 30147 32555
rect 30147 32521 30156 32555
rect 30104 32512 30156 32521
rect 29460 32444 29512 32496
rect 30196 32444 30248 32496
rect 30840 32444 30892 32496
rect 29092 32376 29144 32385
rect 30012 32419 30064 32428
rect 30012 32385 30021 32419
rect 30021 32385 30055 32419
rect 30055 32385 30064 32419
rect 30012 32376 30064 32385
rect 31208 32376 31260 32428
rect 34888 32376 34940 32428
rect 17316 32172 17368 32224
rect 17776 32215 17828 32224
rect 17776 32181 17785 32215
rect 17785 32181 17819 32215
rect 17819 32181 17828 32215
rect 17776 32172 17828 32181
rect 20628 32172 20680 32224
rect 21180 32215 21232 32224
rect 21180 32181 21189 32215
rect 21189 32181 21223 32215
rect 21223 32181 21232 32215
rect 21180 32172 21232 32181
rect 21824 32215 21876 32224
rect 21824 32181 21833 32215
rect 21833 32181 21867 32215
rect 21867 32181 21876 32215
rect 21824 32172 21876 32181
rect 21916 32172 21968 32224
rect 25504 32172 25556 32224
rect 29460 32240 29512 32292
rect 26700 32215 26752 32224
rect 26700 32181 26709 32215
rect 26709 32181 26743 32215
rect 26743 32181 26752 32215
rect 26700 32172 26752 32181
rect 31116 32172 31168 32224
rect 31392 32172 31444 32224
rect 32036 32172 32088 32224
rect 5170 32070 5222 32122
rect 5234 32070 5286 32122
rect 5298 32070 5350 32122
rect 5362 32070 5414 32122
rect 5426 32070 5478 32122
rect 13611 32070 13663 32122
rect 13675 32070 13727 32122
rect 13739 32070 13791 32122
rect 13803 32070 13855 32122
rect 13867 32070 13919 32122
rect 22052 32070 22104 32122
rect 22116 32070 22168 32122
rect 22180 32070 22232 32122
rect 22244 32070 22296 32122
rect 22308 32070 22360 32122
rect 30493 32070 30545 32122
rect 30557 32070 30609 32122
rect 30621 32070 30673 32122
rect 30685 32070 30737 32122
rect 30749 32070 30801 32122
rect 18144 31968 18196 32020
rect 18696 31968 18748 32020
rect 19800 31968 19852 32020
rect 20444 31968 20496 32020
rect 20996 31968 21048 32020
rect 21180 31968 21232 32020
rect 21732 32011 21784 32020
rect 21732 31977 21741 32011
rect 21741 31977 21775 32011
rect 21775 31977 21784 32011
rect 21732 31968 21784 31977
rect 24308 31968 24360 32020
rect 27068 31968 27120 32020
rect 16672 31764 16724 31816
rect 17132 31764 17184 31816
rect 17316 31807 17368 31816
rect 17316 31773 17350 31807
rect 17350 31773 17368 31807
rect 17316 31764 17368 31773
rect 18512 31764 18564 31816
rect 18972 31807 19024 31816
rect 18972 31773 18981 31807
rect 18981 31773 19015 31807
rect 19015 31773 19024 31807
rect 18972 31764 19024 31773
rect 19800 31696 19852 31748
rect 16672 31628 16724 31680
rect 19524 31671 19576 31680
rect 19524 31637 19533 31671
rect 19533 31637 19567 31671
rect 19567 31637 19576 31671
rect 19524 31628 19576 31637
rect 19708 31671 19760 31680
rect 19708 31637 19717 31671
rect 19717 31637 19751 31671
rect 19751 31637 19760 31671
rect 19708 31628 19760 31637
rect 20168 31764 20220 31816
rect 20628 31900 20680 31952
rect 20904 31807 20956 31816
rect 20904 31773 20913 31807
rect 20913 31773 20947 31807
rect 20947 31773 20956 31807
rect 20904 31764 20956 31773
rect 20260 31628 20312 31680
rect 20352 31671 20404 31680
rect 20352 31637 20361 31671
rect 20361 31637 20395 31671
rect 20395 31637 20404 31671
rect 20352 31628 20404 31637
rect 20812 31628 20864 31680
rect 21824 31900 21876 31952
rect 26056 31900 26108 31952
rect 29736 31968 29788 32020
rect 31024 31968 31076 32020
rect 21456 31764 21508 31816
rect 21548 31807 21600 31816
rect 21548 31773 21557 31807
rect 21557 31773 21591 31807
rect 21591 31773 21600 31807
rect 21548 31764 21600 31773
rect 21824 31807 21876 31816
rect 21824 31773 21833 31807
rect 21833 31773 21867 31807
rect 21867 31773 21876 31807
rect 21824 31764 21876 31773
rect 21916 31764 21968 31816
rect 25872 31832 25924 31884
rect 26148 31875 26200 31884
rect 26148 31841 26157 31875
rect 26157 31841 26191 31875
rect 26191 31841 26200 31875
rect 26148 31832 26200 31841
rect 26700 31832 26752 31884
rect 27620 31832 27672 31884
rect 29460 31832 29512 31884
rect 30012 31832 30064 31884
rect 31392 31968 31444 32020
rect 23940 31764 23992 31816
rect 28908 31807 28960 31816
rect 28908 31773 28917 31807
rect 28917 31773 28951 31807
rect 28951 31773 28960 31807
rect 28908 31764 28960 31773
rect 31208 31764 31260 31816
rect 31668 31832 31720 31884
rect 32220 31875 32272 31884
rect 32220 31841 32229 31875
rect 32229 31841 32263 31875
rect 32263 31841 32272 31875
rect 32220 31832 32272 31841
rect 31852 31807 31904 31816
rect 31852 31773 31861 31807
rect 31861 31773 31895 31807
rect 31895 31773 31904 31807
rect 31852 31764 31904 31773
rect 32036 31807 32088 31816
rect 32036 31773 32059 31807
rect 32059 31773 32088 31807
rect 32036 31764 32088 31773
rect 21916 31671 21968 31680
rect 21916 31637 21925 31671
rect 21925 31637 21959 31671
rect 21959 31637 21968 31671
rect 21916 31628 21968 31637
rect 30288 31671 30340 31680
rect 30288 31637 30297 31671
rect 30297 31637 30331 31671
rect 30331 31637 30340 31671
rect 30288 31628 30340 31637
rect 32128 31628 32180 31680
rect 9390 31526 9442 31578
rect 9454 31526 9506 31578
rect 9518 31526 9570 31578
rect 9582 31526 9634 31578
rect 9646 31526 9698 31578
rect 17831 31526 17883 31578
rect 17895 31526 17947 31578
rect 17959 31526 18011 31578
rect 18023 31526 18075 31578
rect 18087 31526 18139 31578
rect 26272 31526 26324 31578
rect 26336 31526 26388 31578
rect 26400 31526 26452 31578
rect 26464 31526 26516 31578
rect 26528 31526 26580 31578
rect 34713 31526 34765 31578
rect 34777 31526 34829 31578
rect 34841 31526 34893 31578
rect 34905 31526 34957 31578
rect 34969 31526 35021 31578
rect 18236 31467 18288 31476
rect 18236 31433 18245 31467
rect 18245 31433 18279 31467
rect 18279 31433 18288 31467
rect 18236 31424 18288 31433
rect 18880 31424 18932 31476
rect 18972 31424 19024 31476
rect 17684 31356 17736 31408
rect 20628 31424 20680 31476
rect 20996 31467 21048 31476
rect 20996 31433 21005 31467
rect 21005 31433 21039 31467
rect 21039 31433 21048 31467
rect 20996 31424 21048 31433
rect 23388 31424 23440 31476
rect 30288 31424 30340 31476
rect 16764 31288 16816 31340
rect 18420 31331 18472 31340
rect 18420 31297 18429 31331
rect 18429 31297 18463 31331
rect 18463 31297 18472 31331
rect 18420 31288 18472 31297
rect 19708 31288 19760 31340
rect 16672 31263 16724 31272
rect 16672 31229 16681 31263
rect 16681 31229 16715 31263
rect 16715 31229 16724 31263
rect 16672 31220 16724 31229
rect 18328 31220 18380 31272
rect 20168 31331 20220 31340
rect 20168 31297 20177 31331
rect 20177 31297 20211 31331
rect 20211 31297 20220 31331
rect 20168 31288 20220 31297
rect 20260 31288 20312 31340
rect 20444 31356 20496 31408
rect 20720 31356 20772 31408
rect 21916 31356 21968 31408
rect 24492 31356 24544 31408
rect 21548 31288 21600 31340
rect 23296 31331 23348 31340
rect 23296 31297 23305 31331
rect 23305 31297 23339 31331
rect 23339 31297 23348 31331
rect 23296 31288 23348 31297
rect 20720 31263 20772 31272
rect 20720 31229 20729 31263
rect 20729 31229 20763 31263
rect 20763 31229 20772 31263
rect 20720 31220 20772 31229
rect 21272 31220 21324 31272
rect 21824 31220 21876 31272
rect 27436 31288 27488 31340
rect 20352 31152 20404 31204
rect 28816 31288 28868 31340
rect 31116 31356 31168 31408
rect 30748 31288 30800 31340
rect 31392 31288 31444 31340
rect 31668 31356 31720 31408
rect 31944 31288 31996 31340
rect 32680 31288 32732 31340
rect 30380 31152 30432 31204
rect 17960 31084 18012 31136
rect 19156 31084 19208 31136
rect 19524 31084 19576 31136
rect 19984 31127 20036 31136
rect 19984 31093 19993 31127
rect 19993 31093 20027 31127
rect 20027 31093 20036 31127
rect 19984 31084 20036 31093
rect 20444 31084 20496 31136
rect 24676 31084 24728 31136
rect 24768 31127 24820 31136
rect 24768 31093 24777 31127
rect 24777 31093 24811 31127
rect 24811 31093 24820 31127
rect 24768 31084 24820 31093
rect 25504 31127 25556 31136
rect 25504 31093 25513 31127
rect 25513 31093 25547 31127
rect 25547 31093 25556 31127
rect 25504 31084 25556 31093
rect 27988 31084 28040 31136
rect 28080 31127 28132 31136
rect 28080 31093 28089 31127
rect 28089 31093 28123 31127
rect 28123 31093 28132 31127
rect 28080 31084 28132 31093
rect 29828 31084 29880 31136
rect 30104 31127 30156 31136
rect 30104 31093 30113 31127
rect 30113 31093 30147 31127
rect 30147 31093 30156 31127
rect 30104 31084 30156 31093
rect 30932 31127 30984 31136
rect 30932 31093 30941 31127
rect 30941 31093 30975 31127
rect 30975 31093 30984 31127
rect 30932 31084 30984 31093
rect 31024 31084 31076 31136
rect 31300 31084 31352 31136
rect 5170 30982 5222 31034
rect 5234 30982 5286 31034
rect 5298 30982 5350 31034
rect 5362 30982 5414 31034
rect 5426 30982 5478 31034
rect 13611 30982 13663 31034
rect 13675 30982 13727 31034
rect 13739 30982 13791 31034
rect 13803 30982 13855 31034
rect 13867 30982 13919 31034
rect 22052 30982 22104 31034
rect 22116 30982 22168 31034
rect 22180 30982 22232 31034
rect 22244 30982 22296 31034
rect 22308 30982 22360 31034
rect 30493 30982 30545 31034
rect 30557 30982 30609 31034
rect 30621 30982 30673 31034
rect 30685 30982 30737 31034
rect 30749 30982 30801 31034
rect 16764 30923 16816 30932
rect 16764 30889 16773 30923
rect 16773 30889 16807 30923
rect 16807 30889 16816 30923
rect 16764 30880 16816 30889
rect 17592 30923 17644 30932
rect 17592 30889 17601 30923
rect 17601 30889 17635 30923
rect 17635 30889 17644 30923
rect 17592 30880 17644 30889
rect 17684 30880 17736 30932
rect 17132 30719 17184 30728
rect 17132 30685 17141 30719
rect 17141 30685 17175 30719
rect 17175 30685 17184 30719
rect 17132 30676 17184 30685
rect 18420 30880 18472 30932
rect 18512 30812 18564 30864
rect 18880 30812 18932 30864
rect 19064 30744 19116 30796
rect 18696 30676 18748 30728
rect 17960 30608 18012 30660
rect 18880 30676 18932 30728
rect 19340 30676 19392 30728
rect 19524 30719 19576 30728
rect 19524 30685 19533 30719
rect 19533 30685 19567 30719
rect 19567 30685 19576 30719
rect 19524 30676 19576 30685
rect 19800 30812 19852 30864
rect 19984 30744 20036 30796
rect 20260 30744 20312 30796
rect 23388 30880 23440 30932
rect 24676 30923 24728 30932
rect 24676 30889 24685 30923
rect 24685 30889 24719 30923
rect 24719 30889 24728 30923
rect 24676 30880 24728 30889
rect 24492 30812 24544 30864
rect 22652 30608 22704 30660
rect 23664 30719 23716 30728
rect 23664 30685 23673 30719
rect 23673 30685 23707 30719
rect 23707 30685 23716 30719
rect 23664 30676 23716 30685
rect 23848 30676 23900 30728
rect 24216 30676 24268 30728
rect 24768 30676 24820 30728
rect 25504 30880 25556 30932
rect 27344 30880 27396 30932
rect 17500 30540 17552 30592
rect 18236 30540 18288 30592
rect 19248 30540 19300 30592
rect 23112 30540 23164 30592
rect 23204 30540 23256 30592
rect 24308 30608 24360 30660
rect 23480 30583 23532 30592
rect 23480 30549 23489 30583
rect 23489 30549 23523 30583
rect 23523 30549 23532 30583
rect 23480 30540 23532 30549
rect 23572 30540 23624 30592
rect 25412 30676 25464 30728
rect 25596 30676 25648 30728
rect 26884 30744 26936 30796
rect 27988 30812 28040 30864
rect 28172 30787 28224 30796
rect 28172 30753 28181 30787
rect 28181 30753 28215 30787
rect 28215 30753 28224 30787
rect 28172 30744 28224 30753
rect 25780 30719 25832 30728
rect 25780 30685 25789 30719
rect 25789 30685 25823 30719
rect 25823 30685 25832 30719
rect 25780 30676 25832 30685
rect 24952 30608 25004 30660
rect 26608 30719 26660 30728
rect 26608 30685 26617 30719
rect 26617 30685 26651 30719
rect 26651 30685 26660 30719
rect 26608 30676 26660 30685
rect 27436 30719 27488 30728
rect 27436 30685 27445 30719
rect 27445 30685 27479 30719
rect 27479 30685 27488 30719
rect 27436 30676 27488 30685
rect 27528 30676 27580 30728
rect 27712 30719 27764 30728
rect 27712 30685 27721 30719
rect 27721 30685 27755 30719
rect 27755 30685 27764 30719
rect 27712 30676 27764 30685
rect 27804 30676 27856 30728
rect 31024 30880 31076 30932
rect 31668 30880 31720 30932
rect 32680 30923 32732 30932
rect 32680 30889 32689 30923
rect 32689 30889 32723 30923
rect 32723 30889 32732 30923
rect 32680 30880 32732 30889
rect 32128 30812 32180 30864
rect 28816 30719 28868 30728
rect 28816 30685 28825 30719
rect 28825 30685 28859 30719
rect 28859 30685 28868 30719
rect 28816 30676 28868 30685
rect 29552 30719 29604 30728
rect 29552 30685 29561 30719
rect 29561 30685 29595 30719
rect 29595 30685 29604 30719
rect 29552 30676 29604 30685
rect 29828 30719 29880 30728
rect 29828 30685 29862 30719
rect 29862 30685 29880 30719
rect 29828 30676 29880 30685
rect 25688 30540 25740 30592
rect 26884 30540 26936 30592
rect 27896 30540 27948 30592
rect 28172 30540 28224 30592
rect 28540 30583 28592 30592
rect 28540 30549 28549 30583
rect 28549 30549 28583 30583
rect 28583 30549 28592 30583
rect 28540 30540 28592 30549
rect 30012 30540 30064 30592
rect 30656 30540 30708 30592
rect 31392 30608 31444 30660
rect 34152 30540 34204 30592
rect 9390 30438 9442 30490
rect 9454 30438 9506 30490
rect 9518 30438 9570 30490
rect 9582 30438 9634 30490
rect 9646 30438 9698 30490
rect 17831 30438 17883 30490
rect 17895 30438 17947 30490
rect 17959 30438 18011 30490
rect 18023 30438 18075 30490
rect 18087 30438 18139 30490
rect 26272 30438 26324 30490
rect 26336 30438 26388 30490
rect 26400 30438 26452 30490
rect 26464 30438 26516 30490
rect 26528 30438 26580 30490
rect 34713 30438 34765 30490
rect 34777 30438 34829 30490
rect 34841 30438 34893 30490
rect 34905 30438 34957 30490
rect 34969 30438 35021 30490
rect 17592 30336 17644 30388
rect 18236 30268 18288 30320
rect 19064 30336 19116 30388
rect 20260 30336 20312 30388
rect 23112 30336 23164 30388
rect 23388 30336 23440 30388
rect 25780 30336 25832 30388
rect 19524 30268 19576 30320
rect 940 29996 992 30048
rect 16396 29996 16448 30048
rect 16488 30039 16540 30048
rect 16488 30005 16497 30039
rect 16497 30005 16531 30039
rect 16531 30005 16540 30039
rect 16488 29996 16540 30005
rect 16764 30200 16816 30252
rect 18328 30243 18380 30252
rect 18328 30209 18337 30243
rect 18337 30209 18371 30243
rect 18371 30209 18380 30243
rect 18328 30200 18380 30209
rect 16672 30175 16724 30184
rect 16672 30141 16681 30175
rect 16681 30141 16715 30175
rect 16715 30141 16724 30175
rect 16672 30132 16724 30141
rect 19156 30200 19208 30252
rect 19248 30243 19300 30252
rect 19248 30209 19257 30243
rect 19257 30209 19291 30243
rect 19291 30209 19300 30243
rect 19248 30200 19300 30209
rect 20260 30243 20312 30252
rect 20260 30209 20269 30243
rect 20269 30209 20303 30243
rect 20303 30209 20312 30243
rect 20260 30200 20312 30209
rect 20444 30243 20496 30252
rect 20444 30209 20453 30243
rect 20453 30209 20487 30243
rect 20487 30209 20496 30243
rect 20444 30200 20496 30209
rect 20812 30200 20864 30252
rect 20904 30243 20956 30252
rect 20904 30209 20913 30243
rect 20913 30209 20947 30243
rect 20947 30209 20956 30243
rect 20904 30200 20956 30209
rect 21180 30200 21232 30252
rect 26608 30336 26660 30388
rect 27528 30336 27580 30388
rect 20536 30132 20588 30184
rect 20996 30175 21048 30184
rect 20996 30141 21005 30175
rect 21005 30141 21039 30175
rect 21039 30141 21048 30175
rect 20996 30132 21048 30141
rect 20352 30064 20404 30116
rect 20628 30107 20680 30116
rect 20628 30073 20637 30107
rect 20637 30073 20671 30107
rect 20671 30073 20680 30107
rect 20628 30064 20680 30073
rect 23388 30200 23440 30252
rect 24032 30200 24084 30252
rect 25136 30243 25188 30252
rect 25136 30209 25145 30243
rect 25145 30209 25179 30243
rect 25179 30209 25188 30243
rect 25136 30200 25188 30209
rect 25320 30243 25372 30252
rect 25320 30209 25329 30243
rect 25329 30209 25363 30243
rect 25363 30209 25372 30243
rect 25320 30200 25372 30209
rect 25596 30200 25648 30252
rect 25688 30243 25740 30252
rect 25688 30209 25697 30243
rect 25697 30209 25731 30243
rect 25731 30209 25740 30243
rect 25688 30200 25740 30209
rect 24952 30132 25004 30184
rect 26332 30243 26384 30252
rect 26332 30209 26341 30243
rect 26341 30209 26375 30243
rect 26375 30209 26384 30243
rect 26332 30200 26384 30209
rect 26608 30200 26660 30252
rect 21548 30064 21600 30116
rect 26884 30132 26936 30184
rect 17040 29996 17092 30048
rect 19156 30039 19208 30048
rect 19156 30005 19165 30039
rect 19165 30005 19199 30039
rect 19199 30005 19208 30039
rect 19156 29996 19208 30005
rect 20076 29996 20128 30048
rect 21272 29996 21324 30048
rect 24676 30039 24728 30048
rect 24676 30005 24685 30039
rect 24685 30005 24719 30039
rect 24719 30005 24728 30039
rect 24676 29996 24728 30005
rect 26700 30039 26752 30048
rect 26700 30005 26709 30039
rect 26709 30005 26743 30039
rect 26743 30005 26752 30039
rect 26700 29996 26752 30005
rect 27528 30200 27580 30252
rect 27620 30243 27672 30252
rect 27620 30209 27629 30243
rect 27629 30209 27663 30243
rect 27663 30209 27672 30243
rect 27620 30200 27672 30209
rect 27804 30243 27856 30252
rect 27804 30209 27813 30243
rect 27813 30209 27847 30243
rect 27847 30209 27856 30243
rect 27804 30200 27856 30209
rect 27896 30200 27948 30252
rect 28080 30200 28132 30252
rect 28264 30175 28316 30184
rect 28264 30141 28273 30175
rect 28273 30141 28307 30175
rect 28307 30141 28316 30175
rect 28264 30132 28316 30141
rect 28540 30243 28592 30252
rect 28540 30209 28549 30243
rect 28549 30209 28583 30243
rect 28583 30209 28592 30243
rect 28540 30200 28592 30209
rect 30104 30336 30156 30388
rect 30932 30336 30984 30388
rect 31392 30379 31444 30388
rect 31392 30345 31401 30379
rect 31401 30345 31435 30379
rect 31435 30345 31444 30379
rect 31392 30336 31444 30345
rect 30012 30200 30064 30252
rect 27988 30064 28040 30116
rect 28540 30064 28592 30116
rect 28632 30064 28684 30116
rect 30656 30243 30708 30252
rect 30656 30209 30665 30243
rect 30665 30209 30699 30243
rect 30699 30209 30708 30243
rect 30656 30200 30708 30209
rect 31852 30243 31904 30252
rect 31852 30209 31861 30243
rect 31861 30209 31895 30243
rect 31895 30209 31904 30243
rect 31852 30200 31904 30209
rect 27436 29996 27488 30048
rect 28172 30039 28224 30048
rect 28172 30005 28181 30039
rect 28181 30005 28215 30039
rect 28215 30005 28224 30039
rect 28172 29996 28224 30005
rect 28448 29996 28500 30048
rect 31208 30064 31260 30116
rect 29828 30039 29880 30048
rect 29828 30005 29837 30039
rect 29837 30005 29871 30039
rect 29871 30005 29880 30039
rect 29828 29996 29880 30005
rect 31576 29996 31628 30048
rect 5170 29894 5222 29946
rect 5234 29894 5286 29946
rect 5298 29894 5350 29946
rect 5362 29894 5414 29946
rect 5426 29894 5478 29946
rect 13611 29894 13663 29946
rect 13675 29894 13727 29946
rect 13739 29894 13791 29946
rect 13803 29894 13855 29946
rect 13867 29894 13919 29946
rect 22052 29894 22104 29946
rect 22116 29894 22168 29946
rect 22180 29894 22232 29946
rect 22244 29894 22296 29946
rect 22308 29894 22360 29946
rect 30493 29894 30545 29946
rect 30557 29894 30609 29946
rect 30621 29894 30673 29946
rect 30685 29894 30737 29946
rect 30749 29894 30801 29946
rect 16488 29792 16540 29844
rect 16764 29792 16816 29844
rect 17132 29792 17184 29844
rect 18328 29792 18380 29844
rect 19156 29792 19208 29844
rect 19248 29792 19300 29844
rect 17592 29699 17644 29708
rect 17592 29665 17601 29699
rect 17601 29665 17635 29699
rect 17635 29665 17644 29699
rect 17592 29656 17644 29665
rect 18604 29631 18656 29640
rect 18604 29597 18613 29631
rect 18613 29597 18647 29631
rect 18647 29597 18656 29631
rect 18604 29588 18656 29597
rect 18696 29631 18748 29640
rect 18696 29597 18705 29631
rect 18705 29597 18739 29631
rect 18739 29597 18748 29631
rect 18696 29588 18748 29597
rect 18880 29631 18932 29640
rect 18880 29597 18889 29631
rect 18889 29597 18923 29631
rect 18923 29597 18932 29631
rect 18880 29588 18932 29597
rect 19892 29724 19944 29776
rect 20536 29724 20588 29776
rect 20076 29656 20128 29708
rect 20352 29699 20404 29708
rect 20352 29665 20361 29699
rect 20361 29665 20395 29699
rect 20395 29665 20404 29699
rect 20352 29656 20404 29665
rect 20904 29792 20956 29844
rect 21272 29792 21324 29844
rect 21548 29792 21600 29844
rect 22652 29835 22704 29844
rect 22652 29801 22661 29835
rect 22661 29801 22695 29835
rect 22695 29801 22704 29835
rect 22652 29792 22704 29801
rect 23388 29792 23440 29844
rect 23480 29792 23532 29844
rect 24032 29835 24084 29844
rect 24032 29801 24041 29835
rect 24041 29801 24075 29835
rect 24075 29801 24084 29835
rect 24032 29792 24084 29801
rect 24216 29835 24268 29844
rect 24216 29801 24225 29835
rect 24225 29801 24259 29835
rect 24259 29801 24268 29835
rect 24216 29792 24268 29801
rect 24676 29792 24728 29844
rect 24952 29835 25004 29844
rect 24952 29801 24961 29835
rect 24961 29801 24995 29835
rect 24995 29801 25004 29835
rect 24952 29792 25004 29801
rect 25136 29835 25188 29844
rect 25136 29801 25145 29835
rect 25145 29801 25179 29835
rect 25179 29801 25188 29835
rect 25136 29792 25188 29801
rect 25320 29792 25372 29844
rect 20168 29520 20220 29572
rect 17408 29452 17460 29504
rect 20812 29631 20864 29640
rect 20812 29597 20821 29631
rect 20821 29597 20855 29631
rect 20855 29597 20864 29631
rect 20812 29588 20864 29597
rect 21456 29631 21508 29640
rect 21456 29597 21465 29631
rect 21465 29597 21499 29631
rect 21499 29597 21508 29631
rect 21456 29588 21508 29597
rect 23204 29724 23256 29776
rect 22836 29631 22888 29640
rect 22836 29597 22845 29631
rect 22845 29597 22879 29631
rect 22879 29597 22888 29631
rect 22836 29588 22888 29597
rect 23664 29656 23716 29708
rect 23572 29588 23624 29640
rect 20352 29452 20404 29504
rect 26608 29792 26660 29844
rect 27712 29792 27764 29844
rect 27896 29792 27948 29844
rect 27988 29792 28040 29844
rect 28172 29792 28224 29844
rect 28632 29792 28684 29844
rect 25688 29631 25740 29640
rect 25688 29597 25696 29631
rect 25696 29597 25730 29631
rect 25730 29597 25740 29631
rect 25688 29588 25740 29597
rect 25780 29631 25832 29640
rect 25780 29597 25789 29631
rect 25789 29597 25823 29631
rect 25823 29597 25832 29631
rect 25780 29588 25832 29597
rect 26700 29588 26752 29640
rect 27436 29631 27488 29640
rect 27436 29597 27445 29631
rect 27445 29597 27479 29631
rect 27479 29597 27488 29631
rect 27436 29588 27488 29597
rect 29552 29699 29604 29708
rect 29552 29665 29561 29699
rect 29561 29665 29595 29699
rect 29595 29665 29604 29699
rect 29552 29656 29604 29665
rect 29828 29631 29880 29640
rect 29828 29597 29862 29631
rect 29862 29597 29880 29631
rect 25504 29563 25556 29572
rect 25504 29529 25513 29563
rect 25513 29529 25547 29563
rect 25547 29529 25556 29563
rect 25504 29520 25556 29529
rect 28908 29520 28960 29572
rect 29828 29588 29880 29597
rect 31944 29792 31996 29844
rect 31576 29631 31628 29640
rect 31576 29597 31610 29631
rect 31610 29597 31628 29631
rect 31576 29588 31628 29597
rect 27804 29452 27856 29504
rect 28632 29452 28684 29504
rect 30840 29452 30892 29504
rect 31576 29452 31628 29504
rect 32404 29452 32456 29504
rect 9390 29350 9442 29402
rect 9454 29350 9506 29402
rect 9518 29350 9570 29402
rect 9582 29350 9634 29402
rect 9646 29350 9698 29402
rect 17831 29350 17883 29402
rect 17895 29350 17947 29402
rect 17959 29350 18011 29402
rect 18023 29350 18075 29402
rect 18087 29350 18139 29402
rect 26272 29350 26324 29402
rect 26336 29350 26388 29402
rect 26400 29350 26452 29402
rect 26464 29350 26516 29402
rect 26528 29350 26580 29402
rect 34713 29350 34765 29402
rect 34777 29350 34829 29402
rect 34841 29350 34893 29402
rect 34905 29350 34957 29402
rect 34969 29350 35021 29402
rect 18604 29248 18656 29300
rect 20444 29248 20496 29300
rect 20628 29248 20680 29300
rect 20996 29248 21048 29300
rect 22836 29248 22888 29300
rect 26884 29248 26936 29300
rect 28264 29248 28316 29300
rect 28908 29291 28960 29300
rect 28908 29257 28917 29291
rect 28917 29257 28951 29291
rect 28951 29257 28960 29291
rect 28908 29248 28960 29257
rect 17408 29180 17460 29232
rect 19892 29180 19944 29232
rect 16396 29044 16448 29096
rect 17776 29112 17828 29164
rect 20076 29155 20128 29164
rect 20076 29121 20105 29155
rect 20105 29121 20128 29155
rect 18420 29044 18472 29096
rect 20076 29112 20128 29121
rect 20260 29112 20312 29164
rect 20996 29112 21048 29164
rect 23848 29180 23900 29232
rect 20720 29044 20772 29096
rect 20904 29087 20956 29096
rect 20904 29053 20913 29087
rect 20913 29053 20947 29087
rect 20947 29053 20956 29087
rect 20904 29044 20956 29053
rect 21548 29044 21600 29096
rect 23020 29112 23072 29164
rect 23480 29112 23532 29164
rect 25044 29155 25096 29164
rect 25044 29121 25053 29155
rect 25053 29121 25087 29155
rect 25087 29121 25096 29155
rect 25044 29112 25096 29121
rect 28264 29155 28316 29164
rect 28264 29121 28273 29155
rect 28273 29121 28307 29155
rect 28307 29121 28316 29155
rect 28264 29112 28316 29121
rect 20260 29019 20312 29028
rect 20260 28985 20269 29019
rect 20269 28985 20303 29019
rect 20303 28985 20312 29019
rect 20260 28976 20312 28985
rect 20812 28976 20864 29028
rect 28632 29155 28684 29164
rect 28632 29121 28641 29155
rect 28641 29121 28675 29155
rect 28675 29121 28684 29155
rect 28632 29112 28684 29121
rect 31208 29044 31260 29096
rect 32404 29044 32456 29096
rect 28540 28976 28592 29028
rect 17040 28951 17092 28960
rect 17040 28917 17049 28951
rect 17049 28917 17083 28951
rect 17083 28917 17092 28951
rect 17040 28908 17092 28917
rect 21548 28951 21600 28960
rect 21548 28917 21557 28951
rect 21557 28917 21591 28951
rect 21591 28917 21600 28951
rect 21548 28908 21600 28917
rect 25136 28951 25188 28960
rect 25136 28917 25145 28951
rect 25145 28917 25179 28951
rect 25179 28917 25188 28951
rect 25136 28908 25188 28917
rect 31852 28908 31904 28960
rect 5170 28806 5222 28858
rect 5234 28806 5286 28858
rect 5298 28806 5350 28858
rect 5362 28806 5414 28858
rect 5426 28806 5478 28858
rect 13611 28806 13663 28858
rect 13675 28806 13727 28858
rect 13739 28806 13791 28858
rect 13803 28806 13855 28858
rect 13867 28806 13919 28858
rect 22052 28806 22104 28858
rect 22116 28806 22168 28858
rect 22180 28806 22232 28858
rect 22244 28806 22296 28858
rect 22308 28806 22360 28858
rect 30493 28806 30545 28858
rect 30557 28806 30609 28858
rect 30621 28806 30673 28858
rect 30685 28806 30737 28858
rect 30749 28806 30801 28858
rect 16672 28704 16724 28756
rect 17776 28747 17828 28756
rect 17776 28713 17785 28747
rect 17785 28713 17819 28747
rect 17819 28713 17828 28747
rect 17776 28704 17828 28713
rect 18328 28704 18380 28756
rect 18880 28704 18932 28756
rect 20720 28704 20772 28756
rect 21456 28704 21508 28756
rect 23664 28747 23716 28756
rect 23664 28713 23673 28747
rect 23673 28713 23707 28747
rect 23707 28713 23716 28747
rect 23664 28704 23716 28713
rect 18236 28543 18288 28552
rect 18236 28509 18245 28543
rect 18245 28509 18279 28543
rect 18279 28509 18288 28543
rect 18236 28500 18288 28509
rect 16856 28432 16908 28484
rect 18696 28500 18748 28552
rect 20628 28500 20680 28552
rect 18420 28475 18472 28484
rect 18420 28441 18429 28475
rect 18429 28441 18463 28475
rect 18463 28441 18472 28475
rect 18420 28432 18472 28441
rect 21456 28500 21508 28552
rect 21548 28500 21600 28552
rect 17500 28364 17552 28416
rect 21088 28432 21140 28484
rect 23020 28543 23072 28552
rect 23020 28509 23029 28543
rect 23029 28509 23063 28543
rect 23063 28509 23072 28543
rect 23020 28500 23072 28509
rect 25044 28636 25096 28688
rect 25136 28636 25188 28688
rect 25780 28704 25832 28756
rect 27896 28704 27948 28756
rect 25504 28611 25556 28620
rect 25504 28577 25513 28611
rect 25513 28577 25547 28611
rect 25547 28577 25556 28611
rect 25504 28568 25556 28577
rect 27712 28568 27764 28620
rect 29000 28568 29052 28620
rect 25136 28543 25188 28552
rect 25136 28509 25145 28543
rect 25145 28509 25179 28543
rect 25179 28509 25188 28543
rect 25136 28500 25188 28509
rect 25320 28543 25372 28552
rect 25320 28509 25329 28543
rect 25329 28509 25363 28543
rect 25363 28509 25372 28543
rect 25320 28500 25372 28509
rect 24032 28475 24084 28484
rect 24032 28441 24041 28475
rect 24041 28441 24075 28475
rect 24075 28441 24084 28475
rect 24032 28432 24084 28441
rect 25688 28543 25740 28552
rect 25688 28509 25697 28543
rect 25697 28509 25731 28543
rect 25731 28509 25740 28543
rect 25688 28500 25740 28509
rect 25504 28432 25556 28484
rect 27344 28543 27396 28552
rect 27344 28509 27353 28543
rect 27353 28509 27387 28543
rect 27387 28509 27396 28543
rect 27344 28500 27396 28509
rect 31024 28500 31076 28552
rect 31852 28543 31904 28552
rect 31852 28509 31886 28543
rect 31886 28509 31904 28543
rect 31852 28500 31904 28509
rect 30380 28432 30432 28484
rect 18604 28364 18656 28416
rect 23112 28407 23164 28416
rect 23112 28373 23121 28407
rect 23121 28373 23155 28407
rect 23155 28373 23164 28407
rect 23112 28364 23164 28373
rect 23204 28364 23256 28416
rect 23848 28407 23900 28416
rect 23848 28373 23865 28407
rect 23865 28373 23900 28407
rect 23848 28364 23900 28373
rect 27160 28364 27212 28416
rect 27528 28407 27580 28416
rect 27528 28373 27537 28407
rect 27537 28373 27571 28407
rect 27571 28373 27580 28407
rect 27528 28364 27580 28373
rect 27620 28364 27672 28416
rect 27896 28364 27948 28416
rect 28080 28407 28132 28416
rect 28080 28373 28089 28407
rect 28089 28373 28123 28407
rect 28123 28373 28132 28407
rect 28080 28364 28132 28373
rect 31392 28407 31444 28416
rect 31392 28373 31401 28407
rect 31401 28373 31435 28407
rect 31435 28373 31444 28407
rect 31392 28364 31444 28373
rect 32128 28364 32180 28416
rect 9390 28262 9442 28314
rect 9454 28262 9506 28314
rect 9518 28262 9570 28314
rect 9582 28262 9634 28314
rect 9646 28262 9698 28314
rect 17831 28262 17883 28314
rect 17895 28262 17947 28314
rect 17959 28262 18011 28314
rect 18023 28262 18075 28314
rect 18087 28262 18139 28314
rect 26272 28262 26324 28314
rect 26336 28262 26388 28314
rect 26400 28262 26452 28314
rect 26464 28262 26516 28314
rect 26528 28262 26580 28314
rect 34713 28262 34765 28314
rect 34777 28262 34829 28314
rect 34841 28262 34893 28314
rect 34905 28262 34957 28314
rect 34969 28262 35021 28314
rect 16856 28203 16908 28212
rect 16856 28169 16865 28203
rect 16865 28169 16899 28203
rect 16899 28169 16908 28203
rect 16856 28160 16908 28169
rect 18420 28160 18472 28212
rect 23664 28203 23716 28212
rect 23664 28169 23673 28203
rect 23673 28169 23707 28203
rect 23707 28169 23716 28203
rect 23664 28160 23716 28169
rect 24032 28160 24084 28212
rect 25044 28160 25096 28212
rect 25504 28160 25556 28212
rect 17040 28067 17092 28076
rect 17040 28033 17049 28067
rect 17049 28033 17083 28067
rect 17083 28033 17092 28067
rect 17040 28024 17092 28033
rect 17500 28024 17552 28076
rect 18144 28024 18196 28076
rect 17960 27956 18012 28008
rect 18328 28024 18380 28076
rect 18972 28024 19024 28076
rect 19340 28067 19392 28076
rect 19340 28033 19349 28067
rect 19349 28033 19383 28067
rect 19383 28033 19392 28067
rect 19340 28024 19392 28033
rect 22928 28024 22980 28076
rect 23296 28024 23348 28076
rect 23572 28024 23624 28076
rect 24032 28067 24084 28076
rect 24032 28033 24066 28067
rect 24066 28033 24084 28067
rect 24032 28024 24084 28033
rect 25964 28024 26016 28076
rect 27528 28160 27580 28212
rect 27712 28160 27764 28212
rect 28816 28160 28868 28212
rect 29000 28203 29052 28212
rect 29000 28169 29009 28203
rect 29009 28169 29043 28203
rect 29043 28169 29052 28203
rect 29000 28160 29052 28169
rect 30380 28203 30432 28212
rect 30380 28169 30389 28203
rect 30389 28169 30423 28203
rect 30423 28169 30432 28203
rect 30380 28160 30432 28169
rect 27160 28067 27212 28076
rect 27160 28033 27169 28067
rect 27169 28033 27203 28067
rect 27203 28033 27212 28067
rect 27160 28024 27212 28033
rect 18696 27956 18748 28008
rect 20076 27956 20128 28008
rect 25412 27999 25464 28008
rect 25412 27965 25421 27999
rect 25421 27965 25455 27999
rect 25455 27965 25464 27999
rect 25412 27956 25464 27965
rect 20260 27888 20312 27940
rect 18052 27863 18104 27872
rect 18052 27829 18061 27863
rect 18061 27829 18095 27863
rect 18095 27829 18104 27863
rect 18052 27820 18104 27829
rect 27620 27956 27672 28008
rect 29000 28024 29052 28076
rect 29184 28067 29236 28076
rect 29184 28033 29193 28067
rect 29193 28033 29227 28067
rect 29227 28033 29236 28067
rect 29184 28024 29236 28033
rect 31208 28160 31260 28212
rect 31760 28160 31812 28212
rect 32404 28160 32456 28212
rect 31392 28092 31444 28144
rect 30932 28024 30984 28076
rect 27896 27999 27948 28008
rect 27896 27965 27905 27999
rect 27905 27965 27939 27999
rect 27939 27965 27948 27999
rect 27896 27956 27948 27965
rect 31116 28067 31168 28076
rect 31116 28033 31125 28067
rect 31125 28033 31159 28067
rect 31159 28033 31168 28067
rect 31116 28024 31168 28033
rect 32128 28067 32180 28076
rect 32128 28033 32137 28067
rect 32137 28033 32171 28067
rect 32171 28033 32180 28067
rect 32128 28024 32180 28033
rect 32404 28067 32456 28076
rect 32404 28033 32413 28067
rect 32413 28033 32447 28067
rect 32447 28033 32456 28067
rect 32404 28024 32456 28033
rect 27436 27888 27488 27940
rect 27988 27888 28040 27940
rect 29368 27888 29420 27940
rect 27712 27820 27764 27872
rect 31300 27863 31352 27872
rect 31300 27829 31309 27863
rect 31309 27829 31343 27863
rect 31343 27829 31352 27863
rect 31300 27820 31352 27829
rect 31668 27863 31720 27872
rect 31668 27829 31677 27863
rect 31677 27829 31711 27863
rect 31711 27829 31720 27863
rect 31668 27820 31720 27829
rect 32496 27820 32548 27872
rect 32772 27820 32824 27872
rect 5170 27718 5222 27770
rect 5234 27718 5286 27770
rect 5298 27718 5350 27770
rect 5362 27718 5414 27770
rect 5426 27718 5478 27770
rect 13611 27718 13663 27770
rect 13675 27718 13727 27770
rect 13739 27718 13791 27770
rect 13803 27718 13855 27770
rect 13867 27718 13919 27770
rect 22052 27718 22104 27770
rect 22116 27718 22168 27770
rect 22180 27718 22232 27770
rect 22244 27718 22296 27770
rect 22308 27718 22360 27770
rect 30493 27718 30545 27770
rect 30557 27718 30609 27770
rect 30621 27718 30673 27770
rect 30685 27718 30737 27770
rect 30749 27718 30801 27770
rect 17960 27659 18012 27668
rect 17960 27625 17969 27659
rect 17969 27625 18003 27659
rect 18003 27625 18012 27659
rect 17960 27616 18012 27625
rect 18144 27616 18196 27668
rect 18052 27548 18104 27600
rect 16672 27412 16724 27464
rect 18880 27480 18932 27532
rect 17960 27412 18012 27464
rect 21088 27616 21140 27668
rect 21824 27616 21876 27668
rect 22928 27659 22980 27668
rect 22928 27625 22937 27659
rect 22937 27625 22971 27659
rect 22971 27625 22980 27659
rect 22928 27616 22980 27625
rect 24032 27616 24084 27668
rect 20628 27548 20680 27600
rect 23756 27548 23808 27600
rect 18420 27344 18472 27396
rect 17500 27276 17552 27328
rect 20260 27412 20312 27464
rect 20996 27523 21048 27532
rect 20996 27489 21005 27523
rect 21005 27489 21039 27523
rect 21039 27489 21048 27523
rect 20996 27480 21048 27489
rect 18972 27319 19024 27328
rect 18972 27285 18981 27319
rect 18981 27285 19015 27319
rect 19015 27285 19024 27319
rect 18972 27276 19024 27285
rect 19340 27276 19392 27328
rect 19432 27319 19484 27328
rect 19432 27285 19441 27319
rect 19441 27285 19475 27319
rect 19475 27285 19484 27319
rect 19432 27276 19484 27285
rect 20444 27344 20496 27396
rect 21088 27412 21140 27464
rect 23112 27455 23164 27464
rect 23112 27421 23121 27455
rect 23121 27421 23155 27455
rect 23155 27421 23164 27455
rect 23112 27412 23164 27421
rect 23664 27412 23716 27464
rect 20352 27276 20404 27328
rect 20812 27276 20864 27328
rect 23756 27276 23808 27328
rect 25044 27616 25096 27668
rect 25136 27616 25188 27668
rect 25964 27659 26016 27668
rect 25964 27625 25973 27659
rect 25973 27625 26007 27659
rect 26007 27625 26016 27659
rect 25964 27616 26016 27625
rect 24124 27344 24176 27396
rect 25320 27412 25372 27464
rect 25504 27455 25556 27464
rect 25504 27421 25513 27455
rect 25513 27421 25547 27455
rect 25547 27421 25556 27455
rect 25504 27412 25556 27421
rect 25780 27455 25832 27464
rect 25780 27421 25789 27455
rect 25789 27421 25823 27455
rect 25823 27421 25832 27455
rect 25780 27412 25832 27421
rect 27896 27548 27948 27600
rect 24768 27387 24820 27396
rect 24768 27353 24777 27387
rect 24777 27353 24811 27387
rect 24811 27353 24820 27387
rect 24768 27344 24820 27353
rect 24952 27387 25004 27396
rect 24952 27353 24961 27387
rect 24961 27353 24995 27387
rect 24995 27353 25004 27387
rect 24952 27344 25004 27353
rect 26884 27412 26936 27464
rect 26976 27412 27028 27464
rect 27436 27455 27488 27464
rect 27436 27421 27445 27455
rect 27445 27421 27479 27455
rect 27479 27421 27488 27455
rect 27436 27412 27488 27421
rect 27712 27344 27764 27396
rect 27896 27455 27948 27464
rect 27896 27421 27905 27455
rect 27905 27421 27939 27455
rect 27939 27421 27948 27455
rect 27896 27412 27948 27421
rect 28080 27616 28132 27668
rect 32404 27659 32456 27668
rect 32404 27625 32413 27659
rect 32413 27625 32447 27659
rect 32447 27625 32456 27659
rect 32404 27616 32456 27625
rect 29000 27548 29052 27600
rect 28264 27412 28316 27464
rect 28724 27455 28776 27464
rect 28724 27421 28733 27455
rect 28733 27421 28767 27455
rect 28767 27421 28776 27455
rect 28724 27412 28776 27421
rect 28908 27455 28960 27464
rect 28908 27421 28917 27455
rect 28917 27421 28951 27455
rect 28951 27421 28960 27455
rect 28908 27412 28960 27421
rect 28816 27344 28868 27396
rect 31024 27455 31076 27464
rect 31024 27421 31033 27455
rect 31033 27421 31067 27455
rect 31067 27421 31076 27455
rect 31024 27412 31076 27421
rect 31300 27455 31352 27464
rect 31300 27421 31334 27455
rect 31334 27421 31352 27455
rect 31300 27412 31352 27421
rect 29092 27276 29144 27328
rect 31484 27276 31536 27328
rect 9390 27174 9442 27226
rect 9454 27174 9506 27226
rect 9518 27174 9570 27226
rect 9582 27174 9634 27226
rect 9646 27174 9698 27226
rect 17831 27174 17883 27226
rect 17895 27174 17947 27226
rect 17959 27174 18011 27226
rect 18023 27174 18075 27226
rect 18087 27174 18139 27226
rect 26272 27174 26324 27226
rect 26336 27174 26388 27226
rect 26400 27174 26452 27226
rect 26464 27174 26516 27226
rect 26528 27174 26580 27226
rect 34713 27174 34765 27226
rect 34777 27174 34829 27226
rect 34841 27174 34893 27226
rect 34905 27174 34957 27226
rect 34969 27174 35021 27226
rect 16856 27072 16908 27124
rect 18236 27115 18288 27124
rect 18236 27081 18245 27115
rect 18245 27081 18279 27115
rect 18279 27081 18288 27115
rect 18236 27072 18288 27081
rect 19340 27072 19392 27124
rect 18972 27004 19024 27056
rect 17316 26936 17368 26988
rect 17684 26979 17736 26988
rect 17684 26945 17694 26979
rect 17694 26945 17728 26979
rect 17728 26945 17736 26979
rect 17684 26936 17736 26945
rect 17868 26979 17920 26988
rect 17868 26945 17877 26979
rect 17877 26945 17911 26979
rect 17911 26945 17920 26979
rect 17868 26936 17920 26945
rect 18420 26936 18472 26988
rect 19432 27047 19484 27056
rect 19432 27013 19450 27047
rect 19450 27013 19484 27047
rect 19432 27004 19484 27013
rect 18236 26868 18288 26920
rect 19708 26911 19760 26920
rect 19708 26877 19717 26911
rect 19717 26877 19751 26911
rect 19751 26877 19760 26911
rect 20352 27004 20404 27056
rect 20904 27072 20956 27124
rect 21088 27115 21140 27124
rect 21088 27081 21097 27115
rect 21097 27081 21131 27115
rect 21131 27081 21140 27115
rect 21088 27072 21140 27081
rect 21272 27072 21324 27124
rect 19708 26868 19760 26877
rect 20076 26911 20128 26920
rect 20076 26877 20085 26911
rect 20085 26877 20119 26911
rect 20119 26877 20128 26911
rect 20076 26868 20128 26877
rect 20536 26979 20588 26988
rect 20536 26945 20545 26979
rect 20545 26945 20579 26979
rect 20579 26945 20588 26979
rect 20536 26936 20588 26945
rect 21180 26979 21232 26988
rect 20720 26868 20772 26920
rect 17500 26800 17552 26852
rect 21180 26945 21189 26979
rect 21189 26945 21223 26979
rect 21223 26945 21232 26979
rect 21180 26936 21232 26945
rect 21364 26979 21416 26988
rect 21364 26945 21373 26979
rect 21373 26945 21407 26979
rect 21407 26945 21416 26979
rect 21364 26936 21416 26945
rect 21272 26911 21324 26920
rect 21272 26877 21281 26911
rect 21281 26877 21315 26911
rect 21315 26877 21324 26911
rect 21272 26868 21324 26877
rect 16948 26732 17000 26784
rect 18512 26732 18564 26784
rect 19432 26732 19484 26784
rect 20720 26732 20772 26784
rect 21088 26732 21140 26784
rect 21180 26732 21232 26784
rect 21732 26732 21784 26784
rect 22468 26936 22520 26988
rect 23572 27072 23624 27124
rect 24768 27072 24820 27124
rect 23204 26979 23256 26988
rect 23204 26945 23213 26979
rect 23213 26945 23247 26979
rect 23247 26945 23256 26979
rect 23204 26936 23256 26945
rect 24124 27004 24176 27056
rect 24492 27004 24544 27056
rect 25780 27072 25832 27124
rect 28908 27072 28960 27124
rect 29184 27072 29236 27124
rect 29368 27072 29420 27124
rect 31116 27072 31168 27124
rect 23204 26800 23256 26852
rect 24768 26936 24820 26988
rect 24952 26936 25004 26988
rect 25320 26979 25372 26988
rect 25320 26945 25329 26979
rect 25329 26945 25363 26979
rect 25363 26945 25372 26979
rect 25320 26936 25372 26945
rect 25504 26979 25556 26988
rect 25504 26945 25513 26979
rect 25513 26945 25547 26979
rect 25547 26945 25556 26979
rect 25504 26936 25556 26945
rect 28816 26936 28868 26988
rect 27344 26868 27396 26920
rect 29000 26936 29052 26988
rect 32404 27072 32456 27124
rect 29092 26868 29144 26920
rect 30932 26979 30984 26988
rect 30932 26945 30941 26979
rect 30941 26945 30975 26979
rect 30975 26945 30984 26979
rect 30932 26936 30984 26945
rect 31208 26936 31260 26988
rect 33048 26800 33100 26852
rect 22836 26732 22888 26784
rect 32220 26732 32272 26784
rect 5170 26630 5222 26682
rect 5234 26630 5286 26682
rect 5298 26630 5350 26682
rect 5362 26630 5414 26682
rect 5426 26630 5478 26682
rect 13611 26630 13663 26682
rect 13675 26630 13727 26682
rect 13739 26630 13791 26682
rect 13803 26630 13855 26682
rect 13867 26630 13919 26682
rect 22052 26630 22104 26682
rect 22116 26630 22168 26682
rect 22180 26630 22232 26682
rect 22244 26630 22296 26682
rect 22308 26630 22360 26682
rect 30493 26630 30545 26682
rect 30557 26630 30609 26682
rect 30621 26630 30673 26682
rect 30685 26630 30737 26682
rect 30749 26630 30801 26682
rect 17684 26571 17736 26580
rect 17684 26537 17693 26571
rect 17693 26537 17727 26571
rect 17727 26537 17736 26571
rect 17684 26528 17736 26537
rect 17868 26528 17920 26580
rect 18512 26528 18564 26580
rect 19708 26528 19760 26580
rect 20076 26528 20128 26580
rect 20904 26571 20956 26580
rect 20904 26537 20913 26571
rect 20913 26537 20947 26571
rect 20947 26537 20956 26571
rect 20904 26528 20956 26537
rect 22468 26528 22520 26580
rect 18880 26460 18932 26512
rect 20812 26460 20864 26512
rect 21088 26460 21140 26512
rect 20720 26435 20772 26444
rect 20720 26401 20729 26435
rect 20729 26401 20763 26435
rect 20763 26401 20772 26435
rect 20720 26392 20772 26401
rect 21916 26460 21968 26512
rect 23756 26528 23808 26580
rect 24584 26571 24636 26580
rect 24584 26537 24593 26571
rect 24593 26537 24627 26571
rect 24627 26537 24636 26571
rect 24584 26528 24636 26537
rect 25320 26528 25372 26580
rect 25504 26528 25556 26580
rect 26976 26528 27028 26580
rect 27436 26528 27488 26580
rect 29092 26528 29144 26580
rect 16856 26324 16908 26376
rect 17592 26324 17644 26376
rect 19432 26367 19484 26376
rect 19432 26333 19441 26367
rect 19441 26333 19475 26367
rect 19475 26333 19484 26367
rect 19432 26324 19484 26333
rect 20536 26324 20588 26376
rect 20904 26324 20956 26376
rect 21272 26367 21324 26376
rect 21272 26333 21281 26367
rect 21281 26333 21315 26367
rect 21315 26333 21324 26367
rect 21272 26324 21324 26333
rect 21364 26367 21416 26376
rect 21364 26333 21373 26367
rect 21373 26333 21407 26367
rect 21407 26333 21416 26367
rect 21364 26324 21416 26333
rect 16672 26256 16724 26308
rect 18512 26256 18564 26308
rect 20260 26299 20312 26308
rect 20260 26265 20269 26299
rect 20269 26265 20303 26299
rect 20303 26265 20312 26299
rect 20260 26256 20312 26265
rect 21732 26367 21784 26376
rect 21732 26333 21741 26367
rect 21741 26333 21775 26367
rect 21775 26333 21784 26367
rect 21732 26324 21784 26333
rect 21824 26256 21876 26308
rect 22468 26299 22520 26308
rect 22468 26265 22477 26299
rect 22477 26265 22511 26299
rect 22511 26265 22520 26299
rect 22468 26256 22520 26265
rect 22836 26367 22888 26376
rect 22836 26333 22845 26367
rect 22845 26333 22879 26367
rect 22879 26333 22888 26367
rect 22836 26324 22888 26333
rect 23480 26256 23532 26308
rect 24768 26299 24820 26308
rect 24768 26265 24777 26299
rect 24777 26265 24811 26299
rect 24811 26265 24820 26299
rect 24768 26256 24820 26265
rect 17408 26188 17460 26240
rect 21272 26188 21324 26240
rect 23572 26188 23624 26240
rect 24216 26231 24268 26240
rect 24216 26197 24225 26231
rect 24225 26197 24259 26231
rect 24259 26197 24268 26231
rect 24216 26188 24268 26197
rect 24952 26231 25004 26240
rect 24952 26197 24961 26231
rect 24961 26197 24995 26231
rect 24995 26197 25004 26231
rect 24952 26188 25004 26197
rect 26148 26324 26200 26376
rect 26240 26367 26292 26376
rect 26240 26333 26249 26367
rect 26249 26333 26283 26367
rect 26283 26333 26292 26367
rect 26240 26324 26292 26333
rect 26884 26460 26936 26512
rect 28724 26460 28776 26512
rect 29552 26460 29604 26512
rect 32956 26460 33008 26512
rect 27252 26392 27304 26444
rect 27804 26392 27856 26444
rect 27344 26367 27396 26376
rect 27344 26333 27353 26367
rect 27353 26333 27387 26367
rect 27387 26333 27396 26367
rect 27344 26324 27396 26333
rect 27436 26367 27488 26376
rect 27436 26333 27445 26367
rect 27445 26333 27479 26367
rect 27479 26333 27488 26367
rect 27436 26324 27488 26333
rect 28632 26324 28684 26376
rect 28816 26367 28868 26376
rect 28816 26333 28825 26367
rect 28825 26333 28859 26367
rect 28859 26333 28868 26367
rect 28816 26324 28868 26333
rect 30840 26392 30892 26444
rect 29828 26324 29880 26376
rect 31024 26324 31076 26376
rect 31760 26324 31812 26376
rect 32220 26367 32272 26376
rect 32220 26333 32254 26367
rect 32254 26333 32272 26367
rect 32220 26324 32272 26333
rect 28908 26256 28960 26308
rect 25688 26188 25740 26240
rect 26240 26188 26292 26240
rect 26700 26188 26752 26240
rect 27712 26188 27764 26240
rect 27804 26231 27856 26240
rect 27804 26197 27813 26231
rect 27813 26197 27847 26231
rect 27847 26197 27856 26231
rect 27804 26188 27856 26197
rect 30012 26231 30064 26240
rect 30012 26197 30021 26231
rect 30021 26197 30055 26231
rect 30055 26197 30064 26231
rect 30012 26188 30064 26197
rect 9390 26086 9442 26138
rect 9454 26086 9506 26138
rect 9518 26086 9570 26138
rect 9582 26086 9634 26138
rect 9646 26086 9698 26138
rect 17831 26086 17883 26138
rect 17895 26086 17947 26138
rect 17959 26086 18011 26138
rect 18023 26086 18075 26138
rect 18087 26086 18139 26138
rect 26272 26086 26324 26138
rect 26336 26086 26388 26138
rect 26400 26086 26452 26138
rect 26464 26086 26516 26138
rect 26528 26086 26580 26138
rect 34713 26086 34765 26138
rect 34777 26086 34829 26138
rect 34841 26086 34893 26138
rect 34905 26086 34957 26138
rect 34969 26086 35021 26138
rect 17500 26027 17552 26036
rect 17500 25993 17509 26027
rect 17509 25993 17543 26027
rect 17543 25993 17552 26027
rect 17500 25984 17552 25993
rect 17776 25916 17828 25968
rect 17132 25891 17184 25900
rect 17132 25857 17141 25891
rect 17141 25857 17175 25891
rect 17175 25857 17184 25891
rect 17132 25848 17184 25857
rect 17316 25780 17368 25832
rect 17960 25848 18012 25900
rect 20904 25984 20956 26036
rect 19156 25891 19208 25900
rect 19156 25857 19165 25891
rect 19165 25857 19199 25891
rect 19199 25857 19208 25891
rect 19156 25848 19208 25857
rect 21180 25916 21232 25968
rect 24584 25984 24636 26036
rect 19984 25848 20036 25900
rect 21456 25891 21508 25900
rect 21456 25857 21465 25891
rect 21465 25857 21499 25891
rect 21499 25857 21508 25891
rect 21456 25848 21508 25857
rect 22744 25848 22796 25900
rect 22836 25848 22888 25900
rect 23572 25848 23624 25900
rect 24216 25916 24268 25968
rect 24308 25916 24360 25968
rect 25044 25916 25096 25968
rect 26700 26027 26752 26036
rect 26700 25993 26709 26027
rect 26709 25993 26743 26027
rect 26743 25993 26752 26027
rect 26700 25984 26752 25993
rect 27344 25984 27396 26036
rect 27620 26027 27672 26036
rect 27620 25993 27629 26027
rect 27629 25993 27663 26027
rect 27663 25993 27672 26027
rect 27620 25984 27672 25993
rect 26148 25959 26200 25968
rect 26148 25925 26157 25959
rect 26157 25925 26191 25959
rect 26191 25925 26200 25959
rect 26148 25916 26200 25925
rect 24676 25848 24728 25900
rect 25412 25848 25464 25900
rect 17224 25644 17276 25696
rect 18420 25712 18472 25764
rect 19156 25712 19208 25764
rect 19892 25780 19944 25832
rect 20996 25780 21048 25832
rect 21548 25780 21600 25832
rect 23480 25780 23532 25832
rect 18328 25644 18380 25696
rect 18696 25687 18748 25696
rect 18696 25653 18705 25687
rect 18705 25653 18739 25687
rect 18739 25653 18748 25687
rect 18696 25644 18748 25653
rect 19800 25644 19852 25696
rect 23572 25687 23624 25696
rect 23572 25653 23581 25687
rect 23581 25653 23615 25687
rect 23615 25653 23624 25687
rect 23572 25644 23624 25653
rect 24860 25644 24912 25696
rect 25688 25891 25740 25900
rect 25688 25857 25697 25891
rect 25697 25857 25731 25891
rect 25731 25857 25740 25891
rect 25688 25848 25740 25857
rect 25872 25687 25924 25696
rect 25872 25653 25881 25687
rect 25881 25653 25915 25687
rect 25915 25653 25924 25687
rect 25872 25644 25924 25653
rect 26056 25644 26108 25696
rect 26700 25848 26752 25900
rect 28816 25984 28868 26036
rect 29552 25984 29604 26036
rect 27896 25891 27948 25900
rect 27896 25857 27905 25891
rect 27905 25857 27939 25891
rect 27939 25857 27948 25891
rect 27896 25848 27948 25857
rect 28632 25891 28684 25900
rect 28632 25857 28641 25891
rect 28641 25857 28675 25891
rect 28675 25857 28684 25891
rect 28632 25848 28684 25857
rect 27436 25780 27488 25832
rect 27712 25780 27764 25832
rect 28908 25780 28960 25832
rect 27252 25644 27304 25696
rect 29368 25644 29420 25696
rect 29736 25780 29788 25832
rect 30012 25848 30064 25900
rect 30104 25848 30156 25900
rect 31208 25984 31260 26036
rect 32588 26027 32640 26036
rect 32588 25993 32597 26027
rect 32597 25993 32631 26027
rect 32631 25993 32640 26027
rect 32588 25984 32640 25993
rect 31484 25891 31536 25900
rect 31484 25857 31493 25891
rect 31493 25857 31527 25891
rect 31527 25857 31536 25891
rect 31484 25848 31536 25857
rect 32956 25848 33008 25900
rect 32312 25823 32364 25832
rect 32312 25789 32321 25823
rect 32321 25789 32355 25823
rect 32355 25789 32364 25823
rect 32312 25780 32364 25789
rect 32680 25823 32732 25832
rect 32680 25789 32689 25823
rect 32689 25789 32723 25823
rect 32723 25789 32732 25823
rect 32680 25780 32732 25789
rect 32772 25823 32824 25832
rect 32772 25789 32781 25823
rect 32781 25789 32815 25823
rect 32815 25789 32824 25823
rect 32772 25780 32824 25789
rect 30380 25712 30432 25764
rect 29920 25644 29972 25696
rect 30104 25644 30156 25696
rect 30840 25644 30892 25696
rect 31576 25644 31628 25696
rect 31760 25644 31812 25696
rect 32128 25687 32180 25696
rect 32128 25653 32137 25687
rect 32137 25653 32171 25687
rect 32171 25653 32180 25687
rect 32128 25644 32180 25653
rect 5170 25542 5222 25594
rect 5234 25542 5286 25594
rect 5298 25542 5350 25594
rect 5362 25542 5414 25594
rect 5426 25542 5478 25594
rect 13611 25542 13663 25594
rect 13675 25542 13727 25594
rect 13739 25542 13791 25594
rect 13803 25542 13855 25594
rect 13867 25542 13919 25594
rect 22052 25542 22104 25594
rect 22116 25542 22168 25594
rect 22180 25542 22232 25594
rect 22244 25542 22296 25594
rect 22308 25542 22360 25594
rect 30493 25542 30545 25594
rect 30557 25542 30609 25594
rect 30621 25542 30673 25594
rect 30685 25542 30737 25594
rect 30749 25542 30801 25594
rect 17132 25440 17184 25492
rect 18236 25440 18288 25492
rect 18328 25440 18380 25492
rect 18696 25440 18748 25492
rect 19800 25483 19852 25492
rect 19800 25449 19809 25483
rect 19809 25449 19843 25483
rect 19843 25449 19852 25483
rect 19800 25440 19852 25449
rect 19892 25440 19944 25492
rect 19984 25440 20036 25492
rect 17316 25372 17368 25424
rect 16948 25236 17000 25288
rect 19340 25415 19392 25424
rect 19340 25381 19349 25415
rect 19349 25381 19383 25415
rect 19383 25381 19392 25415
rect 19340 25372 19392 25381
rect 19524 25279 19576 25288
rect 19524 25245 19533 25279
rect 19533 25245 19567 25279
rect 19567 25245 19576 25279
rect 19524 25236 19576 25245
rect 22744 25440 22796 25492
rect 24676 25483 24728 25492
rect 24676 25449 24685 25483
rect 24685 25449 24719 25483
rect 24719 25449 24728 25483
rect 24676 25440 24728 25449
rect 20904 25372 20956 25424
rect 20996 25372 21048 25424
rect 21272 25372 21324 25424
rect 20260 25304 20312 25356
rect 20260 25168 20312 25220
rect 20444 25236 20496 25288
rect 20996 25168 21048 25220
rect 21824 25236 21876 25288
rect 22468 25236 22520 25288
rect 23940 25304 23992 25356
rect 21456 25168 21508 25220
rect 22744 25168 22796 25220
rect 23572 25168 23624 25220
rect 25872 25440 25924 25492
rect 26700 25440 26752 25492
rect 27896 25440 27948 25492
rect 28632 25440 28684 25492
rect 29368 25483 29420 25492
rect 29368 25449 29377 25483
rect 29377 25449 29411 25483
rect 29411 25449 29420 25483
rect 29368 25440 29420 25449
rect 29736 25440 29788 25492
rect 30104 25440 30156 25492
rect 32312 25440 32364 25492
rect 24952 25372 25004 25424
rect 25688 25372 25740 25424
rect 29828 25415 29880 25424
rect 29828 25381 29837 25415
rect 29837 25381 29871 25415
rect 29871 25381 29880 25415
rect 29828 25372 29880 25381
rect 28908 25304 28960 25356
rect 25412 25236 25464 25288
rect 25504 25168 25556 25220
rect 25964 25211 26016 25220
rect 25964 25177 25998 25211
rect 25998 25177 26016 25211
rect 25964 25168 26016 25177
rect 27804 25236 27856 25288
rect 29184 25279 29236 25288
rect 29184 25245 29193 25279
rect 29193 25245 29227 25279
rect 29227 25245 29236 25279
rect 29184 25236 29236 25245
rect 29368 25279 29420 25288
rect 29368 25245 29389 25279
rect 29389 25245 29420 25279
rect 29368 25236 29420 25245
rect 30104 25236 30156 25288
rect 29092 25168 29144 25220
rect 29552 25211 29604 25220
rect 29552 25177 29561 25211
rect 29561 25177 29595 25211
rect 29595 25177 29604 25211
rect 29552 25168 29604 25177
rect 30840 25236 30892 25288
rect 31576 25236 31628 25288
rect 31760 25168 31812 25220
rect 16948 25143 17000 25152
rect 16948 25109 16957 25143
rect 16957 25109 16991 25143
rect 16991 25109 17000 25143
rect 16948 25100 17000 25109
rect 17224 25100 17276 25152
rect 18236 25100 18288 25152
rect 20352 25100 20404 25152
rect 20720 25143 20772 25152
rect 20720 25109 20729 25143
rect 20729 25109 20763 25143
rect 20763 25109 20772 25143
rect 20720 25100 20772 25109
rect 21272 25100 21324 25152
rect 23756 25100 23808 25152
rect 31576 25143 31628 25152
rect 31576 25109 31585 25143
rect 31585 25109 31619 25143
rect 31619 25109 31628 25143
rect 31576 25100 31628 25109
rect 9390 24998 9442 25050
rect 9454 24998 9506 25050
rect 9518 24998 9570 25050
rect 9582 24998 9634 25050
rect 9646 24998 9698 25050
rect 17831 24998 17883 25050
rect 17895 24998 17947 25050
rect 17959 24998 18011 25050
rect 18023 24998 18075 25050
rect 18087 24998 18139 25050
rect 26272 24998 26324 25050
rect 26336 24998 26388 25050
rect 26400 24998 26452 25050
rect 26464 24998 26516 25050
rect 26528 24998 26580 25050
rect 34713 24998 34765 25050
rect 34777 24998 34829 25050
rect 34841 24998 34893 25050
rect 34905 24998 34957 25050
rect 34969 24998 35021 25050
rect 17132 24896 17184 24948
rect 16948 24871 17000 24880
rect 16948 24837 16982 24871
rect 16982 24837 17000 24871
rect 16948 24828 17000 24837
rect 18236 24896 18288 24948
rect 18420 24896 18472 24948
rect 19524 24896 19576 24948
rect 20444 24896 20496 24948
rect 20536 24939 20588 24948
rect 20536 24905 20545 24939
rect 20545 24905 20579 24939
rect 20579 24905 20588 24939
rect 20536 24896 20588 24905
rect 19248 24760 19300 24812
rect 21916 24896 21968 24948
rect 23756 24896 23808 24948
rect 25044 24939 25096 24948
rect 25044 24905 25053 24939
rect 25053 24905 25087 24939
rect 25087 24905 25096 24939
rect 25044 24896 25096 24905
rect 25964 24896 26016 24948
rect 18236 24692 18288 24744
rect 18512 24735 18564 24744
rect 18512 24701 18521 24735
rect 18521 24701 18555 24735
rect 18555 24701 18564 24735
rect 18512 24692 18564 24701
rect 20720 24692 20772 24744
rect 16948 24556 17000 24608
rect 20352 24624 20404 24676
rect 21548 24760 21600 24812
rect 22560 24760 22612 24812
rect 24952 24803 25004 24812
rect 24952 24769 24961 24803
rect 24961 24769 24995 24803
rect 24995 24769 25004 24803
rect 24952 24760 25004 24769
rect 26056 24803 26108 24812
rect 26056 24769 26065 24803
rect 26065 24769 26099 24803
rect 26099 24769 26108 24803
rect 26056 24760 26108 24769
rect 26700 24760 26752 24812
rect 27436 24760 27488 24812
rect 26148 24624 26200 24676
rect 29184 24896 29236 24948
rect 28908 24803 28960 24812
rect 28908 24769 28942 24803
rect 28942 24769 28960 24803
rect 28908 24760 28960 24769
rect 29552 24828 29604 24880
rect 30380 24896 30432 24948
rect 31760 24939 31812 24948
rect 31760 24905 31769 24939
rect 31769 24905 31803 24939
rect 31803 24905 31812 24939
rect 31760 24896 31812 24905
rect 29736 24692 29788 24744
rect 30840 24803 30892 24812
rect 30840 24769 30849 24803
rect 30849 24769 30883 24803
rect 30883 24769 30892 24803
rect 30840 24760 30892 24769
rect 30932 24692 30984 24744
rect 31116 24803 31168 24812
rect 31116 24769 31125 24803
rect 31125 24769 31159 24803
rect 31159 24769 31168 24803
rect 31116 24760 31168 24769
rect 31208 24760 31260 24812
rect 21088 24599 21140 24608
rect 21088 24565 21097 24599
rect 21097 24565 21131 24599
rect 21131 24565 21140 24599
rect 21088 24556 21140 24565
rect 21272 24599 21324 24608
rect 21272 24565 21281 24599
rect 21281 24565 21315 24599
rect 21315 24565 21324 24599
rect 21272 24556 21324 24565
rect 22652 24599 22704 24608
rect 22652 24565 22661 24599
rect 22661 24565 22695 24599
rect 22695 24565 22704 24599
rect 22652 24556 22704 24565
rect 23112 24556 23164 24608
rect 23204 24556 23256 24608
rect 24308 24599 24360 24608
rect 24308 24565 24317 24599
rect 24317 24565 24351 24599
rect 24351 24565 24360 24599
rect 24308 24556 24360 24565
rect 25136 24556 25188 24608
rect 28540 24599 28592 24608
rect 28540 24565 28549 24599
rect 28549 24565 28583 24599
rect 28583 24565 28592 24599
rect 28540 24556 28592 24565
rect 31208 24624 31260 24676
rect 31576 24760 31628 24812
rect 32312 24760 32364 24812
rect 32496 24803 32548 24812
rect 32496 24769 32505 24803
rect 32505 24769 32539 24803
rect 32539 24769 32548 24803
rect 32496 24760 32548 24769
rect 32220 24692 32272 24744
rect 32680 24760 32732 24812
rect 32864 24803 32916 24812
rect 32864 24769 32873 24803
rect 32873 24769 32907 24803
rect 32907 24769 32916 24803
rect 32864 24760 32916 24769
rect 33048 24760 33100 24812
rect 32128 24624 32180 24676
rect 29552 24556 29604 24608
rect 31024 24599 31076 24608
rect 31024 24565 31033 24599
rect 31033 24565 31067 24599
rect 31067 24565 31076 24599
rect 31024 24556 31076 24565
rect 31484 24556 31536 24608
rect 32680 24599 32732 24608
rect 32680 24565 32689 24599
rect 32689 24565 32723 24599
rect 32723 24565 32732 24599
rect 32680 24556 32732 24565
rect 33324 24556 33376 24608
rect 5170 24454 5222 24506
rect 5234 24454 5286 24506
rect 5298 24454 5350 24506
rect 5362 24454 5414 24506
rect 5426 24454 5478 24506
rect 13611 24454 13663 24506
rect 13675 24454 13727 24506
rect 13739 24454 13791 24506
rect 13803 24454 13855 24506
rect 13867 24454 13919 24506
rect 22052 24454 22104 24506
rect 22116 24454 22168 24506
rect 22180 24454 22232 24506
rect 22244 24454 22296 24506
rect 22308 24454 22360 24506
rect 30493 24454 30545 24506
rect 30557 24454 30609 24506
rect 30621 24454 30673 24506
rect 30685 24454 30737 24506
rect 30749 24454 30801 24506
rect 18420 24395 18472 24404
rect 18420 24361 18429 24395
rect 18429 24361 18463 24395
rect 18463 24361 18472 24395
rect 18420 24352 18472 24361
rect 19248 24395 19300 24404
rect 19248 24361 19257 24395
rect 19257 24361 19291 24395
rect 19291 24361 19300 24395
rect 19248 24352 19300 24361
rect 21088 24352 21140 24404
rect 21548 24352 21600 24404
rect 22560 24352 22612 24404
rect 22744 24352 22796 24404
rect 23112 24352 23164 24404
rect 24308 24352 24360 24404
rect 28540 24352 28592 24404
rect 28908 24352 28960 24404
rect 30840 24352 30892 24404
rect 31024 24352 31076 24404
rect 31208 24352 31260 24404
rect 33324 24395 33376 24404
rect 33324 24361 33333 24395
rect 33333 24361 33367 24395
rect 33367 24361 33376 24395
rect 33324 24352 33376 24361
rect 16948 24216 17000 24268
rect 18236 24216 18288 24268
rect 18880 24216 18932 24268
rect 19524 24216 19576 24268
rect 21916 24284 21968 24336
rect 17316 24191 17368 24200
rect 17316 24157 17350 24191
rect 17350 24157 17368 24191
rect 17316 24148 17368 24157
rect 19340 24148 19392 24200
rect 20168 24055 20220 24064
rect 20168 24021 20177 24055
rect 20177 24021 20211 24055
rect 20211 24021 20220 24055
rect 20168 24012 20220 24021
rect 20720 24148 20772 24200
rect 20904 24191 20956 24200
rect 20904 24157 20913 24191
rect 20913 24157 20947 24191
rect 20947 24157 20956 24191
rect 20904 24148 20956 24157
rect 22652 24284 22704 24336
rect 20996 24012 21048 24064
rect 21456 24012 21508 24064
rect 22928 24191 22980 24200
rect 22928 24157 22937 24191
rect 22937 24157 22971 24191
rect 22971 24157 22980 24191
rect 22928 24148 22980 24157
rect 22744 24012 22796 24064
rect 23112 24012 23164 24064
rect 23572 24191 23624 24200
rect 23572 24157 23581 24191
rect 23581 24157 23615 24191
rect 23615 24157 23624 24191
rect 23572 24148 23624 24157
rect 23848 24191 23900 24200
rect 23848 24157 23857 24191
rect 23857 24157 23891 24191
rect 23891 24157 23900 24191
rect 23848 24148 23900 24157
rect 24676 24191 24728 24200
rect 24676 24157 24685 24191
rect 24685 24157 24719 24191
rect 24719 24157 24728 24191
rect 24676 24148 24728 24157
rect 29552 24080 29604 24132
rect 32036 24080 32088 24132
rect 32588 24080 32640 24132
rect 24124 24055 24176 24064
rect 24124 24021 24133 24055
rect 24133 24021 24167 24055
rect 24167 24021 24176 24055
rect 24124 24012 24176 24021
rect 25412 24012 25464 24064
rect 26056 24055 26108 24064
rect 26056 24021 26065 24055
rect 26065 24021 26099 24055
rect 26099 24021 26108 24055
rect 26056 24012 26108 24021
rect 31024 24055 31076 24064
rect 31024 24021 31033 24055
rect 31033 24021 31067 24055
rect 31067 24021 31076 24055
rect 31024 24012 31076 24021
rect 31300 24055 31352 24064
rect 31300 24021 31309 24055
rect 31309 24021 31343 24055
rect 31343 24021 31352 24055
rect 31300 24012 31352 24021
rect 9390 23910 9442 23962
rect 9454 23910 9506 23962
rect 9518 23910 9570 23962
rect 9582 23910 9634 23962
rect 9646 23910 9698 23962
rect 17831 23910 17883 23962
rect 17895 23910 17947 23962
rect 17959 23910 18011 23962
rect 18023 23910 18075 23962
rect 18087 23910 18139 23962
rect 26272 23910 26324 23962
rect 26336 23910 26388 23962
rect 26400 23910 26452 23962
rect 26464 23910 26516 23962
rect 26528 23910 26580 23962
rect 34713 23910 34765 23962
rect 34777 23910 34829 23962
rect 34841 23910 34893 23962
rect 34905 23910 34957 23962
rect 34969 23910 35021 23962
rect 20168 23808 20220 23860
rect 21456 23851 21508 23860
rect 21456 23817 21465 23851
rect 21465 23817 21499 23851
rect 21499 23817 21508 23851
rect 21456 23808 21508 23817
rect 22744 23808 22796 23860
rect 23204 23851 23256 23860
rect 23204 23817 23213 23851
rect 23213 23817 23247 23851
rect 23247 23817 23256 23851
rect 23204 23808 23256 23817
rect 22928 23740 22980 23792
rect 23572 23808 23624 23860
rect 25136 23851 25188 23860
rect 25136 23817 25145 23851
rect 25145 23817 25179 23851
rect 25179 23817 25188 23851
rect 25136 23808 25188 23817
rect 25596 23808 25648 23860
rect 22376 23672 22428 23724
rect 25412 23740 25464 23792
rect 26148 23783 26200 23792
rect 26148 23749 26157 23783
rect 26157 23749 26191 23783
rect 26191 23749 26200 23783
rect 26148 23740 26200 23749
rect 29828 23808 29880 23860
rect 24400 23672 24452 23724
rect 24492 23672 24544 23724
rect 26516 23715 26568 23724
rect 26516 23681 26525 23715
rect 26525 23681 26559 23715
rect 26559 23681 26568 23715
rect 26516 23672 26568 23681
rect 26792 23672 26844 23724
rect 23664 23647 23716 23656
rect 23664 23613 23673 23647
rect 23673 23613 23707 23647
rect 23707 23613 23716 23647
rect 23664 23604 23716 23613
rect 23388 23536 23440 23588
rect 24860 23604 24912 23656
rect 25872 23604 25924 23656
rect 29276 23672 29328 23724
rect 29644 23715 29696 23724
rect 29644 23681 29653 23715
rect 29653 23681 29687 23715
rect 29687 23681 29696 23715
rect 29644 23672 29696 23681
rect 30196 23672 30248 23724
rect 31024 23808 31076 23860
rect 31300 23808 31352 23860
rect 32588 23851 32640 23860
rect 32588 23817 32597 23851
rect 32597 23817 32631 23851
rect 32631 23817 32640 23851
rect 32588 23808 32640 23817
rect 31944 23672 31996 23724
rect 32220 23604 32272 23656
rect 22928 23468 22980 23520
rect 23296 23511 23348 23520
rect 23296 23477 23305 23511
rect 23305 23477 23339 23511
rect 23339 23477 23348 23511
rect 23296 23468 23348 23477
rect 26332 23511 26384 23520
rect 26332 23477 26341 23511
rect 26341 23477 26375 23511
rect 26375 23477 26384 23511
rect 26332 23468 26384 23477
rect 27896 23468 27948 23520
rect 29920 23511 29972 23520
rect 29920 23477 29929 23511
rect 29929 23477 29963 23511
rect 29963 23477 29972 23511
rect 29920 23468 29972 23477
rect 5170 23366 5222 23418
rect 5234 23366 5286 23418
rect 5298 23366 5350 23418
rect 5362 23366 5414 23418
rect 5426 23366 5478 23418
rect 13611 23366 13663 23418
rect 13675 23366 13727 23418
rect 13739 23366 13791 23418
rect 13803 23366 13855 23418
rect 13867 23366 13919 23418
rect 22052 23366 22104 23418
rect 22116 23366 22168 23418
rect 22180 23366 22232 23418
rect 22244 23366 22296 23418
rect 22308 23366 22360 23418
rect 30493 23366 30545 23418
rect 30557 23366 30609 23418
rect 30621 23366 30673 23418
rect 30685 23366 30737 23418
rect 30749 23366 30801 23418
rect 22376 23264 22428 23316
rect 23112 23264 23164 23316
rect 23572 23307 23624 23316
rect 23572 23273 23581 23307
rect 23581 23273 23615 23307
rect 23615 23273 23624 23307
rect 23572 23264 23624 23273
rect 24400 23307 24452 23316
rect 24400 23273 24409 23307
rect 24409 23273 24443 23307
rect 24443 23273 24452 23307
rect 24400 23264 24452 23273
rect 25504 23307 25556 23316
rect 25504 23273 25513 23307
rect 25513 23273 25547 23307
rect 25547 23273 25556 23307
rect 25504 23264 25556 23273
rect 26056 23264 26108 23316
rect 23756 23239 23808 23248
rect 23756 23205 23765 23239
rect 23765 23205 23799 23239
rect 23799 23205 23808 23239
rect 23756 23196 23808 23205
rect 23848 23128 23900 23180
rect 30196 23264 30248 23316
rect 30932 23307 30984 23316
rect 30932 23273 30941 23307
rect 30941 23273 30975 23307
rect 30975 23273 30984 23307
rect 30932 23264 30984 23273
rect 17040 23060 17092 23112
rect 18328 23060 18380 23112
rect 20628 23103 20680 23112
rect 20628 23069 20637 23103
rect 20637 23069 20671 23103
rect 20671 23069 20680 23103
rect 20628 23060 20680 23069
rect 20720 23060 20772 23112
rect 20904 23060 20956 23112
rect 21732 23103 21784 23112
rect 21732 23069 21741 23103
rect 21741 23069 21775 23103
rect 21775 23069 21784 23103
rect 21732 23060 21784 23069
rect 23296 23060 23348 23112
rect 23756 23060 23808 23112
rect 19800 22992 19852 23044
rect 22376 22992 22428 23044
rect 24124 23060 24176 23112
rect 25412 23103 25464 23112
rect 25412 23069 25421 23103
rect 25421 23069 25455 23103
rect 25455 23069 25464 23103
rect 25412 23060 25464 23069
rect 25872 23103 25924 23112
rect 25872 23069 25881 23103
rect 25881 23069 25915 23103
rect 25915 23069 25924 23103
rect 25872 23060 25924 23069
rect 24860 22992 24912 23044
rect 26332 22992 26384 23044
rect 27896 23060 27948 23112
rect 29276 23171 29328 23180
rect 29276 23137 29285 23171
rect 29285 23137 29319 23171
rect 29319 23137 29328 23171
rect 29276 23128 29328 23137
rect 30380 23060 30432 23112
rect 31208 23103 31260 23112
rect 31208 23069 31217 23103
rect 31217 23069 31251 23103
rect 31251 23069 31260 23103
rect 31208 23060 31260 23069
rect 17408 22967 17460 22976
rect 17408 22933 17417 22967
rect 17417 22933 17451 22967
rect 17451 22933 17460 22967
rect 17408 22924 17460 22933
rect 19064 22924 19116 22976
rect 19984 22924 20036 22976
rect 21824 22967 21876 22976
rect 21824 22933 21833 22967
rect 21833 22933 21867 22967
rect 21867 22933 21876 22967
rect 21824 22924 21876 22933
rect 27252 22967 27304 22976
rect 27252 22933 27261 22967
rect 27261 22933 27295 22967
rect 27295 22933 27304 22967
rect 27252 22924 27304 22933
rect 27344 22967 27396 22976
rect 27344 22933 27353 22967
rect 27353 22933 27387 22967
rect 27387 22933 27396 22967
rect 27344 22924 27396 22933
rect 29000 23035 29052 23044
rect 29000 23001 29018 23035
rect 29018 23001 29052 23035
rect 29000 22992 29052 23001
rect 29184 22992 29236 23044
rect 29920 22992 29972 23044
rect 27988 22924 28040 22976
rect 31024 22967 31076 22976
rect 31024 22933 31033 22967
rect 31033 22933 31067 22967
rect 31067 22933 31076 22967
rect 31024 22924 31076 22933
rect 9390 22822 9442 22874
rect 9454 22822 9506 22874
rect 9518 22822 9570 22874
rect 9582 22822 9634 22874
rect 9646 22822 9698 22874
rect 17831 22822 17883 22874
rect 17895 22822 17947 22874
rect 17959 22822 18011 22874
rect 18023 22822 18075 22874
rect 18087 22822 18139 22874
rect 26272 22822 26324 22874
rect 26336 22822 26388 22874
rect 26400 22822 26452 22874
rect 26464 22822 26516 22874
rect 26528 22822 26580 22874
rect 34713 22822 34765 22874
rect 34777 22822 34829 22874
rect 34841 22822 34893 22874
rect 34905 22822 34957 22874
rect 34969 22822 35021 22874
rect 17408 22720 17460 22772
rect 18328 22763 18380 22772
rect 18328 22729 18337 22763
rect 18337 22729 18371 22763
rect 18371 22729 18380 22763
rect 18328 22720 18380 22729
rect 19800 22720 19852 22772
rect 21732 22720 21784 22772
rect 23020 22720 23072 22772
rect 16948 22559 17000 22568
rect 16948 22525 16957 22559
rect 16957 22525 16991 22559
rect 16991 22525 17000 22559
rect 16948 22516 17000 22525
rect 18788 22584 18840 22636
rect 19064 22627 19116 22636
rect 19064 22593 19073 22627
rect 19073 22593 19107 22627
rect 19107 22593 19116 22627
rect 19064 22584 19116 22593
rect 21364 22627 21416 22636
rect 21364 22593 21373 22627
rect 21373 22593 21407 22627
rect 21407 22593 21416 22627
rect 21364 22584 21416 22593
rect 22100 22627 22152 22636
rect 22100 22593 22109 22627
rect 22109 22593 22143 22627
rect 22143 22593 22152 22627
rect 22100 22584 22152 22593
rect 22376 22652 22428 22704
rect 23388 22763 23440 22772
rect 23388 22729 23397 22763
rect 23397 22729 23431 22763
rect 23431 22729 23440 22763
rect 23388 22720 23440 22729
rect 24952 22720 25004 22772
rect 25412 22720 25464 22772
rect 26148 22720 26200 22772
rect 26608 22720 26660 22772
rect 27988 22720 28040 22772
rect 18880 22559 18932 22568
rect 18880 22525 18889 22559
rect 18889 22525 18923 22559
rect 18923 22525 18932 22559
rect 18880 22516 18932 22525
rect 18604 22448 18656 22500
rect 22928 22584 22980 22636
rect 23388 22584 23440 22636
rect 23664 22516 23716 22568
rect 25412 22584 25464 22636
rect 26056 22584 26108 22636
rect 26700 22584 26752 22636
rect 27896 22627 27948 22636
rect 27896 22593 27905 22627
rect 27905 22593 27939 22627
rect 27939 22593 27948 22627
rect 27896 22584 27948 22593
rect 29000 22763 29052 22772
rect 29000 22729 29009 22763
rect 29009 22729 29043 22763
rect 29043 22729 29052 22763
rect 29000 22720 29052 22729
rect 31024 22720 31076 22772
rect 32036 22720 32088 22772
rect 29552 22695 29604 22704
rect 29552 22661 29561 22695
rect 29561 22661 29595 22695
rect 29595 22661 29604 22695
rect 29552 22652 29604 22661
rect 32864 22695 32916 22704
rect 32864 22661 32873 22695
rect 32873 22661 32907 22695
rect 32907 22661 32916 22695
rect 32864 22652 32916 22661
rect 24768 22559 24820 22568
rect 24768 22525 24777 22559
rect 24777 22525 24811 22559
rect 24811 22525 24820 22559
rect 24768 22516 24820 22525
rect 26240 22516 26292 22568
rect 32772 22584 32824 22636
rect 30380 22516 30432 22568
rect 25044 22448 25096 22500
rect 27252 22491 27304 22500
rect 27252 22457 27261 22491
rect 27261 22457 27295 22491
rect 27295 22457 27304 22491
rect 27252 22448 27304 22457
rect 32220 22448 32272 22500
rect 20812 22380 20864 22432
rect 21456 22423 21508 22432
rect 21456 22389 21465 22423
rect 21465 22389 21499 22423
rect 21499 22389 21508 22423
rect 21456 22380 21508 22389
rect 21824 22423 21876 22432
rect 21824 22389 21833 22423
rect 21833 22389 21867 22423
rect 21867 22389 21876 22423
rect 21824 22380 21876 22389
rect 24308 22380 24360 22432
rect 25136 22423 25188 22432
rect 25136 22389 25145 22423
rect 25145 22389 25179 22423
rect 25179 22389 25188 22423
rect 25136 22380 25188 22389
rect 27804 22423 27856 22432
rect 27804 22389 27813 22423
rect 27813 22389 27847 22423
rect 27847 22389 27856 22423
rect 27804 22380 27856 22389
rect 28356 22423 28408 22432
rect 28356 22389 28365 22423
rect 28365 22389 28399 22423
rect 28399 22389 28408 22423
rect 28356 22380 28408 22389
rect 28724 22380 28776 22432
rect 31116 22380 31168 22432
rect 31392 22380 31444 22432
rect 31760 22380 31812 22432
rect 5170 22278 5222 22330
rect 5234 22278 5286 22330
rect 5298 22278 5350 22330
rect 5362 22278 5414 22330
rect 5426 22278 5478 22330
rect 13611 22278 13663 22330
rect 13675 22278 13727 22330
rect 13739 22278 13791 22330
rect 13803 22278 13855 22330
rect 13867 22278 13919 22330
rect 22052 22278 22104 22330
rect 22116 22278 22168 22330
rect 22180 22278 22232 22330
rect 22244 22278 22296 22330
rect 22308 22278 22360 22330
rect 30493 22278 30545 22330
rect 30557 22278 30609 22330
rect 30621 22278 30673 22330
rect 30685 22278 30737 22330
rect 30749 22278 30801 22330
rect 17224 22176 17276 22228
rect 19984 22176 20036 22228
rect 20628 22176 20680 22228
rect 21364 22219 21416 22228
rect 21364 22185 21373 22219
rect 21373 22185 21407 22219
rect 21407 22185 21416 22219
rect 21364 22176 21416 22185
rect 17132 21972 17184 22024
rect 23112 22176 23164 22228
rect 25872 22176 25924 22228
rect 26700 22219 26752 22228
rect 26700 22185 26709 22219
rect 26709 22185 26743 22219
rect 26743 22185 26752 22219
rect 26700 22176 26752 22185
rect 30380 22176 30432 22228
rect 31208 22176 31260 22228
rect 32772 22176 32824 22228
rect 18604 22015 18656 22024
rect 18604 21981 18616 22015
rect 18616 21981 18650 22015
rect 18650 21981 18656 22015
rect 18604 21972 18656 21981
rect 18788 21972 18840 22024
rect 18972 21972 19024 22024
rect 26332 22040 26384 22092
rect 18328 21904 18380 21956
rect 17684 21836 17736 21888
rect 18512 21836 18564 21888
rect 19432 21904 19484 21956
rect 20352 21904 20404 21956
rect 18788 21836 18840 21888
rect 19892 21836 19944 21888
rect 20720 21836 20772 21888
rect 21824 21972 21876 22024
rect 24308 21972 24360 22024
rect 26148 22015 26200 22024
rect 26148 21981 26157 22015
rect 26157 21981 26191 22015
rect 26191 21981 26200 22015
rect 26148 21972 26200 21981
rect 26792 22040 26844 22092
rect 27252 22040 27304 22092
rect 28172 22015 28224 22024
rect 28172 21981 28181 22015
rect 28181 21981 28215 22015
rect 28215 21981 28224 22015
rect 28172 21972 28224 21981
rect 29920 22015 29972 22024
rect 29920 21981 29929 22015
rect 29929 21981 29963 22015
rect 29963 21981 29972 22015
rect 29920 21972 29972 21981
rect 21548 21879 21600 21888
rect 21548 21845 21557 21879
rect 21557 21845 21591 21879
rect 21591 21845 21600 21879
rect 21548 21836 21600 21845
rect 21916 21836 21968 21888
rect 22560 21836 22612 21888
rect 23388 21836 23440 21888
rect 24400 21879 24452 21888
rect 24400 21845 24409 21879
rect 24409 21845 24443 21879
rect 24443 21845 24452 21879
rect 24400 21836 24452 21845
rect 25320 21836 25372 21888
rect 25780 21947 25832 21956
rect 25780 21913 25798 21947
rect 25798 21913 25832 21947
rect 25780 21904 25832 21913
rect 26332 21904 26384 21956
rect 27528 21904 27580 21956
rect 29644 21904 29696 21956
rect 30472 22015 30524 22024
rect 30472 21981 30481 22015
rect 30481 21981 30515 22015
rect 30515 21981 30524 22015
rect 30472 21972 30524 21981
rect 31116 22015 31168 22024
rect 31116 21981 31125 22015
rect 31125 21981 31159 22015
rect 31159 21981 31168 22015
rect 31116 21972 31168 21981
rect 31208 22015 31260 22024
rect 31208 21981 31217 22015
rect 31217 21981 31251 22015
rect 31251 21981 31260 22015
rect 31208 21972 31260 21981
rect 31392 22015 31444 22024
rect 31392 21981 31401 22015
rect 31401 21981 31435 22015
rect 31435 21981 31444 22015
rect 31392 21972 31444 21981
rect 31760 22040 31812 22092
rect 31944 21972 31996 22024
rect 32220 21972 32272 22024
rect 34888 21972 34940 22024
rect 26884 21836 26936 21888
rect 28356 21879 28408 21888
rect 28356 21845 28365 21879
rect 28365 21845 28399 21879
rect 28399 21845 28408 21879
rect 28356 21836 28408 21845
rect 30196 21836 30248 21888
rect 30840 21836 30892 21888
rect 31300 21836 31352 21888
rect 33508 21879 33560 21888
rect 33508 21845 33517 21879
rect 33517 21845 33551 21879
rect 33551 21845 33560 21879
rect 33508 21836 33560 21845
rect 9390 21734 9442 21786
rect 9454 21734 9506 21786
rect 9518 21734 9570 21786
rect 9582 21734 9634 21786
rect 9646 21734 9698 21786
rect 17831 21734 17883 21786
rect 17895 21734 17947 21786
rect 17959 21734 18011 21786
rect 18023 21734 18075 21786
rect 18087 21734 18139 21786
rect 26272 21734 26324 21786
rect 26336 21734 26388 21786
rect 26400 21734 26452 21786
rect 26464 21734 26516 21786
rect 26528 21734 26580 21786
rect 34713 21734 34765 21786
rect 34777 21734 34829 21786
rect 34841 21734 34893 21786
rect 34905 21734 34957 21786
rect 34969 21734 35021 21786
rect 17684 21675 17736 21684
rect 17684 21641 17693 21675
rect 17693 21641 17727 21675
rect 17727 21641 17736 21675
rect 17684 21632 17736 21641
rect 18328 21675 18380 21684
rect 18328 21641 18355 21675
rect 18355 21641 18380 21675
rect 18328 21632 18380 21641
rect 17224 21564 17276 21616
rect 18512 21607 18564 21616
rect 18512 21573 18521 21607
rect 18521 21573 18555 21607
rect 18555 21573 18564 21607
rect 19616 21632 19668 21684
rect 20352 21675 20404 21684
rect 20352 21641 20361 21675
rect 20361 21641 20395 21675
rect 20395 21641 20404 21675
rect 20352 21632 20404 21641
rect 21640 21675 21692 21684
rect 21640 21641 21649 21675
rect 21649 21641 21683 21675
rect 21683 21641 21692 21675
rect 21640 21632 21692 21641
rect 22376 21675 22428 21684
rect 22376 21641 22385 21675
rect 22385 21641 22419 21675
rect 22419 21641 22428 21675
rect 22376 21632 22428 21641
rect 18512 21564 18564 21573
rect 18972 21564 19024 21616
rect 18696 21496 18748 21548
rect 19432 21539 19484 21548
rect 19432 21505 19441 21539
rect 19441 21505 19475 21539
rect 19475 21505 19484 21539
rect 19432 21496 19484 21505
rect 19708 21539 19760 21548
rect 19708 21505 19717 21539
rect 19717 21505 19751 21539
rect 19751 21505 19760 21539
rect 19708 21496 19760 21505
rect 19892 21539 19944 21548
rect 19892 21505 19901 21539
rect 19901 21505 19935 21539
rect 19935 21505 19944 21539
rect 19892 21496 19944 21505
rect 20260 21564 20312 21616
rect 18052 21292 18104 21344
rect 19800 21471 19852 21480
rect 19800 21437 19809 21471
rect 19809 21437 19843 21471
rect 19843 21437 19852 21471
rect 19800 21428 19852 21437
rect 20996 21496 21048 21548
rect 20720 21428 20772 21480
rect 21180 21539 21232 21548
rect 21180 21505 21189 21539
rect 21189 21505 21223 21539
rect 21223 21505 21232 21539
rect 21180 21496 21232 21505
rect 21916 21564 21968 21616
rect 24400 21564 24452 21616
rect 22560 21496 22612 21548
rect 23020 21539 23072 21548
rect 23020 21505 23029 21539
rect 23029 21505 23063 21539
rect 23063 21505 23072 21539
rect 23020 21496 23072 21505
rect 23940 21496 23992 21548
rect 24768 21632 24820 21684
rect 25596 21632 25648 21684
rect 25780 21632 25832 21684
rect 31116 21632 31168 21684
rect 33508 21632 33560 21684
rect 25044 21607 25096 21616
rect 25044 21573 25053 21607
rect 25053 21573 25087 21607
rect 25087 21573 25096 21607
rect 25044 21564 25096 21573
rect 25320 21564 25372 21616
rect 25136 21496 25188 21548
rect 28356 21564 28408 21616
rect 30196 21607 30248 21616
rect 30196 21573 30230 21607
rect 30230 21573 30248 21607
rect 30196 21564 30248 21573
rect 31208 21564 31260 21616
rect 21548 21428 21600 21480
rect 21916 21428 21968 21480
rect 23112 21471 23164 21480
rect 19616 21335 19668 21344
rect 19616 21301 19625 21335
rect 19625 21301 19659 21335
rect 19659 21301 19668 21335
rect 19616 21292 19668 21301
rect 20260 21335 20312 21344
rect 20260 21301 20269 21335
rect 20269 21301 20303 21335
rect 20303 21301 20312 21335
rect 20260 21292 20312 21301
rect 20444 21292 20496 21344
rect 20812 21292 20864 21344
rect 23112 21437 23121 21471
rect 23121 21437 23155 21471
rect 23155 21437 23164 21471
rect 23112 21428 23164 21437
rect 24768 21403 24820 21412
rect 24768 21369 24777 21403
rect 24777 21369 24811 21403
rect 24811 21369 24820 21403
rect 24768 21360 24820 21369
rect 25228 21403 25280 21412
rect 25228 21369 25237 21403
rect 25237 21369 25271 21403
rect 25271 21369 25280 21403
rect 25228 21360 25280 21369
rect 25596 21471 25648 21480
rect 25596 21437 25605 21471
rect 25605 21437 25639 21471
rect 25639 21437 25648 21471
rect 25596 21428 25648 21437
rect 26056 21471 26108 21480
rect 26056 21437 26065 21471
rect 26065 21437 26099 21471
rect 26099 21437 26108 21471
rect 26056 21428 26108 21437
rect 27068 21496 27120 21548
rect 29276 21496 29328 21548
rect 30012 21496 30064 21548
rect 32404 21539 32456 21548
rect 32404 21505 32413 21539
rect 32413 21505 32447 21539
rect 32447 21505 32456 21539
rect 32404 21496 32456 21505
rect 32772 21496 32824 21548
rect 31300 21403 31352 21412
rect 31300 21369 31309 21403
rect 31309 21369 31343 21403
rect 31343 21369 31352 21403
rect 31300 21360 31352 21369
rect 31760 21360 31812 21412
rect 33600 21471 33652 21480
rect 33600 21437 33609 21471
rect 33609 21437 33643 21471
rect 33643 21437 33652 21471
rect 33600 21428 33652 21437
rect 22836 21292 22888 21344
rect 24492 21335 24544 21344
rect 24492 21301 24501 21335
rect 24501 21301 24535 21335
rect 24535 21301 24544 21335
rect 24492 21292 24544 21301
rect 25136 21335 25188 21344
rect 25136 21301 25145 21335
rect 25145 21301 25179 21335
rect 25179 21301 25188 21335
rect 25136 21292 25188 21301
rect 26976 21335 27028 21344
rect 26976 21301 26985 21335
rect 26985 21301 27019 21335
rect 27019 21301 27028 21335
rect 26976 21292 27028 21301
rect 27988 21292 28040 21344
rect 32496 21335 32548 21344
rect 32496 21301 32505 21335
rect 32505 21301 32539 21335
rect 32539 21301 32548 21335
rect 32496 21292 32548 21301
rect 33508 21292 33560 21344
rect 5170 21190 5222 21242
rect 5234 21190 5286 21242
rect 5298 21190 5350 21242
rect 5362 21190 5414 21242
rect 5426 21190 5478 21242
rect 13611 21190 13663 21242
rect 13675 21190 13727 21242
rect 13739 21190 13791 21242
rect 13803 21190 13855 21242
rect 13867 21190 13919 21242
rect 22052 21190 22104 21242
rect 22116 21190 22168 21242
rect 22180 21190 22232 21242
rect 22244 21190 22296 21242
rect 22308 21190 22360 21242
rect 30493 21190 30545 21242
rect 30557 21190 30609 21242
rect 30621 21190 30673 21242
rect 30685 21190 30737 21242
rect 30749 21190 30801 21242
rect 19800 21088 19852 21140
rect 20444 21131 20496 21140
rect 20444 21097 20453 21131
rect 20453 21097 20487 21131
rect 20487 21097 20496 21131
rect 20444 21088 20496 21097
rect 21916 21131 21968 21140
rect 21916 21097 21925 21131
rect 21925 21097 21959 21131
rect 21959 21097 21968 21131
rect 21916 21088 21968 21097
rect 23020 21088 23072 21140
rect 18880 20952 18932 21004
rect 17684 20884 17736 20936
rect 17592 20816 17644 20868
rect 18052 20884 18104 20936
rect 20720 20952 20772 21004
rect 22560 20952 22612 21004
rect 27068 21131 27120 21140
rect 27068 21097 27077 21131
rect 27077 21097 27111 21131
rect 27111 21097 27120 21131
rect 27068 21088 27120 21097
rect 27344 21088 27396 21140
rect 29920 21088 29972 21140
rect 23940 21020 23992 21072
rect 24032 20952 24084 21004
rect 23940 20927 23992 20936
rect 23940 20893 23949 20927
rect 23949 20893 23983 20927
rect 23983 20893 23992 20927
rect 23940 20884 23992 20893
rect 24308 20952 24360 21004
rect 25136 20952 25188 21004
rect 26056 21020 26108 21072
rect 27712 21063 27764 21072
rect 27712 21029 27721 21063
rect 27721 21029 27755 21063
rect 27755 21029 27764 21063
rect 27712 21020 27764 21029
rect 25320 20927 25372 20936
rect 25320 20893 25329 20927
rect 25329 20893 25363 20927
rect 25363 20893 25372 20927
rect 25320 20884 25372 20893
rect 18236 20748 18288 20800
rect 18512 20748 18564 20800
rect 21180 20748 21232 20800
rect 21548 20748 21600 20800
rect 24584 20748 24636 20800
rect 25596 20884 25648 20936
rect 26608 20927 26660 20936
rect 26608 20893 26617 20927
rect 26617 20893 26651 20927
rect 26651 20893 26660 20927
rect 26608 20884 26660 20893
rect 30012 20952 30064 21004
rect 31944 21131 31996 21140
rect 31944 21097 31953 21131
rect 31953 21097 31987 21131
rect 31987 21097 31996 21131
rect 31944 21088 31996 21097
rect 32404 21088 32456 21140
rect 32772 21088 32824 21140
rect 26792 20927 26844 20936
rect 26792 20893 26801 20927
rect 26801 20893 26835 20927
rect 26835 20893 26844 20927
rect 26792 20884 26844 20893
rect 26976 20884 27028 20936
rect 27436 20927 27488 20936
rect 27436 20893 27445 20927
rect 27445 20893 27479 20927
rect 27479 20893 27488 20927
rect 27436 20884 27488 20893
rect 27804 20884 27856 20936
rect 27988 20884 28040 20936
rect 29276 20884 29328 20936
rect 30840 20927 30892 20936
rect 30840 20893 30874 20927
rect 30874 20893 30892 20927
rect 26700 20748 26752 20800
rect 28724 20748 28776 20800
rect 29000 20816 29052 20868
rect 30380 20816 30432 20868
rect 30840 20884 30892 20893
rect 30932 20816 30984 20868
rect 33324 20816 33376 20868
rect 31944 20748 31996 20800
rect 9390 20646 9442 20698
rect 9454 20646 9506 20698
rect 9518 20646 9570 20698
rect 9582 20646 9634 20698
rect 9646 20646 9698 20698
rect 17831 20646 17883 20698
rect 17895 20646 17947 20698
rect 17959 20646 18011 20698
rect 18023 20646 18075 20698
rect 18087 20646 18139 20698
rect 26272 20646 26324 20698
rect 26336 20646 26388 20698
rect 26400 20646 26452 20698
rect 26464 20646 26516 20698
rect 26528 20646 26580 20698
rect 34713 20646 34765 20698
rect 34777 20646 34829 20698
rect 34841 20646 34893 20698
rect 34905 20646 34957 20698
rect 34969 20646 35021 20698
rect 17132 20544 17184 20596
rect 17776 20544 17828 20596
rect 18236 20544 18288 20596
rect 19616 20544 19668 20596
rect 19708 20544 19760 20596
rect 17592 20408 17644 20460
rect 17684 20272 17736 20324
rect 17960 20383 18012 20392
rect 17960 20349 17969 20383
rect 17969 20349 18003 20383
rect 18003 20349 18012 20383
rect 17960 20340 18012 20349
rect 19708 20451 19760 20460
rect 19708 20417 19717 20451
rect 19717 20417 19751 20451
rect 19751 20417 19760 20451
rect 19708 20408 19760 20417
rect 23020 20544 23072 20596
rect 26608 20544 26660 20596
rect 27712 20587 27764 20596
rect 27712 20553 27721 20587
rect 27721 20553 27755 20587
rect 27755 20553 27764 20587
rect 27712 20544 27764 20553
rect 27804 20587 27856 20596
rect 27804 20553 27813 20587
rect 27813 20553 27847 20587
rect 27847 20553 27856 20587
rect 27804 20544 27856 20553
rect 29000 20544 29052 20596
rect 22468 20476 22520 20528
rect 20260 20408 20312 20460
rect 22652 20408 22704 20460
rect 23204 20408 23256 20460
rect 23480 20451 23532 20460
rect 23480 20417 23489 20451
rect 23489 20417 23523 20451
rect 23523 20417 23532 20451
rect 23480 20408 23532 20417
rect 23664 20408 23716 20460
rect 26884 20476 26936 20528
rect 26148 20451 26200 20460
rect 26148 20417 26157 20451
rect 26157 20417 26191 20451
rect 26191 20417 26200 20451
rect 26148 20408 26200 20417
rect 27160 20451 27212 20460
rect 27160 20417 27169 20451
rect 27169 20417 27203 20451
rect 27203 20417 27212 20451
rect 27160 20408 27212 20417
rect 27436 20451 27488 20460
rect 27436 20417 27445 20451
rect 27445 20417 27479 20451
rect 27479 20417 27488 20451
rect 27436 20408 27488 20417
rect 27896 20451 27948 20460
rect 27896 20417 27905 20451
rect 27905 20417 27939 20451
rect 27939 20417 27948 20451
rect 27896 20408 27948 20417
rect 30564 20476 30616 20528
rect 32496 20544 32548 20596
rect 33324 20587 33376 20596
rect 33324 20553 33333 20587
rect 33333 20553 33367 20587
rect 33367 20553 33376 20587
rect 33324 20544 33376 20553
rect 32864 20519 32916 20528
rect 28172 20451 28224 20460
rect 28172 20417 28181 20451
rect 28181 20417 28215 20451
rect 28215 20417 28224 20451
rect 28172 20408 28224 20417
rect 32864 20485 32873 20519
rect 32873 20485 32907 20519
rect 32907 20485 32916 20519
rect 32864 20476 32916 20485
rect 31208 20408 31260 20460
rect 31944 20408 31996 20460
rect 32404 20451 32456 20460
rect 32404 20417 32413 20451
rect 32413 20417 32447 20451
rect 32447 20417 32456 20451
rect 32404 20408 32456 20417
rect 33232 20451 33284 20460
rect 33232 20417 33241 20451
rect 33241 20417 33275 20451
rect 33275 20417 33284 20451
rect 33232 20408 33284 20417
rect 33508 20451 33560 20460
rect 33508 20417 33517 20451
rect 33517 20417 33551 20451
rect 33551 20417 33560 20451
rect 33508 20408 33560 20417
rect 27988 20272 28040 20324
rect 18144 20204 18196 20256
rect 19340 20247 19392 20256
rect 19340 20213 19349 20247
rect 19349 20213 19383 20247
rect 19383 20213 19392 20247
rect 19340 20204 19392 20213
rect 19432 20247 19484 20256
rect 19432 20213 19441 20247
rect 19441 20213 19475 20247
rect 19475 20213 19484 20247
rect 19432 20204 19484 20213
rect 22744 20247 22796 20256
rect 22744 20213 22753 20247
rect 22753 20213 22787 20247
rect 22787 20213 22796 20247
rect 22744 20204 22796 20213
rect 23112 20247 23164 20256
rect 23112 20213 23121 20247
rect 23121 20213 23155 20247
rect 23155 20213 23164 20247
rect 23112 20204 23164 20213
rect 26424 20247 26476 20256
rect 26424 20213 26433 20247
rect 26433 20213 26467 20247
rect 26467 20213 26476 20247
rect 26424 20204 26476 20213
rect 26976 20247 27028 20256
rect 26976 20213 26985 20247
rect 26985 20213 27019 20247
rect 27019 20213 27028 20247
rect 26976 20204 27028 20213
rect 31392 20247 31444 20256
rect 31392 20213 31401 20247
rect 31401 20213 31435 20247
rect 31435 20213 31444 20247
rect 31392 20204 31444 20213
rect 32220 20383 32272 20392
rect 32220 20349 32229 20383
rect 32229 20349 32263 20383
rect 32263 20349 32272 20383
rect 32220 20340 32272 20349
rect 32312 20272 32364 20324
rect 32588 20204 32640 20256
rect 33048 20247 33100 20256
rect 33048 20213 33057 20247
rect 33057 20213 33091 20247
rect 33091 20213 33100 20247
rect 33048 20204 33100 20213
rect 5170 20102 5222 20154
rect 5234 20102 5286 20154
rect 5298 20102 5350 20154
rect 5362 20102 5414 20154
rect 5426 20102 5478 20154
rect 13611 20102 13663 20154
rect 13675 20102 13727 20154
rect 13739 20102 13791 20154
rect 13803 20102 13855 20154
rect 13867 20102 13919 20154
rect 22052 20102 22104 20154
rect 22116 20102 22168 20154
rect 22180 20102 22232 20154
rect 22244 20102 22296 20154
rect 22308 20102 22360 20154
rect 30493 20102 30545 20154
rect 30557 20102 30609 20154
rect 30621 20102 30673 20154
rect 30685 20102 30737 20154
rect 30749 20102 30801 20154
rect 17684 20000 17736 20052
rect 18144 20043 18196 20052
rect 18144 20009 18153 20043
rect 18153 20009 18187 20043
rect 18187 20009 18196 20043
rect 18144 20000 18196 20009
rect 19340 20000 19392 20052
rect 19708 20000 19760 20052
rect 22468 20000 22520 20052
rect 22744 20000 22796 20052
rect 23204 20000 23256 20052
rect 26424 20000 26476 20052
rect 26792 20043 26844 20052
rect 26792 20009 26801 20043
rect 26801 20009 26835 20043
rect 26835 20009 26844 20043
rect 26792 20000 26844 20009
rect 27804 20000 27856 20052
rect 29184 20000 29236 20052
rect 29552 20043 29604 20052
rect 29552 20009 29561 20043
rect 29561 20009 29595 20043
rect 29595 20009 29604 20043
rect 29552 20000 29604 20009
rect 31208 20000 31260 20052
rect 940 19796 992 19848
rect 17684 19839 17736 19848
rect 17684 19805 17693 19839
rect 17693 19805 17727 19839
rect 17727 19805 17736 19839
rect 17684 19796 17736 19805
rect 18512 19771 18564 19780
rect 18512 19737 18539 19771
rect 18539 19737 18564 19771
rect 18512 19728 18564 19737
rect 18696 19771 18748 19780
rect 18696 19737 18705 19771
rect 18705 19737 18739 19771
rect 18739 19737 18748 19771
rect 18696 19728 18748 19737
rect 19800 19932 19852 19984
rect 21916 19932 21968 19984
rect 22192 19907 22244 19916
rect 20076 19839 20128 19848
rect 20076 19805 20085 19839
rect 20085 19805 20119 19839
rect 20119 19805 20128 19839
rect 20076 19796 20128 19805
rect 21180 19839 21232 19848
rect 21180 19805 21189 19839
rect 21189 19805 21223 19839
rect 21223 19805 21232 19839
rect 21180 19796 21232 19805
rect 18236 19660 18288 19712
rect 18328 19703 18380 19712
rect 18328 19669 18337 19703
rect 18337 19669 18371 19703
rect 18371 19669 18380 19703
rect 18328 19660 18380 19669
rect 19248 19703 19300 19712
rect 19248 19669 19257 19703
rect 19257 19669 19291 19703
rect 19291 19669 19300 19703
rect 19248 19660 19300 19669
rect 20720 19660 20772 19712
rect 21364 19703 21416 19712
rect 21364 19669 21373 19703
rect 21373 19669 21407 19703
rect 21407 19669 21416 19703
rect 21364 19660 21416 19669
rect 22192 19873 22201 19907
rect 22201 19873 22235 19907
rect 22235 19873 22244 19907
rect 22192 19864 22244 19873
rect 22376 19796 22428 19848
rect 22836 19907 22888 19916
rect 22836 19873 22845 19907
rect 22845 19873 22879 19907
rect 22879 19873 22888 19907
rect 22836 19864 22888 19873
rect 23112 19839 23164 19848
rect 23112 19805 23146 19839
rect 23146 19805 23164 19839
rect 23112 19796 23164 19805
rect 32404 19975 32456 19984
rect 32404 19941 32413 19975
rect 32413 19941 32447 19975
rect 32447 19941 32456 19975
rect 32404 19932 32456 19941
rect 30932 19907 30984 19916
rect 30932 19873 30941 19907
rect 30941 19873 30975 19907
rect 30975 19873 30984 19907
rect 30932 19864 30984 19873
rect 32128 19864 32180 19916
rect 25872 19728 25924 19780
rect 26976 19796 27028 19848
rect 32220 19796 32272 19848
rect 33140 19839 33192 19848
rect 33140 19805 33149 19839
rect 33149 19805 33183 19839
rect 33183 19805 33192 19839
rect 33140 19796 33192 19805
rect 33508 20043 33560 20052
rect 33508 20009 33517 20043
rect 33517 20009 33551 20043
rect 33551 20009 33560 20043
rect 33508 20000 33560 20009
rect 33600 19796 33652 19848
rect 29368 19728 29420 19780
rect 31392 19728 31444 19780
rect 21732 19660 21784 19712
rect 22928 19660 22980 19712
rect 32588 19660 32640 19712
rect 32864 19703 32916 19712
rect 32864 19669 32873 19703
rect 32873 19669 32907 19703
rect 32907 19669 32916 19703
rect 32864 19660 32916 19669
rect 9390 19558 9442 19610
rect 9454 19558 9506 19610
rect 9518 19558 9570 19610
rect 9582 19558 9634 19610
rect 9646 19558 9698 19610
rect 17831 19558 17883 19610
rect 17895 19558 17947 19610
rect 17959 19558 18011 19610
rect 18023 19558 18075 19610
rect 18087 19558 18139 19610
rect 26272 19558 26324 19610
rect 26336 19558 26388 19610
rect 26400 19558 26452 19610
rect 26464 19558 26516 19610
rect 26528 19558 26580 19610
rect 34713 19558 34765 19610
rect 34777 19558 34829 19610
rect 34841 19558 34893 19610
rect 34905 19558 34957 19610
rect 34969 19558 35021 19610
rect 19248 19456 19300 19508
rect 19432 19456 19484 19508
rect 20076 19456 20128 19508
rect 17132 19184 17184 19236
rect 18328 19320 18380 19372
rect 18696 19320 18748 19372
rect 18236 19252 18288 19304
rect 18972 19363 19024 19372
rect 18972 19329 18981 19363
rect 18981 19329 19015 19363
rect 19015 19329 19024 19363
rect 18972 19320 19024 19329
rect 19340 19252 19392 19304
rect 20904 19388 20956 19440
rect 19708 19320 19760 19372
rect 20168 19320 20220 19372
rect 21364 19456 21416 19508
rect 21916 19456 21968 19508
rect 21824 19388 21876 19440
rect 21088 19320 21140 19372
rect 21456 19320 21508 19372
rect 23020 19388 23072 19440
rect 24860 19456 24912 19508
rect 25688 19456 25740 19508
rect 27160 19456 27212 19508
rect 29368 19499 29420 19508
rect 29368 19465 29377 19499
rect 29377 19465 29411 19499
rect 29411 19465 29420 19499
rect 29368 19456 29420 19465
rect 22376 19320 22428 19372
rect 22744 19320 22796 19372
rect 23388 19363 23440 19372
rect 23388 19329 23397 19363
rect 23397 19329 23431 19363
rect 23431 19329 23440 19363
rect 23388 19320 23440 19329
rect 23848 19320 23900 19372
rect 24860 19363 24912 19372
rect 24860 19329 24869 19363
rect 24869 19329 24903 19363
rect 24903 19329 24912 19363
rect 24860 19320 24912 19329
rect 25044 19320 25096 19372
rect 25504 19320 25556 19372
rect 26792 19320 26844 19372
rect 28172 19388 28224 19440
rect 21364 19295 21416 19304
rect 21364 19261 21373 19295
rect 21373 19261 21407 19295
rect 21407 19261 21416 19295
rect 21364 19252 21416 19261
rect 22192 19184 22244 19236
rect 18236 19116 18288 19168
rect 19156 19116 19208 19168
rect 22468 19116 22520 19168
rect 22560 19159 22612 19168
rect 22560 19125 22569 19159
rect 22569 19125 22603 19159
rect 22603 19125 22612 19159
rect 22560 19116 22612 19125
rect 23664 19116 23716 19168
rect 25596 19116 25648 19168
rect 26148 19116 26200 19168
rect 28264 19363 28316 19372
rect 28264 19329 28273 19363
rect 28273 19329 28307 19363
rect 28307 19329 28316 19363
rect 28264 19320 28316 19329
rect 28724 19363 28776 19372
rect 28724 19329 28733 19363
rect 28733 19329 28767 19363
rect 28767 19329 28776 19363
rect 28724 19320 28776 19329
rect 29276 19388 29328 19440
rect 31944 19499 31996 19508
rect 31944 19465 31953 19499
rect 31953 19465 31987 19499
rect 31987 19465 31996 19499
rect 31944 19456 31996 19465
rect 32864 19456 32916 19508
rect 33140 19456 33192 19508
rect 33048 19388 33100 19440
rect 29000 19363 29052 19372
rect 29000 19329 29009 19363
rect 29009 19329 29043 19363
rect 29043 19329 29052 19363
rect 29000 19320 29052 19329
rect 29092 19363 29144 19372
rect 29092 19329 29101 19363
rect 29101 19329 29135 19363
rect 29135 19329 29144 19363
rect 29092 19320 29144 19329
rect 31208 19320 31260 19372
rect 32312 19295 32364 19304
rect 28448 19159 28500 19168
rect 28448 19125 28457 19159
rect 28457 19125 28491 19159
rect 28491 19125 28500 19159
rect 28448 19116 28500 19125
rect 30840 19116 30892 19168
rect 32312 19261 32321 19295
rect 32321 19261 32355 19295
rect 32355 19261 32364 19295
rect 32312 19252 32364 19261
rect 5170 19014 5222 19066
rect 5234 19014 5286 19066
rect 5298 19014 5350 19066
rect 5362 19014 5414 19066
rect 5426 19014 5478 19066
rect 13611 19014 13663 19066
rect 13675 19014 13727 19066
rect 13739 19014 13791 19066
rect 13803 19014 13855 19066
rect 13867 19014 13919 19066
rect 22052 19014 22104 19066
rect 22116 19014 22168 19066
rect 22180 19014 22232 19066
rect 22244 19014 22296 19066
rect 22308 19014 22360 19066
rect 30493 19014 30545 19066
rect 30557 19014 30609 19066
rect 30621 19014 30673 19066
rect 30685 19014 30737 19066
rect 30749 19014 30801 19066
rect 18328 18912 18380 18964
rect 18972 18955 19024 18964
rect 18972 18921 18981 18955
rect 18981 18921 19015 18955
rect 19015 18921 19024 18955
rect 18972 18912 19024 18921
rect 19708 18912 19760 18964
rect 20168 18955 20220 18964
rect 20168 18921 20177 18955
rect 20177 18921 20211 18955
rect 20211 18921 20220 18955
rect 20168 18912 20220 18921
rect 20536 18912 20588 18964
rect 20812 18912 20864 18964
rect 21456 18912 21508 18964
rect 21732 18955 21784 18964
rect 21732 18921 21741 18955
rect 21741 18921 21775 18955
rect 21775 18921 21784 18955
rect 21732 18912 21784 18921
rect 22928 18955 22980 18964
rect 22928 18921 22937 18955
rect 22937 18921 22971 18955
rect 22971 18921 22980 18955
rect 22928 18912 22980 18921
rect 23572 18912 23624 18964
rect 23848 18955 23900 18964
rect 23848 18921 23857 18955
rect 23857 18921 23891 18955
rect 23891 18921 23900 18955
rect 23848 18912 23900 18921
rect 28264 18912 28316 18964
rect 29000 18912 29052 18964
rect 29644 18912 29696 18964
rect 16212 18708 16264 18760
rect 18972 18776 19024 18828
rect 17224 18708 17276 18760
rect 17684 18572 17736 18624
rect 19156 18708 19208 18760
rect 19340 18708 19392 18760
rect 19616 18751 19668 18760
rect 19616 18717 19625 18751
rect 19625 18717 19659 18751
rect 19659 18717 19668 18751
rect 19616 18708 19668 18717
rect 19800 18751 19852 18760
rect 19800 18717 19809 18751
rect 19809 18717 19843 18751
rect 19843 18717 19852 18751
rect 19800 18708 19852 18717
rect 21088 18776 21140 18828
rect 21456 18819 21508 18828
rect 21456 18785 21465 18819
rect 21465 18785 21499 18819
rect 21499 18785 21508 18819
rect 21456 18776 21508 18785
rect 21548 18819 21600 18828
rect 21548 18785 21557 18819
rect 21557 18785 21591 18819
rect 21591 18785 21600 18819
rect 21548 18776 21600 18785
rect 20536 18751 20588 18760
rect 20536 18717 20545 18751
rect 20545 18717 20579 18751
rect 20579 18717 20588 18751
rect 20536 18708 20588 18717
rect 20720 18708 20772 18760
rect 21824 18751 21876 18760
rect 21824 18717 21833 18751
rect 21833 18717 21867 18751
rect 21867 18717 21876 18751
rect 21824 18708 21876 18717
rect 22560 18776 22612 18828
rect 22652 18708 22704 18760
rect 26608 18776 26660 18828
rect 29092 18776 29144 18828
rect 31208 18955 31260 18964
rect 31208 18921 31217 18955
rect 31217 18921 31251 18955
rect 31251 18921 31260 18955
rect 31208 18912 31260 18921
rect 33232 18912 33284 18964
rect 23480 18751 23532 18760
rect 23480 18717 23489 18751
rect 23489 18717 23523 18751
rect 23523 18717 23532 18751
rect 23480 18708 23532 18717
rect 23664 18708 23716 18760
rect 26884 18708 26936 18760
rect 23940 18640 23992 18692
rect 19984 18615 20036 18624
rect 19984 18581 19993 18615
rect 19993 18581 20027 18615
rect 20027 18581 20036 18615
rect 19984 18572 20036 18581
rect 20720 18572 20772 18624
rect 21180 18572 21232 18624
rect 21640 18572 21692 18624
rect 21916 18572 21968 18624
rect 23664 18572 23716 18624
rect 27436 18708 27488 18760
rect 29552 18708 29604 18760
rect 27620 18683 27672 18692
rect 27620 18649 27654 18683
rect 27654 18649 27672 18683
rect 27620 18640 27672 18649
rect 29184 18640 29236 18692
rect 30104 18751 30156 18760
rect 30104 18717 30113 18751
rect 30113 18717 30147 18751
rect 30147 18717 30156 18751
rect 30104 18708 30156 18717
rect 32128 18776 32180 18828
rect 28540 18572 28592 18624
rect 29460 18572 29512 18624
rect 30932 18708 30984 18760
rect 31300 18708 31352 18760
rect 31944 18708 31996 18760
rect 30380 18615 30432 18624
rect 30380 18581 30389 18615
rect 30389 18581 30423 18615
rect 30423 18581 30432 18615
rect 30380 18572 30432 18581
rect 9390 18470 9442 18522
rect 9454 18470 9506 18522
rect 9518 18470 9570 18522
rect 9582 18470 9634 18522
rect 9646 18470 9698 18522
rect 17831 18470 17883 18522
rect 17895 18470 17947 18522
rect 17959 18470 18011 18522
rect 18023 18470 18075 18522
rect 18087 18470 18139 18522
rect 26272 18470 26324 18522
rect 26336 18470 26388 18522
rect 26400 18470 26452 18522
rect 26464 18470 26516 18522
rect 26528 18470 26580 18522
rect 34713 18470 34765 18522
rect 34777 18470 34829 18522
rect 34841 18470 34893 18522
rect 34905 18470 34957 18522
rect 34969 18470 35021 18522
rect 17224 18368 17276 18420
rect 17132 18232 17184 18284
rect 18328 18368 18380 18420
rect 19616 18368 19668 18420
rect 19984 18368 20036 18420
rect 20720 18368 20772 18420
rect 21640 18368 21692 18420
rect 25504 18411 25556 18420
rect 25504 18377 25513 18411
rect 25513 18377 25547 18411
rect 25547 18377 25556 18411
rect 25504 18368 25556 18377
rect 27620 18368 27672 18420
rect 18236 18232 18288 18284
rect 18788 18275 18840 18284
rect 18788 18241 18797 18275
rect 18797 18241 18831 18275
rect 18831 18241 18840 18275
rect 18788 18232 18840 18241
rect 17684 18207 17736 18216
rect 17684 18173 17693 18207
rect 17693 18173 17727 18207
rect 17727 18173 17736 18207
rect 17684 18164 17736 18173
rect 19340 18300 19392 18352
rect 19800 18300 19852 18352
rect 20720 18232 20772 18284
rect 21548 18232 21600 18284
rect 22376 18232 22428 18284
rect 22468 18232 22520 18284
rect 24952 18275 25004 18284
rect 24952 18241 24961 18275
rect 24961 18241 24995 18275
rect 24995 18241 25004 18275
rect 24952 18232 25004 18241
rect 17500 18028 17552 18080
rect 20812 18096 20864 18148
rect 25872 18275 25924 18284
rect 25872 18241 25881 18275
rect 25881 18241 25915 18275
rect 25915 18241 25924 18275
rect 25872 18232 25924 18241
rect 26056 18232 26108 18284
rect 26516 18232 26568 18284
rect 26700 18232 26752 18284
rect 26976 18275 27028 18284
rect 26976 18241 26985 18275
rect 26985 18241 27019 18275
rect 27019 18241 27028 18275
rect 26976 18232 27028 18241
rect 27528 18232 27580 18284
rect 29460 18368 29512 18420
rect 29644 18411 29696 18420
rect 29644 18377 29653 18411
rect 29653 18377 29687 18411
rect 29687 18377 29696 18411
rect 29644 18368 29696 18377
rect 29736 18411 29788 18420
rect 29736 18377 29745 18411
rect 29745 18377 29779 18411
rect 29779 18377 29788 18411
rect 29736 18368 29788 18377
rect 30104 18368 30156 18420
rect 28448 18300 28500 18352
rect 30380 18232 30432 18284
rect 25780 18096 25832 18148
rect 18420 18028 18472 18080
rect 18512 18071 18564 18080
rect 18512 18037 18521 18071
rect 18521 18037 18555 18071
rect 18555 18037 18564 18071
rect 18512 18028 18564 18037
rect 22744 18071 22796 18080
rect 22744 18037 22753 18071
rect 22753 18037 22787 18071
rect 22787 18037 22796 18071
rect 22744 18028 22796 18037
rect 24676 18028 24728 18080
rect 26240 18071 26292 18080
rect 26240 18037 26249 18071
rect 26249 18037 26283 18071
rect 26283 18037 26292 18071
rect 26240 18028 26292 18037
rect 27896 18028 27948 18080
rect 30840 18028 30892 18080
rect 31392 18028 31444 18080
rect 5170 17926 5222 17978
rect 5234 17926 5286 17978
rect 5298 17926 5350 17978
rect 5362 17926 5414 17978
rect 5426 17926 5478 17978
rect 13611 17926 13663 17978
rect 13675 17926 13727 17978
rect 13739 17926 13791 17978
rect 13803 17926 13855 17978
rect 13867 17926 13919 17978
rect 22052 17926 22104 17978
rect 22116 17926 22168 17978
rect 22180 17926 22232 17978
rect 22244 17926 22296 17978
rect 22308 17926 22360 17978
rect 30493 17926 30545 17978
rect 30557 17926 30609 17978
rect 30621 17926 30673 17978
rect 30685 17926 30737 17978
rect 30749 17926 30801 17978
rect 17500 17867 17552 17876
rect 17500 17833 17509 17867
rect 17509 17833 17543 17867
rect 17543 17833 17552 17867
rect 17500 17824 17552 17833
rect 18144 17824 18196 17876
rect 19340 17867 19392 17876
rect 19340 17833 19349 17867
rect 19349 17833 19383 17867
rect 19383 17833 19392 17867
rect 19340 17824 19392 17833
rect 16120 17688 16172 17740
rect 15568 17663 15620 17672
rect 15568 17629 15577 17663
rect 15577 17629 15611 17663
rect 15611 17629 15620 17663
rect 15568 17620 15620 17629
rect 22100 17824 22152 17876
rect 16120 17552 16172 17604
rect 17132 17527 17184 17536
rect 17132 17493 17141 17527
rect 17141 17493 17175 17527
rect 17175 17493 17184 17527
rect 17132 17484 17184 17493
rect 21456 17688 21508 17740
rect 22560 17824 22612 17876
rect 22744 17824 22796 17876
rect 23112 17867 23164 17876
rect 23112 17833 23121 17867
rect 23121 17833 23155 17867
rect 23155 17833 23164 17867
rect 23112 17824 23164 17833
rect 23940 17867 23992 17876
rect 23940 17833 23949 17867
rect 23949 17833 23983 17867
rect 23983 17833 23992 17867
rect 23940 17824 23992 17833
rect 25780 17867 25832 17876
rect 25780 17833 25789 17867
rect 25789 17833 25823 17867
rect 25823 17833 25832 17867
rect 25780 17824 25832 17833
rect 29460 17824 29512 17876
rect 30380 17824 30432 17876
rect 22468 17756 22520 17808
rect 23296 17756 23348 17808
rect 30288 17756 30340 17808
rect 20260 17663 20312 17672
rect 20260 17629 20269 17663
rect 20269 17629 20303 17663
rect 20303 17629 20312 17663
rect 20260 17620 20312 17629
rect 20628 17620 20680 17672
rect 20812 17663 20864 17672
rect 20812 17629 20821 17663
rect 20821 17629 20855 17663
rect 20855 17629 20864 17663
rect 20812 17620 20864 17629
rect 20996 17663 21048 17672
rect 20996 17629 21005 17663
rect 21005 17629 21039 17663
rect 21039 17629 21048 17663
rect 20996 17620 21048 17629
rect 18236 17484 18288 17536
rect 18420 17484 18472 17536
rect 19708 17484 19760 17536
rect 20076 17527 20128 17536
rect 20076 17493 20085 17527
rect 20085 17493 20119 17527
rect 20119 17493 20128 17527
rect 20076 17484 20128 17493
rect 20168 17484 20220 17536
rect 20352 17527 20404 17536
rect 20352 17493 20361 17527
rect 20361 17493 20395 17527
rect 20395 17493 20404 17527
rect 20352 17484 20404 17493
rect 20904 17552 20956 17604
rect 21732 17620 21784 17672
rect 21916 17620 21968 17672
rect 22376 17620 22428 17672
rect 22928 17663 22980 17672
rect 22928 17629 22937 17663
rect 22937 17629 22971 17663
rect 22971 17629 22980 17663
rect 22928 17620 22980 17629
rect 23204 17663 23256 17672
rect 23204 17629 23213 17663
rect 23213 17629 23247 17663
rect 23247 17629 23256 17663
rect 23204 17620 23256 17629
rect 23296 17663 23348 17672
rect 23296 17629 23305 17663
rect 23305 17629 23339 17663
rect 23339 17629 23348 17663
rect 23296 17620 23348 17629
rect 23572 17620 23624 17672
rect 24308 17620 24360 17672
rect 24676 17663 24728 17672
rect 24676 17629 24710 17663
rect 24710 17629 24728 17663
rect 24676 17620 24728 17629
rect 25044 17552 25096 17604
rect 27896 17620 27948 17672
rect 25964 17552 26016 17604
rect 31392 17620 31444 17672
rect 30840 17552 30892 17604
rect 21456 17527 21508 17536
rect 21456 17493 21465 17527
rect 21465 17493 21499 17527
rect 21499 17493 21508 17527
rect 21456 17484 21508 17493
rect 21824 17484 21876 17536
rect 22284 17527 22336 17536
rect 22284 17493 22293 17527
rect 22293 17493 22327 17527
rect 22327 17493 22336 17527
rect 22284 17484 22336 17493
rect 22744 17527 22796 17536
rect 22744 17493 22753 17527
rect 22753 17493 22787 17527
rect 22787 17493 22796 17527
rect 22744 17484 22796 17493
rect 27252 17527 27304 17536
rect 27252 17493 27261 17527
rect 27261 17493 27295 17527
rect 27295 17493 27304 17527
rect 27252 17484 27304 17493
rect 27344 17527 27396 17536
rect 27344 17493 27353 17527
rect 27353 17493 27387 17527
rect 27387 17493 27396 17527
rect 27344 17484 27396 17493
rect 28540 17484 28592 17536
rect 9390 17382 9442 17434
rect 9454 17382 9506 17434
rect 9518 17382 9570 17434
rect 9582 17382 9634 17434
rect 9646 17382 9698 17434
rect 17831 17382 17883 17434
rect 17895 17382 17947 17434
rect 17959 17382 18011 17434
rect 18023 17382 18075 17434
rect 18087 17382 18139 17434
rect 26272 17382 26324 17434
rect 26336 17382 26388 17434
rect 26400 17382 26452 17434
rect 26464 17382 26516 17434
rect 26528 17382 26580 17434
rect 34713 17382 34765 17434
rect 34777 17382 34829 17434
rect 34841 17382 34893 17434
rect 34905 17382 34957 17434
rect 34969 17382 35021 17434
rect 15568 17280 15620 17332
rect 16120 17280 16172 17332
rect 17132 17280 17184 17332
rect 18236 17280 18288 17332
rect 16028 17212 16080 17264
rect 18512 17212 18564 17264
rect 16212 17144 16264 17196
rect 18420 17187 18472 17196
rect 18420 17153 18425 17187
rect 18425 17153 18459 17187
rect 18459 17153 18472 17187
rect 18420 17144 18472 17153
rect 18788 17280 18840 17332
rect 19984 17280 20036 17332
rect 20260 17280 20312 17332
rect 20352 17280 20404 17332
rect 20812 17280 20864 17332
rect 19432 17144 19484 17196
rect 19708 17187 19760 17196
rect 19708 17153 19717 17187
rect 19717 17153 19751 17187
rect 19751 17153 19760 17187
rect 19708 17144 19760 17153
rect 20076 17187 20128 17196
rect 18972 17119 19024 17128
rect 18972 17085 18981 17119
rect 18981 17085 19015 17119
rect 19015 17085 19024 17119
rect 18972 17076 19024 17085
rect 20076 17153 20085 17187
rect 20085 17153 20119 17187
rect 20119 17153 20128 17187
rect 20076 17144 20128 17153
rect 20444 17144 20496 17196
rect 20536 17187 20588 17196
rect 20536 17153 20545 17187
rect 20545 17153 20579 17187
rect 20579 17153 20588 17187
rect 20536 17144 20588 17153
rect 21824 17144 21876 17196
rect 18236 16940 18288 16992
rect 19340 16983 19392 16992
rect 19340 16949 19349 16983
rect 19349 16949 19383 16983
rect 19383 16949 19392 16983
rect 19340 16940 19392 16949
rect 19708 16940 19760 16992
rect 21640 17119 21692 17128
rect 21640 17085 21649 17119
rect 21649 17085 21683 17119
rect 21683 17085 21692 17119
rect 22284 17187 22336 17196
rect 22284 17153 22293 17187
rect 22293 17153 22327 17187
rect 22327 17153 22336 17187
rect 22284 17144 22336 17153
rect 22376 17144 22428 17196
rect 22468 17187 22520 17196
rect 22468 17153 22477 17187
rect 22477 17153 22511 17187
rect 22511 17153 22520 17187
rect 22468 17144 22520 17153
rect 22744 17280 22796 17332
rect 22836 17280 22888 17332
rect 24400 17280 24452 17332
rect 24952 17280 25004 17332
rect 25596 17280 25648 17332
rect 22836 17144 22888 17196
rect 23020 17187 23072 17196
rect 23020 17153 23029 17187
rect 23029 17153 23063 17187
rect 23063 17153 23072 17187
rect 23020 17144 23072 17153
rect 23572 17212 23624 17264
rect 25872 17323 25924 17332
rect 25872 17289 25881 17323
rect 25881 17289 25915 17323
rect 25915 17289 25924 17323
rect 25872 17280 25924 17289
rect 25964 17280 26016 17332
rect 26148 17280 26200 17332
rect 26608 17280 26660 17332
rect 26976 17323 27028 17332
rect 26976 17289 26985 17323
rect 26985 17289 27019 17323
rect 27019 17289 27028 17323
rect 26976 17280 27028 17289
rect 27252 17280 27304 17332
rect 29276 17323 29328 17332
rect 29276 17289 29285 17323
rect 29285 17289 29319 17323
rect 29319 17289 29328 17323
rect 29276 17280 29328 17289
rect 29552 17280 29604 17332
rect 29644 17280 29696 17332
rect 29736 17323 29788 17332
rect 29736 17289 29745 17323
rect 29745 17289 29779 17323
rect 29779 17289 29788 17323
rect 29736 17280 29788 17289
rect 30840 17323 30892 17332
rect 30840 17289 30849 17323
rect 30849 17289 30883 17323
rect 30883 17289 30892 17323
rect 30840 17280 30892 17289
rect 23388 17144 23440 17196
rect 24860 17144 24912 17196
rect 25228 17187 25280 17196
rect 25228 17153 25237 17187
rect 25237 17153 25271 17187
rect 25271 17153 25280 17187
rect 25228 17144 25280 17153
rect 26148 17187 26200 17196
rect 26148 17153 26157 17187
rect 26157 17153 26191 17187
rect 26191 17153 26200 17187
rect 26148 17144 26200 17153
rect 26240 17144 26292 17196
rect 26976 17144 27028 17196
rect 21640 17076 21692 17085
rect 21088 16940 21140 16992
rect 21732 16940 21784 16992
rect 22376 17051 22428 17060
rect 22376 17017 22385 17051
rect 22385 17017 22419 17051
rect 22419 17017 22428 17051
rect 22376 17008 22428 17017
rect 22928 17008 22980 17060
rect 26424 17076 26476 17128
rect 30380 17144 30432 17196
rect 29920 17119 29972 17128
rect 29920 17085 29929 17119
rect 29929 17085 29963 17119
rect 29963 17085 29972 17119
rect 29920 17076 29972 17085
rect 25688 17008 25740 17060
rect 26148 17008 26200 17060
rect 26700 17008 26752 17060
rect 29460 17008 29512 17060
rect 22836 16940 22888 16992
rect 26332 16940 26384 16992
rect 27344 16940 27396 16992
rect 5170 16838 5222 16890
rect 5234 16838 5286 16890
rect 5298 16838 5350 16890
rect 5362 16838 5414 16890
rect 5426 16838 5478 16890
rect 13611 16838 13663 16890
rect 13675 16838 13727 16890
rect 13739 16838 13791 16890
rect 13803 16838 13855 16890
rect 13867 16838 13919 16890
rect 22052 16838 22104 16890
rect 22116 16838 22168 16890
rect 22180 16838 22232 16890
rect 22244 16838 22296 16890
rect 22308 16838 22360 16890
rect 30493 16838 30545 16890
rect 30557 16838 30609 16890
rect 30621 16838 30673 16890
rect 30685 16838 30737 16890
rect 30749 16838 30801 16890
rect 18972 16736 19024 16788
rect 19340 16736 19392 16788
rect 19892 16736 19944 16788
rect 20996 16736 21048 16788
rect 21732 16779 21784 16788
rect 21732 16745 21741 16779
rect 21741 16745 21775 16779
rect 21775 16745 21784 16779
rect 21732 16736 21784 16745
rect 21824 16736 21876 16788
rect 16212 16600 16264 16652
rect 18512 16532 18564 16584
rect 19708 16600 19760 16652
rect 20904 16711 20956 16720
rect 20904 16677 20913 16711
rect 20913 16677 20947 16711
rect 20947 16677 20956 16711
rect 20904 16668 20956 16677
rect 22376 16736 22428 16788
rect 22468 16736 22520 16788
rect 23020 16736 23072 16788
rect 23204 16736 23256 16788
rect 26056 16736 26108 16788
rect 26148 16736 26200 16788
rect 26424 16736 26476 16788
rect 29368 16779 29420 16788
rect 29368 16745 29377 16779
rect 29377 16745 29411 16779
rect 29411 16745 29420 16779
rect 29368 16736 29420 16745
rect 20444 16575 20496 16584
rect 20444 16541 20453 16575
rect 20453 16541 20487 16575
rect 20487 16541 20496 16575
rect 20444 16532 20496 16541
rect 20628 16532 20680 16584
rect 22560 16600 22612 16652
rect 17684 16396 17736 16448
rect 19708 16507 19760 16516
rect 19708 16473 19717 16507
rect 19717 16473 19751 16507
rect 19751 16473 19760 16507
rect 19708 16464 19760 16473
rect 19432 16396 19484 16448
rect 19892 16439 19944 16448
rect 19892 16405 19901 16439
rect 19901 16405 19935 16439
rect 19935 16405 19944 16439
rect 19892 16396 19944 16405
rect 20168 16396 20220 16448
rect 21088 16396 21140 16448
rect 21456 16532 21508 16584
rect 21916 16464 21968 16516
rect 22836 16575 22888 16584
rect 22836 16541 22845 16575
rect 22845 16541 22879 16575
rect 22879 16541 22888 16575
rect 22836 16532 22888 16541
rect 22928 16532 22980 16584
rect 23112 16532 23164 16584
rect 23296 16575 23348 16584
rect 23296 16541 23305 16575
rect 23305 16541 23339 16575
rect 23339 16541 23348 16575
rect 23296 16532 23348 16541
rect 23664 16600 23716 16652
rect 26240 16668 26292 16720
rect 26240 16532 26292 16584
rect 26608 16575 26660 16584
rect 26608 16541 26617 16575
rect 26617 16541 26651 16575
rect 26651 16541 26660 16575
rect 26608 16532 26660 16541
rect 28264 16575 28316 16584
rect 28264 16541 28273 16575
rect 28273 16541 28307 16575
rect 28307 16541 28316 16575
rect 28264 16532 28316 16541
rect 29092 16575 29144 16584
rect 29092 16541 29101 16575
rect 29101 16541 29135 16575
rect 29135 16541 29144 16575
rect 29092 16532 29144 16541
rect 29920 16736 29972 16788
rect 30380 16736 30432 16788
rect 30932 16736 30984 16788
rect 23388 16464 23440 16516
rect 26332 16464 26384 16516
rect 30380 16575 30432 16584
rect 30380 16541 30389 16575
rect 30389 16541 30423 16575
rect 30423 16541 30432 16575
rect 30380 16532 30432 16541
rect 30656 16532 30708 16584
rect 31392 16532 31444 16584
rect 26792 16439 26844 16448
rect 26792 16405 26801 16439
rect 26801 16405 26835 16439
rect 26835 16405 26844 16439
rect 26792 16396 26844 16405
rect 28448 16439 28500 16448
rect 28448 16405 28457 16439
rect 28457 16405 28491 16439
rect 28491 16405 28500 16439
rect 28448 16396 28500 16405
rect 29184 16396 29236 16448
rect 31484 16464 31536 16516
rect 29920 16439 29972 16448
rect 29920 16405 29929 16439
rect 29929 16405 29963 16439
rect 29963 16405 29972 16439
rect 29920 16396 29972 16405
rect 30012 16396 30064 16448
rect 32220 16396 32272 16448
rect 9390 16294 9442 16346
rect 9454 16294 9506 16346
rect 9518 16294 9570 16346
rect 9582 16294 9634 16346
rect 9646 16294 9698 16346
rect 17831 16294 17883 16346
rect 17895 16294 17947 16346
rect 17959 16294 18011 16346
rect 18023 16294 18075 16346
rect 18087 16294 18139 16346
rect 26272 16294 26324 16346
rect 26336 16294 26388 16346
rect 26400 16294 26452 16346
rect 26464 16294 26516 16346
rect 26528 16294 26580 16346
rect 34713 16294 34765 16346
rect 34777 16294 34829 16346
rect 34841 16294 34893 16346
rect 34905 16294 34957 16346
rect 34969 16294 35021 16346
rect 17684 16192 17736 16244
rect 18972 16192 19024 16244
rect 19432 16192 19484 16244
rect 25228 16192 25280 16244
rect 18236 16056 18288 16108
rect 19892 16124 19944 16176
rect 18512 15988 18564 16040
rect 20628 15988 20680 16040
rect 18420 15920 18472 15972
rect 20168 15963 20220 15972
rect 20168 15929 20177 15963
rect 20177 15929 20211 15963
rect 20211 15929 20220 15963
rect 20168 15920 20220 15929
rect 25780 16099 25832 16108
rect 25780 16065 25789 16099
rect 25789 16065 25823 16099
rect 25823 16065 25832 16099
rect 25780 16056 25832 16065
rect 25964 16099 26016 16108
rect 25964 16065 25973 16099
rect 25973 16065 26007 16099
rect 26007 16065 26016 16099
rect 25964 16056 26016 16065
rect 26148 16235 26200 16244
rect 26148 16201 26157 16235
rect 26157 16201 26191 16235
rect 26191 16201 26200 16235
rect 26148 16192 26200 16201
rect 26608 16192 26660 16244
rect 26792 16192 26844 16244
rect 26976 16235 27028 16244
rect 26976 16201 26985 16235
rect 26985 16201 27019 16235
rect 27019 16201 27028 16235
rect 26976 16192 27028 16201
rect 28448 16192 28500 16244
rect 29092 16192 29144 16244
rect 29920 16192 29972 16244
rect 30380 16124 30432 16176
rect 26056 15988 26108 16040
rect 24492 15895 24544 15904
rect 24492 15861 24501 15895
rect 24501 15861 24535 15895
rect 24535 15861 24544 15895
rect 24492 15852 24544 15861
rect 24584 15852 24636 15904
rect 26240 15920 26292 15972
rect 25872 15852 25924 15904
rect 27620 16056 27672 16108
rect 28540 16056 28592 16108
rect 29736 16056 29788 16108
rect 30656 15852 30708 15904
rect 31392 15895 31444 15904
rect 31392 15861 31401 15895
rect 31401 15861 31435 15895
rect 31435 15861 31444 15895
rect 31392 15852 31444 15861
rect 5170 15750 5222 15802
rect 5234 15750 5286 15802
rect 5298 15750 5350 15802
rect 5362 15750 5414 15802
rect 5426 15750 5478 15802
rect 13611 15750 13663 15802
rect 13675 15750 13727 15802
rect 13739 15750 13791 15802
rect 13803 15750 13855 15802
rect 13867 15750 13919 15802
rect 22052 15750 22104 15802
rect 22116 15750 22168 15802
rect 22180 15750 22232 15802
rect 22244 15750 22296 15802
rect 22308 15750 22360 15802
rect 30493 15750 30545 15802
rect 30557 15750 30609 15802
rect 30621 15750 30673 15802
rect 30685 15750 30737 15802
rect 30749 15750 30801 15802
rect 24584 15648 24636 15700
rect 26056 15648 26108 15700
rect 28264 15648 28316 15700
rect 29736 15691 29788 15700
rect 29736 15657 29745 15691
rect 29745 15657 29779 15691
rect 29779 15657 29788 15691
rect 29736 15648 29788 15657
rect 30012 15691 30064 15700
rect 30012 15657 30021 15691
rect 30021 15657 30055 15691
rect 30055 15657 30064 15691
rect 30012 15648 30064 15657
rect 30380 15648 30432 15700
rect 31484 15691 31536 15700
rect 31484 15657 31493 15691
rect 31493 15657 31527 15691
rect 31527 15657 31536 15691
rect 31484 15648 31536 15657
rect 24400 15487 24452 15496
rect 24400 15453 24409 15487
rect 24409 15453 24443 15487
rect 24443 15453 24452 15487
rect 24400 15444 24452 15453
rect 24308 15376 24360 15428
rect 24676 15419 24728 15428
rect 24676 15385 24710 15419
rect 24710 15385 24728 15419
rect 24676 15376 24728 15385
rect 24860 15376 24912 15428
rect 24216 15351 24268 15360
rect 24216 15317 24225 15351
rect 24225 15317 24259 15351
rect 24259 15317 24268 15351
rect 24216 15308 24268 15317
rect 27620 15444 27672 15496
rect 28172 15487 28224 15496
rect 28172 15453 28181 15487
rect 28181 15453 28215 15487
rect 28215 15453 28224 15487
rect 28172 15444 28224 15453
rect 28908 15580 28960 15632
rect 29092 15512 29144 15564
rect 26240 15376 26292 15428
rect 26700 15376 26752 15428
rect 28908 15444 28960 15496
rect 31300 15444 31352 15496
rect 31668 15487 31720 15496
rect 31668 15453 31677 15487
rect 31677 15453 31711 15487
rect 31711 15453 31720 15487
rect 31668 15444 31720 15453
rect 29368 15376 29420 15428
rect 30564 15376 30616 15428
rect 26148 15308 26200 15360
rect 27988 15351 28040 15360
rect 27988 15317 27997 15351
rect 27997 15317 28031 15351
rect 28031 15317 28040 15351
rect 27988 15308 28040 15317
rect 9390 15206 9442 15258
rect 9454 15206 9506 15258
rect 9518 15206 9570 15258
rect 9582 15206 9634 15258
rect 9646 15206 9698 15258
rect 17831 15206 17883 15258
rect 17895 15206 17947 15258
rect 17959 15206 18011 15258
rect 18023 15206 18075 15258
rect 18087 15206 18139 15258
rect 26272 15206 26324 15258
rect 26336 15206 26388 15258
rect 26400 15206 26452 15258
rect 26464 15206 26516 15258
rect 26528 15206 26580 15258
rect 34713 15206 34765 15258
rect 34777 15206 34829 15258
rect 34841 15206 34893 15258
rect 34905 15206 34957 15258
rect 34969 15206 35021 15258
rect 20628 15104 20680 15156
rect 26608 15104 26660 15156
rect 26700 15147 26752 15156
rect 26700 15113 26709 15147
rect 26709 15113 26743 15147
rect 26743 15113 26752 15147
rect 26700 15104 26752 15113
rect 29368 15104 29420 15156
rect 30564 15104 30616 15156
rect 31392 15104 31444 15156
rect 31668 15147 31720 15156
rect 31668 15113 31677 15147
rect 31677 15113 31711 15147
rect 31711 15113 31720 15147
rect 31668 15104 31720 15113
rect 22652 15036 22704 15088
rect 20076 15011 20128 15020
rect 20076 14977 20110 15011
rect 20110 14977 20128 15011
rect 20076 14968 20128 14977
rect 23296 15011 23348 15020
rect 23296 14977 23330 15011
rect 23330 14977 23348 15011
rect 23296 14968 23348 14977
rect 24216 15036 24268 15088
rect 25964 15079 26016 15088
rect 25964 15045 25973 15079
rect 25973 15045 26007 15079
rect 26007 15045 26016 15079
rect 25964 15036 26016 15045
rect 27988 15036 28040 15088
rect 24400 14968 24452 15020
rect 26056 14968 26108 15020
rect 26240 15011 26292 15020
rect 26240 14977 26249 15011
rect 26249 14977 26283 15011
rect 26283 14977 26292 15011
rect 26240 14968 26292 14977
rect 26516 15011 26568 15020
rect 26516 14977 26525 15011
rect 26525 14977 26559 15011
rect 26559 14977 26568 15011
rect 26516 14968 26568 14977
rect 27620 15011 27672 15020
rect 27620 14977 27629 15011
rect 27629 14977 27663 15011
rect 27663 14977 27672 15011
rect 27620 14968 27672 14977
rect 31484 15011 31536 15020
rect 31484 14977 31493 15011
rect 31493 14977 31527 15011
rect 31527 14977 31536 15011
rect 31484 14968 31536 14977
rect 24308 14900 24360 14952
rect 25780 14764 25832 14816
rect 27896 14764 27948 14816
rect 5170 14662 5222 14714
rect 5234 14662 5286 14714
rect 5298 14662 5350 14714
rect 5362 14662 5414 14714
rect 5426 14662 5478 14714
rect 13611 14662 13663 14714
rect 13675 14662 13727 14714
rect 13739 14662 13791 14714
rect 13803 14662 13855 14714
rect 13867 14662 13919 14714
rect 22052 14662 22104 14714
rect 22116 14662 22168 14714
rect 22180 14662 22232 14714
rect 22244 14662 22296 14714
rect 22308 14662 22360 14714
rect 30493 14662 30545 14714
rect 30557 14662 30609 14714
rect 30621 14662 30673 14714
rect 30685 14662 30737 14714
rect 30749 14662 30801 14714
rect 23296 14560 23348 14612
rect 24676 14560 24728 14612
rect 25964 14560 26016 14612
rect 26516 14560 26568 14612
rect 28172 14560 28224 14612
rect 25412 14424 25464 14476
rect 1676 14288 1728 14340
rect 24492 14356 24544 14408
rect 25872 14356 25924 14408
rect 27896 14399 27948 14408
rect 27896 14365 27905 14399
rect 27905 14365 27939 14399
rect 27939 14365 27948 14399
rect 27896 14356 27948 14365
rect 28448 14356 28500 14408
rect 9390 14118 9442 14170
rect 9454 14118 9506 14170
rect 9518 14118 9570 14170
rect 9582 14118 9634 14170
rect 9646 14118 9698 14170
rect 17831 14118 17883 14170
rect 17895 14118 17947 14170
rect 17959 14118 18011 14170
rect 18023 14118 18075 14170
rect 18087 14118 18139 14170
rect 26272 14118 26324 14170
rect 26336 14118 26388 14170
rect 26400 14118 26452 14170
rect 26464 14118 26516 14170
rect 26528 14118 26580 14170
rect 34713 14118 34765 14170
rect 34777 14118 34829 14170
rect 34841 14118 34893 14170
rect 34905 14118 34957 14170
rect 34969 14118 35021 14170
rect 5170 13574 5222 13626
rect 5234 13574 5286 13626
rect 5298 13574 5350 13626
rect 5362 13574 5414 13626
rect 5426 13574 5478 13626
rect 13611 13574 13663 13626
rect 13675 13574 13727 13626
rect 13739 13574 13791 13626
rect 13803 13574 13855 13626
rect 13867 13574 13919 13626
rect 22052 13574 22104 13626
rect 22116 13574 22168 13626
rect 22180 13574 22232 13626
rect 22244 13574 22296 13626
rect 22308 13574 22360 13626
rect 30493 13574 30545 13626
rect 30557 13574 30609 13626
rect 30621 13574 30673 13626
rect 30685 13574 30737 13626
rect 30749 13574 30801 13626
rect 9390 13030 9442 13082
rect 9454 13030 9506 13082
rect 9518 13030 9570 13082
rect 9582 13030 9634 13082
rect 9646 13030 9698 13082
rect 17831 13030 17883 13082
rect 17895 13030 17947 13082
rect 17959 13030 18011 13082
rect 18023 13030 18075 13082
rect 18087 13030 18139 13082
rect 26272 13030 26324 13082
rect 26336 13030 26388 13082
rect 26400 13030 26452 13082
rect 26464 13030 26516 13082
rect 26528 13030 26580 13082
rect 34713 13030 34765 13082
rect 34777 13030 34829 13082
rect 34841 13030 34893 13082
rect 34905 13030 34957 13082
rect 34969 13030 35021 13082
rect 5170 12486 5222 12538
rect 5234 12486 5286 12538
rect 5298 12486 5350 12538
rect 5362 12486 5414 12538
rect 5426 12486 5478 12538
rect 13611 12486 13663 12538
rect 13675 12486 13727 12538
rect 13739 12486 13791 12538
rect 13803 12486 13855 12538
rect 13867 12486 13919 12538
rect 22052 12486 22104 12538
rect 22116 12486 22168 12538
rect 22180 12486 22232 12538
rect 22244 12486 22296 12538
rect 22308 12486 22360 12538
rect 30493 12486 30545 12538
rect 30557 12486 30609 12538
rect 30621 12486 30673 12538
rect 30685 12486 30737 12538
rect 30749 12486 30801 12538
rect 16028 12180 16080 12232
rect 34152 12087 34204 12096
rect 34152 12053 34161 12087
rect 34161 12053 34195 12087
rect 34195 12053 34204 12087
rect 34152 12044 34204 12053
rect 9390 11942 9442 11994
rect 9454 11942 9506 11994
rect 9518 11942 9570 11994
rect 9582 11942 9634 11994
rect 9646 11942 9698 11994
rect 17831 11942 17883 11994
rect 17895 11942 17947 11994
rect 17959 11942 18011 11994
rect 18023 11942 18075 11994
rect 18087 11942 18139 11994
rect 26272 11942 26324 11994
rect 26336 11942 26388 11994
rect 26400 11942 26452 11994
rect 26464 11942 26516 11994
rect 26528 11942 26580 11994
rect 34713 11942 34765 11994
rect 34777 11942 34829 11994
rect 34841 11942 34893 11994
rect 34905 11942 34957 11994
rect 34969 11942 35021 11994
rect 34152 11840 34204 11892
rect 34520 11568 34572 11620
rect 5170 11398 5222 11450
rect 5234 11398 5286 11450
rect 5298 11398 5350 11450
rect 5362 11398 5414 11450
rect 5426 11398 5478 11450
rect 13611 11398 13663 11450
rect 13675 11398 13727 11450
rect 13739 11398 13791 11450
rect 13803 11398 13855 11450
rect 13867 11398 13919 11450
rect 22052 11398 22104 11450
rect 22116 11398 22168 11450
rect 22180 11398 22232 11450
rect 22244 11398 22296 11450
rect 22308 11398 22360 11450
rect 30493 11398 30545 11450
rect 30557 11398 30609 11450
rect 30621 11398 30673 11450
rect 30685 11398 30737 11450
rect 30749 11398 30801 11450
rect 9390 10854 9442 10906
rect 9454 10854 9506 10906
rect 9518 10854 9570 10906
rect 9582 10854 9634 10906
rect 9646 10854 9698 10906
rect 17831 10854 17883 10906
rect 17895 10854 17947 10906
rect 17959 10854 18011 10906
rect 18023 10854 18075 10906
rect 18087 10854 18139 10906
rect 26272 10854 26324 10906
rect 26336 10854 26388 10906
rect 26400 10854 26452 10906
rect 26464 10854 26516 10906
rect 26528 10854 26580 10906
rect 34713 10854 34765 10906
rect 34777 10854 34829 10906
rect 34841 10854 34893 10906
rect 34905 10854 34957 10906
rect 34969 10854 35021 10906
rect 5170 10310 5222 10362
rect 5234 10310 5286 10362
rect 5298 10310 5350 10362
rect 5362 10310 5414 10362
rect 5426 10310 5478 10362
rect 13611 10310 13663 10362
rect 13675 10310 13727 10362
rect 13739 10310 13791 10362
rect 13803 10310 13855 10362
rect 13867 10310 13919 10362
rect 22052 10310 22104 10362
rect 22116 10310 22168 10362
rect 22180 10310 22232 10362
rect 22244 10310 22296 10362
rect 22308 10310 22360 10362
rect 30493 10310 30545 10362
rect 30557 10310 30609 10362
rect 30621 10310 30673 10362
rect 30685 10310 30737 10362
rect 30749 10310 30801 10362
rect 1400 10047 1452 10056
rect 1400 10013 1409 10047
rect 1409 10013 1443 10047
rect 1443 10013 1452 10047
rect 1400 10004 1452 10013
rect 9390 9766 9442 9818
rect 9454 9766 9506 9818
rect 9518 9766 9570 9818
rect 9582 9766 9634 9818
rect 9646 9766 9698 9818
rect 17831 9766 17883 9818
rect 17895 9766 17947 9818
rect 17959 9766 18011 9818
rect 18023 9766 18075 9818
rect 18087 9766 18139 9818
rect 26272 9766 26324 9818
rect 26336 9766 26388 9818
rect 26400 9766 26452 9818
rect 26464 9766 26516 9818
rect 26528 9766 26580 9818
rect 34713 9766 34765 9818
rect 34777 9766 34829 9818
rect 34841 9766 34893 9818
rect 34905 9766 34957 9818
rect 34969 9766 35021 9818
rect 5170 9222 5222 9274
rect 5234 9222 5286 9274
rect 5298 9222 5350 9274
rect 5362 9222 5414 9274
rect 5426 9222 5478 9274
rect 13611 9222 13663 9274
rect 13675 9222 13727 9274
rect 13739 9222 13791 9274
rect 13803 9222 13855 9274
rect 13867 9222 13919 9274
rect 22052 9222 22104 9274
rect 22116 9222 22168 9274
rect 22180 9222 22232 9274
rect 22244 9222 22296 9274
rect 22308 9222 22360 9274
rect 30493 9222 30545 9274
rect 30557 9222 30609 9274
rect 30621 9222 30673 9274
rect 30685 9222 30737 9274
rect 30749 9222 30801 9274
rect 9390 8678 9442 8730
rect 9454 8678 9506 8730
rect 9518 8678 9570 8730
rect 9582 8678 9634 8730
rect 9646 8678 9698 8730
rect 17831 8678 17883 8730
rect 17895 8678 17947 8730
rect 17959 8678 18011 8730
rect 18023 8678 18075 8730
rect 18087 8678 18139 8730
rect 26272 8678 26324 8730
rect 26336 8678 26388 8730
rect 26400 8678 26452 8730
rect 26464 8678 26516 8730
rect 26528 8678 26580 8730
rect 34713 8678 34765 8730
rect 34777 8678 34829 8730
rect 34841 8678 34893 8730
rect 34905 8678 34957 8730
rect 34969 8678 35021 8730
rect 5170 8134 5222 8186
rect 5234 8134 5286 8186
rect 5298 8134 5350 8186
rect 5362 8134 5414 8186
rect 5426 8134 5478 8186
rect 13611 8134 13663 8186
rect 13675 8134 13727 8186
rect 13739 8134 13791 8186
rect 13803 8134 13855 8186
rect 13867 8134 13919 8186
rect 22052 8134 22104 8186
rect 22116 8134 22168 8186
rect 22180 8134 22232 8186
rect 22244 8134 22296 8186
rect 22308 8134 22360 8186
rect 30493 8134 30545 8186
rect 30557 8134 30609 8186
rect 30621 8134 30673 8186
rect 30685 8134 30737 8186
rect 30749 8134 30801 8186
rect 9390 7590 9442 7642
rect 9454 7590 9506 7642
rect 9518 7590 9570 7642
rect 9582 7590 9634 7642
rect 9646 7590 9698 7642
rect 17831 7590 17883 7642
rect 17895 7590 17947 7642
rect 17959 7590 18011 7642
rect 18023 7590 18075 7642
rect 18087 7590 18139 7642
rect 26272 7590 26324 7642
rect 26336 7590 26388 7642
rect 26400 7590 26452 7642
rect 26464 7590 26516 7642
rect 26528 7590 26580 7642
rect 34713 7590 34765 7642
rect 34777 7590 34829 7642
rect 34841 7590 34893 7642
rect 34905 7590 34957 7642
rect 34969 7590 35021 7642
rect 5170 7046 5222 7098
rect 5234 7046 5286 7098
rect 5298 7046 5350 7098
rect 5362 7046 5414 7098
rect 5426 7046 5478 7098
rect 13611 7046 13663 7098
rect 13675 7046 13727 7098
rect 13739 7046 13791 7098
rect 13803 7046 13855 7098
rect 13867 7046 13919 7098
rect 22052 7046 22104 7098
rect 22116 7046 22168 7098
rect 22180 7046 22232 7098
rect 22244 7046 22296 7098
rect 22308 7046 22360 7098
rect 30493 7046 30545 7098
rect 30557 7046 30609 7098
rect 30621 7046 30673 7098
rect 30685 7046 30737 7098
rect 30749 7046 30801 7098
rect 9390 6502 9442 6554
rect 9454 6502 9506 6554
rect 9518 6502 9570 6554
rect 9582 6502 9634 6554
rect 9646 6502 9698 6554
rect 17831 6502 17883 6554
rect 17895 6502 17947 6554
rect 17959 6502 18011 6554
rect 18023 6502 18075 6554
rect 18087 6502 18139 6554
rect 26272 6502 26324 6554
rect 26336 6502 26388 6554
rect 26400 6502 26452 6554
rect 26464 6502 26516 6554
rect 26528 6502 26580 6554
rect 34713 6502 34765 6554
rect 34777 6502 34829 6554
rect 34841 6502 34893 6554
rect 34905 6502 34957 6554
rect 34969 6502 35021 6554
rect 5170 5958 5222 6010
rect 5234 5958 5286 6010
rect 5298 5958 5350 6010
rect 5362 5958 5414 6010
rect 5426 5958 5478 6010
rect 13611 5958 13663 6010
rect 13675 5958 13727 6010
rect 13739 5958 13791 6010
rect 13803 5958 13855 6010
rect 13867 5958 13919 6010
rect 22052 5958 22104 6010
rect 22116 5958 22168 6010
rect 22180 5958 22232 6010
rect 22244 5958 22296 6010
rect 22308 5958 22360 6010
rect 30493 5958 30545 6010
rect 30557 5958 30609 6010
rect 30621 5958 30673 6010
rect 30685 5958 30737 6010
rect 30749 5958 30801 6010
rect 9390 5414 9442 5466
rect 9454 5414 9506 5466
rect 9518 5414 9570 5466
rect 9582 5414 9634 5466
rect 9646 5414 9698 5466
rect 17831 5414 17883 5466
rect 17895 5414 17947 5466
rect 17959 5414 18011 5466
rect 18023 5414 18075 5466
rect 18087 5414 18139 5466
rect 26272 5414 26324 5466
rect 26336 5414 26388 5466
rect 26400 5414 26452 5466
rect 26464 5414 26516 5466
rect 26528 5414 26580 5466
rect 34713 5414 34765 5466
rect 34777 5414 34829 5466
rect 34841 5414 34893 5466
rect 34905 5414 34957 5466
rect 34969 5414 35021 5466
rect 5170 4870 5222 4922
rect 5234 4870 5286 4922
rect 5298 4870 5350 4922
rect 5362 4870 5414 4922
rect 5426 4870 5478 4922
rect 13611 4870 13663 4922
rect 13675 4870 13727 4922
rect 13739 4870 13791 4922
rect 13803 4870 13855 4922
rect 13867 4870 13919 4922
rect 22052 4870 22104 4922
rect 22116 4870 22168 4922
rect 22180 4870 22232 4922
rect 22244 4870 22296 4922
rect 22308 4870 22360 4922
rect 30493 4870 30545 4922
rect 30557 4870 30609 4922
rect 30621 4870 30673 4922
rect 30685 4870 30737 4922
rect 30749 4870 30801 4922
rect 9390 4326 9442 4378
rect 9454 4326 9506 4378
rect 9518 4326 9570 4378
rect 9582 4326 9634 4378
rect 9646 4326 9698 4378
rect 17831 4326 17883 4378
rect 17895 4326 17947 4378
rect 17959 4326 18011 4378
rect 18023 4326 18075 4378
rect 18087 4326 18139 4378
rect 26272 4326 26324 4378
rect 26336 4326 26388 4378
rect 26400 4326 26452 4378
rect 26464 4326 26516 4378
rect 26528 4326 26580 4378
rect 34713 4326 34765 4378
rect 34777 4326 34829 4378
rect 34841 4326 34893 4378
rect 34905 4326 34957 4378
rect 34969 4326 35021 4378
rect 5170 3782 5222 3834
rect 5234 3782 5286 3834
rect 5298 3782 5350 3834
rect 5362 3782 5414 3834
rect 5426 3782 5478 3834
rect 13611 3782 13663 3834
rect 13675 3782 13727 3834
rect 13739 3782 13791 3834
rect 13803 3782 13855 3834
rect 13867 3782 13919 3834
rect 22052 3782 22104 3834
rect 22116 3782 22168 3834
rect 22180 3782 22232 3834
rect 22244 3782 22296 3834
rect 22308 3782 22360 3834
rect 30493 3782 30545 3834
rect 30557 3782 30609 3834
rect 30621 3782 30673 3834
rect 30685 3782 30737 3834
rect 30749 3782 30801 3834
rect 9390 3238 9442 3290
rect 9454 3238 9506 3290
rect 9518 3238 9570 3290
rect 9582 3238 9634 3290
rect 9646 3238 9698 3290
rect 17831 3238 17883 3290
rect 17895 3238 17947 3290
rect 17959 3238 18011 3290
rect 18023 3238 18075 3290
rect 18087 3238 18139 3290
rect 26272 3238 26324 3290
rect 26336 3238 26388 3290
rect 26400 3238 26452 3290
rect 26464 3238 26516 3290
rect 26528 3238 26580 3290
rect 34713 3238 34765 3290
rect 34777 3238 34829 3290
rect 34841 3238 34893 3290
rect 34905 3238 34957 3290
rect 34969 3238 35021 3290
rect 5170 2694 5222 2746
rect 5234 2694 5286 2746
rect 5298 2694 5350 2746
rect 5362 2694 5414 2746
rect 5426 2694 5478 2746
rect 13611 2694 13663 2746
rect 13675 2694 13727 2746
rect 13739 2694 13791 2746
rect 13803 2694 13855 2746
rect 13867 2694 13919 2746
rect 22052 2694 22104 2746
rect 22116 2694 22168 2746
rect 22180 2694 22232 2746
rect 22244 2694 22296 2746
rect 22308 2694 22360 2746
rect 30493 2694 30545 2746
rect 30557 2694 30609 2746
rect 30621 2694 30673 2746
rect 30685 2694 30737 2746
rect 30749 2694 30801 2746
rect 28448 2635 28500 2644
rect 28448 2601 28457 2635
rect 28457 2601 28491 2635
rect 28491 2601 28500 2635
rect 28448 2592 28500 2601
rect 31484 2592 31536 2644
rect 1676 2499 1728 2508
rect 1676 2465 1685 2499
rect 1685 2465 1719 2499
rect 1719 2465 1728 2499
rect 1676 2456 1728 2465
rect 20 2388 72 2440
rect 9128 2431 9180 2440
rect 9128 2397 9137 2431
rect 9137 2397 9171 2431
rect 9171 2397 9180 2431
rect 9128 2388 9180 2397
rect 19616 2431 19668 2440
rect 19616 2397 19625 2431
rect 19625 2397 19659 2431
rect 19659 2397 19668 2431
rect 19616 2388 19668 2397
rect 28356 2388 28408 2440
rect 18788 2252 18840 2304
rect 35164 2252 35216 2304
rect 9390 2150 9442 2202
rect 9454 2150 9506 2202
rect 9518 2150 9570 2202
rect 9582 2150 9634 2202
rect 9646 2150 9698 2202
rect 17831 2150 17883 2202
rect 17895 2150 17947 2202
rect 17959 2150 18011 2202
rect 18023 2150 18075 2202
rect 18087 2150 18139 2202
rect 26272 2150 26324 2202
rect 26336 2150 26388 2202
rect 26400 2150 26452 2202
rect 26464 2150 26516 2202
rect 26528 2150 26580 2202
rect 34713 2150 34765 2202
rect 34777 2150 34829 2202
rect 34841 2150 34893 2202
rect 34905 2150 34957 2202
rect 34969 2150 35021 2202
<< metal2 >>
rect 7074 41200 7186 42000
rect 16734 41200 16846 42000
rect 26394 41200 26506 42000
rect 35410 41200 35522 42000
rect 5170 39740 5478 39749
rect 5170 39738 5176 39740
rect 5232 39738 5256 39740
rect 5312 39738 5336 39740
rect 5392 39738 5416 39740
rect 5472 39738 5478 39740
rect 5232 39686 5234 39738
rect 5414 39686 5416 39738
rect 5170 39684 5176 39686
rect 5232 39684 5256 39686
rect 5312 39684 5336 39686
rect 5392 39684 5416 39686
rect 5472 39684 5478 39686
rect 5170 39675 5478 39684
rect 938 39536 994 39545
rect 938 39471 994 39480
rect 952 39438 980 39471
rect 7116 39438 7144 41200
rect 13611 39740 13919 39749
rect 13611 39738 13617 39740
rect 13673 39738 13697 39740
rect 13753 39738 13777 39740
rect 13833 39738 13857 39740
rect 13913 39738 13919 39740
rect 13673 39686 13675 39738
rect 13855 39686 13857 39738
rect 13611 39684 13617 39686
rect 13673 39684 13697 39686
rect 13753 39684 13777 39686
rect 13833 39684 13857 39686
rect 13913 39684 13919 39686
rect 13611 39675 13919 39684
rect 16776 39438 16804 41200
rect 22052 39740 22360 39749
rect 22052 39738 22058 39740
rect 22114 39738 22138 39740
rect 22194 39738 22218 39740
rect 22274 39738 22298 39740
rect 22354 39738 22360 39740
rect 22114 39686 22116 39738
rect 22296 39686 22298 39738
rect 22052 39684 22058 39686
rect 22114 39684 22138 39686
rect 22194 39684 22218 39686
rect 22274 39684 22298 39686
rect 22354 39684 22360 39686
rect 22052 39675 22360 39684
rect 26436 39642 26464 41200
rect 30493 39740 30801 39749
rect 30493 39738 30499 39740
rect 30555 39738 30579 39740
rect 30635 39738 30659 39740
rect 30715 39738 30739 39740
rect 30795 39738 30801 39740
rect 30555 39686 30557 39738
rect 30737 39686 30739 39738
rect 30493 39684 30499 39686
rect 30555 39684 30579 39686
rect 30635 39684 30659 39686
rect 30715 39684 30739 39686
rect 30795 39684 30801 39686
rect 30493 39675 30801 39684
rect 35452 39642 35480 41200
rect 26424 39636 26476 39642
rect 26424 39578 26476 39584
rect 35440 39636 35492 39642
rect 35440 39578 35492 39584
rect 940 39432 992 39438
rect 940 39374 992 39380
rect 7104 39432 7156 39438
rect 7104 39374 7156 39380
rect 16764 39432 16816 39438
rect 16764 39374 16816 39380
rect 34152 39364 34204 39370
rect 34152 39306 34204 39312
rect 1584 39296 1636 39302
rect 1584 39238 1636 39244
rect 16120 39296 16172 39302
rect 16120 39238 16172 39244
rect 17592 39296 17644 39302
rect 17592 39238 17644 39244
rect 1596 33522 1624 39238
rect 9390 39196 9698 39205
rect 9390 39194 9396 39196
rect 9452 39194 9476 39196
rect 9532 39194 9556 39196
rect 9612 39194 9636 39196
rect 9692 39194 9698 39196
rect 9452 39142 9454 39194
rect 9634 39142 9636 39194
rect 9390 39140 9396 39142
rect 9452 39140 9476 39142
rect 9532 39140 9556 39142
rect 9612 39140 9636 39142
rect 9692 39140 9698 39142
rect 9390 39131 9698 39140
rect 5170 38652 5478 38661
rect 5170 38650 5176 38652
rect 5232 38650 5256 38652
rect 5312 38650 5336 38652
rect 5392 38650 5416 38652
rect 5472 38650 5478 38652
rect 5232 38598 5234 38650
rect 5414 38598 5416 38650
rect 5170 38596 5176 38598
rect 5232 38596 5256 38598
rect 5312 38596 5336 38598
rect 5392 38596 5416 38598
rect 5472 38596 5478 38598
rect 5170 38587 5478 38596
rect 13611 38652 13919 38661
rect 13611 38650 13617 38652
rect 13673 38650 13697 38652
rect 13753 38650 13777 38652
rect 13833 38650 13857 38652
rect 13913 38650 13919 38652
rect 13673 38598 13675 38650
rect 13855 38598 13857 38650
rect 13611 38596 13617 38598
rect 13673 38596 13697 38598
rect 13753 38596 13777 38598
rect 13833 38596 13857 38598
rect 13913 38596 13919 38598
rect 13611 38587 13919 38596
rect 9390 38108 9698 38117
rect 9390 38106 9396 38108
rect 9452 38106 9476 38108
rect 9532 38106 9556 38108
rect 9612 38106 9636 38108
rect 9692 38106 9698 38108
rect 9452 38054 9454 38106
rect 9634 38054 9636 38106
rect 9390 38052 9396 38054
rect 9452 38052 9476 38054
rect 9532 38052 9556 38054
rect 9612 38052 9636 38054
rect 9692 38052 9698 38054
rect 9390 38043 9698 38052
rect 5170 37564 5478 37573
rect 5170 37562 5176 37564
rect 5232 37562 5256 37564
rect 5312 37562 5336 37564
rect 5392 37562 5416 37564
rect 5472 37562 5478 37564
rect 5232 37510 5234 37562
rect 5414 37510 5416 37562
rect 5170 37508 5176 37510
rect 5232 37508 5256 37510
rect 5312 37508 5336 37510
rect 5392 37508 5416 37510
rect 5472 37508 5478 37510
rect 5170 37499 5478 37508
rect 13611 37564 13919 37573
rect 13611 37562 13617 37564
rect 13673 37562 13697 37564
rect 13753 37562 13777 37564
rect 13833 37562 13857 37564
rect 13913 37562 13919 37564
rect 13673 37510 13675 37562
rect 13855 37510 13857 37562
rect 13611 37508 13617 37510
rect 13673 37508 13697 37510
rect 13753 37508 13777 37510
rect 13833 37508 13857 37510
rect 13913 37508 13919 37510
rect 13611 37499 13919 37508
rect 9390 37020 9698 37029
rect 9390 37018 9396 37020
rect 9452 37018 9476 37020
rect 9532 37018 9556 37020
rect 9612 37018 9636 37020
rect 9692 37018 9698 37020
rect 9452 36966 9454 37018
rect 9634 36966 9636 37018
rect 9390 36964 9396 36966
rect 9452 36964 9476 36966
rect 9532 36964 9556 36966
rect 9612 36964 9636 36966
rect 9692 36964 9698 36966
rect 9390 36955 9698 36964
rect 5170 36476 5478 36485
rect 5170 36474 5176 36476
rect 5232 36474 5256 36476
rect 5312 36474 5336 36476
rect 5392 36474 5416 36476
rect 5472 36474 5478 36476
rect 5232 36422 5234 36474
rect 5414 36422 5416 36474
rect 5170 36420 5176 36422
rect 5232 36420 5256 36422
rect 5312 36420 5336 36422
rect 5392 36420 5416 36422
rect 5472 36420 5478 36422
rect 5170 36411 5478 36420
rect 13611 36476 13919 36485
rect 13611 36474 13617 36476
rect 13673 36474 13697 36476
rect 13753 36474 13777 36476
rect 13833 36474 13857 36476
rect 13913 36474 13919 36476
rect 13673 36422 13675 36474
rect 13855 36422 13857 36474
rect 13611 36420 13617 36422
rect 13673 36420 13697 36422
rect 13753 36420 13777 36422
rect 13833 36420 13857 36422
rect 13913 36420 13919 36422
rect 13611 36411 13919 36420
rect 9390 35932 9698 35941
rect 9390 35930 9396 35932
rect 9452 35930 9476 35932
rect 9532 35930 9556 35932
rect 9612 35930 9636 35932
rect 9692 35930 9698 35932
rect 9452 35878 9454 35930
rect 9634 35878 9636 35930
rect 9390 35876 9396 35878
rect 9452 35876 9476 35878
rect 9532 35876 9556 35878
rect 9612 35876 9636 35878
rect 9692 35876 9698 35878
rect 9390 35867 9698 35876
rect 5170 35388 5478 35397
rect 5170 35386 5176 35388
rect 5232 35386 5256 35388
rect 5312 35386 5336 35388
rect 5392 35386 5416 35388
rect 5472 35386 5478 35388
rect 5232 35334 5234 35386
rect 5414 35334 5416 35386
rect 5170 35332 5176 35334
rect 5232 35332 5256 35334
rect 5312 35332 5336 35334
rect 5392 35332 5416 35334
rect 5472 35332 5478 35334
rect 5170 35323 5478 35332
rect 13611 35388 13919 35397
rect 13611 35386 13617 35388
rect 13673 35386 13697 35388
rect 13753 35386 13777 35388
rect 13833 35386 13857 35388
rect 13913 35386 13919 35388
rect 13673 35334 13675 35386
rect 13855 35334 13857 35386
rect 13611 35332 13617 35334
rect 13673 35332 13697 35334
rect 13753 35332 13777 35334
rect 13833 35332 13857 35334
rect 13913 35332 13919 35334
rect 13611 35323 13919 35332
rect 9390 34844 9698 34853
rect 9390 34842 9396 34844
rect 9452 34842 9476 34844
rect 9532 34842 9556 34844
rect 9612 34842 9636 34844
rect 9692 34842 9698 34844
rect 9452 34790 9454 34842
rect 9634 34790 9636 34842
rect 9390 34788 9396 34790
rect 9452 34788 9476 34790
rect 9532 34788 9556 34790
rect 9612 34788 9636 34790
rect 9692 34788 9698 34790
rect 9390 34779 9698 34788
rect 5170 34300 5478 34309
rect 5170 34298 5176 34300
rect 5232 34298 5256 34300
rect 5312 34298 5336 34300
rect 5392 34298 5416 34300
rect 5472 34298 5478 34300
rect 5232 34246 5234 34298
rect 5414 34246 5416 34298
rect 5170 34244 5176 34246
rect 5232 34244 5256 34246
rect 5312 34244 5336 34246
rect 5392 34244 5416 34246
rect 5472 34244 5478 34246
rect 5170 34235 5478 34244
rect 13611 34300 13919 34309
rect 13611 34298 13617 34300
rect 13673 34298 13697 34300
rect 13753 34298 13777 34300
rect 13833 34298 13857 34300
rect 13913 34298 13919 34300
rect 13673 34246 13675 34298
rect 13855 34246 13857 34298
rect 13611 34244 13617 34246
rect 13673 34244 13697 34246
rect 13753 34244 13777 34246
rect 13833 34244 13857 34246
rect 13913 34244 13919 34246
rect 13611 34235 13919 34244
rect 9390 33756 9698 33765
rect 9390 33754 9396 33756
rect 9452 33754 9476 33756
rect 9532 33754 9556 33756
rect 9612 33754 9636 33756
rect 9692 33754 9698 33756
rect 9452 33702 9454 33754
rect 9634 33702 9636 33754
rect 9390 33700 9396 33702
rect 9452 33700 9476 33702
rect 9532 33700 9556 33702
rect 9612 33700 9636 33702
rect 9692 33700 9698 33702
rect 9390 33691 9698 33700
rect 1584 33516 1636 33522
rect 1584 33458 1636 33464
rect 5170 33212 5478 33221
rect 5170 33210 5176 33212
rect 5232 33210 5256 33212
rect 5312 33210 5336 33212
rect 5392 33210 5416 33212
rect 5472 33210 5478 33212
rect 5232 33158 5234 33210
rect 5414 33158 5416 33210
rect 5170 33156 5176 33158
rect 5232 33156 5256 33158
rect 5312 33156 5336 33158
rect 5392 33156 5416 33158
rect 5472 33156 5478 33158
rect 5170 33147 5478 33156
rect 13611 33212 13919 33221
rect 13611 33210 13617 33212
rect 13673 33210 13697 33212
rect 13753 33210 13777 33212
rect 13833 33210 13857 33212
rect 13913 33210 13919 33212
rect 13673 33158 13675 33210
rect 13855 33158 13857 33210
rect 13611 33156 13617 33158
rect 13673 33156 13697 33158
rect 13753 33156 13777 33158
rect 13833 33156 13857 33158
rect 13913 33156 13919 33158
rect 13611 33147 13919 33156
rect 9390 32668 9698 32677
rect 9390 32666 9396 32668
rect 9452 32666 9476 32668
rect 9532 32666 9556 32668
rect 9612 32666 9636 32668
rect 9692 32666 9698 32668
rect 9452 32614 9454 32666
rect 9634 32614 9636 32666
rect 9390 32612 9396 32614
rect 9452 32612 9476 32614
rect 9532 32612 9556 32614
rect 9612 32612 9636 32614
rect 9692 32612 9698 32614
rect 9390 32603 9698 32612
rect 5170 32124 5478 32133
rect 5170 32122 5176 32124
rect 5232 32122 5256 32124
rect 5312 32122 5336 32124
rect 5392 32122 5416 32124
rect 5472 32122 5478 32124
rect 5232 32070 5234 32122
rect 5414 32070 5416 32122
rect 5170 32068 5176 32070
rect 5232 32068 5256 32070
rect 5312 32068 5336 32070
rect 5392 32068 5416 32070
rect 5472 32068 5478 32070
rect 5170 32059 5478 32068
rect 13611 32124 13919 32133
rect 13611 32122 13617 32124
rect 13673 32122 13697 32124
rect 13753 32122 13777 32124
rect 13833 32122 13857 32124
rect 13913 32122 13919 32124
rect 13673 32070 13675 32122
rect 13855 32070 13857 32122
rect 13611 32068 13617 32070
rect 13673 32068 13697 32070
rect 13753 32068 13777 32070
rect 13833 32068 13857 32070
rect 13913 32068 13919 32070
rect 13611 32059 13919 32068
rect 9390 31580 9698 31589
rect 9390 31578 9396 31580
rect 9452 31578 9476 31580
rect 9532 31578 9556 31580
rect 9612 31578 9636 31580
rect 9692 31578 9698 31580
rect 9452 31526 9454 31578
rect 9634 31526 9636 31578
rect 9390 31524 9396 31526
rect 9452 31524 9476 31526
rect 9532 31524 9556 31526
rect 9612 31524 9636 31526
rect 9692 31524 9698 31526
rect 9390 31515 9698 31524
rect 5170 31036 5478 31045
rect 5170 31034 5176 31036
rect 5232 31034 5256 31036
rect 5312 31034 5336 31036
rect 5392 31034 5416 31036
rect 5472 31034 5478 31036
rect 5232 30982 5234 31034
rect 5414 30982 5416 31034
rect 5170 30980 5176 30982
rect 5232 30980 5256 30982
rect 5312 30980 5336 30982
rect 5392 30980 5416 30982
rect 5472 30980 5478 30982
rect 5170 30971 5478 30980
rect 13611 31036 13919 31045
rect 13611 31034 13617 31036
rect 13673 31034 13697 31036
rect 13753 31034 13777 31036
rect 13833 31034 13857 31036
rect 13913 31034 13919 31036
rect 13673 30982 13675 31034
rect 13855 30982 13857 31034
rect 13611 30980 13617 30982
rect 13673 30980 13697 30982
rect 13753 30980 13777 30982
rect 13833 30980 13857 30982
rect 13913 30980 13919 30982
rect 13611 30971 13919 30980
rect 9390 30492 9698 30501
rect 9390 30490 9396 30492
rect 9452 30490 9476 30492
rect 9532 30490 9556 30492
rect 9612 30490 9636 30492
rect 9692 30490 9698 30492
rect 9452 30438 9454 30490
rect 9634 30438 9636 30490
rect 9390 30436 9396 30438
rect 9452 30436 9476 30438
rect 9532 30436 9556 30438
rect 9612 30436 9636 30438
rect 9692 30436 9698 30438
rect 9390 30427 9698 30436
rect 940 30048 992 30054
rect 938 30016 940 30025
rect 992 30016 994 30025
rect 938 29951 994 29960
rect 5170 29948 5478 29957
rect 5170 29946 5176 29948
rect 5232 29946 5256 29948
rect 5312 29946 5336 29948
rect 5392 29946 5416 29948
rect 5472 29946 5478 29948
rect 5232 29894 5234 29946
rect 5414 29894 5416 29946
rect 5170 29892 5176 29894
rect 5232 29892 5256 29894
rect 5312 29892 5336 29894
rect 5392 29892 5416 29894
rect 5472 29892 5478 29894
rect 5170 29883 5478 29892
rect 13611 29948 13919 29957
rect 13611 29946 13617 29948
rect 13673 29946 13697 29948
rect 13753 29946 13777 29948
rect 13833 29946 13857 29948
rect 13913 29946 13919 29948
rect 13673 29894 13675 29946
rect 13855 29894 13857 29946
rect 13611 29892 13617 29894
rect 13673 29892 13697 29894
rect 13753 29892 13777 29894
rect 13833 29892 13857 29894
rect 13913 29892 13919 29894
rect 13611 29883 13919 29892
rect 9390 29404 9698 29413
rect 9390 29402 9396 29404
rect 9452 29402 9476 29404
rect 9532 29402 9556 29404
rect 9612 29402 9636 29404
rect 9692 29402 9698 29404
rect 9452 29350 9454 29402
rect 9634 29350 9636 29402
rect 9390 29348 9396 29350
rect 9452 29348 9476 29350
rect 9532 29348 9556 29350
rect 9612 29348 9636 29350
rect 9692 29348 9698 29350
rect 9390 29339 9698 29348
rect 5170 28860 5478 28869
rect 5170 28858 5176 28860
rect 5232 28858 5256 28860
rect 5312 28858 5336 28860
rect 5392 28858 5416 28860
rect 5472 28858 5478 28860
rect 5232 28806 5234 28858
rect 5414 28806 5416 28858
rect 5170 28804 5176 28806
rect 5232 28804 5256 28806
rect 5312 28804 5336 28806
rect 5392 28804 5416 28806
rect 5472 28804 5478 28806
rect 5170 28795 5478 28804
rect 13611 28860 13919 28869
rect 13611 28858 13617 28860
rect 13673 28858 13697 28860
rect 13753 28858 13777 28860
rect 13833 28858 13857 28860
rect 13913 28858 13919 28860
rect 13673 28806 13675 28858
rect 13855 28806 13857 28858
rect 13611 28804 13617 28806
rect 13673 28804 13697 28806
rect 13753 28804 13777 28806
rect 13833 28804 13857 28806
rect 13913 28804 13919 28806
rect 13611 28795 13919 28804
rect 9390 28316 9698 28325
rect 9390 28314 9396 28316
rect 9452 28314 9476 28316
rect 9532 28314 9556 28316
rect 9612 28314 9636 28316
rect 9692 28314 9698 28316
rect 9452 28262 9454 28314
rect 9634 28262 9636 28314
rect 9390 28260 9396 28262
rect 9452 28260 9476 28262
rect 9532 28260 9556 28262
rect 9612 28260 9636 28262
rect 9692 28260 9698 28262
rect 9390 28251 9698 28260
rect 5170 27772 5478 27781
rect 5170 27770 5176 27772
rect 5232 27770 5256 27772
rect 5312 27770 5336 27772
rect 5392 27770 5416 27772
rect 5472 27770 5478 27772
rect 5232 27718 5234 27770
rect 5414 27718 5416 27770
rect 5170 27716 5176 27718
rect 5232 27716 5256 27718
rect 5312 27716 5336 27718
rect 5392 27716 5416 27718
rect 5472 27716 5478 27718
rect 5170 27707 5478 27716
rect 13611 27772 13919 27781
rect 13611 27770 13617 27772
rect 13673 27770 13697 27772
rect 13753 27770 13777 27772
rect 13833 27770 13857 27772
rect 13913 27770 13919 27772
rect 13673 27718 13675 27770
rect 13855 27718 13857 27770
rect 13611 27716 13617 27718
rect 13673 27716 13697 27718
rect 13753 27716 13777 27718
rect 13833 27716 13857 27718
rect 13913 27716 13919 27718
rect 13611 27707 13919 27716
rect 9390 27228 9698 27237
rect 9390 27226 9396 27228
rect 9452 27226 9476 27228
rect 9532 27226 9556 27228
rect 9612 27226 9636 27228
rect 9692 27226 9698 27228
rect 9452 27174 9454 27226
rect 9634 27174 9636 27226
rect 9390 27172 9396 27174
rect 9452 27172 9476 27174
rect 9532 27172 9556 27174
rect 9612 27172 9636 27174
rect 9692 27172 9698 27174
rect 9390 27163 9698 27172
rect 5170 26684 5478 26693
rect 5170 26682 5176 26684
rect 5232 26682 5256 26684
rect 5312 26682 5336 26684
rect 5392 26682 5416 26684
rect 5472 26682 5478 26684
rect 5232 26630 5234 26682
rect 5414 26630 5416 26682
rect 5170 26628 5176 26630
rect 5232 26628 5256 26630
rect 5312 26628 5336 26630
rect 5392 26628 5416 26630
rect 5472 26628 5478 26630
rect 5170 26619 5478 26628
rect 13611 26684 13919 26693
rect 13611 26682 13617 26684
rect 13673 26682 13697 26684
rect 13753 26682 13777 26684
rect 13833 26682 13857 26684
rect 13913 26682 13919 26684
rect 13673 26630 13675 26682
rect 13855 26630 13857 26682
rect 13611 26628 13617 26630
rect 13673 26628 13697 26630
rect 13753 26628 13777 26630
rect 13833 26628 13857 26630
rect 13913 26628 13919 26630
rect 13611 26619 13919 26628
rect 9390 26140 9698 26149
rect 9390 26138 9396 26140
rect 9452 26138 9476 26140
rect 9532 26138 9556 26140
rect 9612 26138 9636 26140
rect 9692 26138 9698 26140
rect 9452 26086 9454 26138
rect 9634 26086 9636 26138
rect 9390 26084 9396 26086
rect 9452 26084 9476 26086
rect 9532 26084 9556 26086
rect 9612 26084 9636 26086
rect 9692 26084 9698 26086
rect 9390 26075 9698 26084
rect 5170 25596 5478 25605
rect 5170 25594 5176 25596
rect 5232 25594 5256 25596
rect 5312 25594 5336 25596
rect 5392 25594 5416 25596
rect 5472 25594 5478 25596
rect 5232 25542 5234 25594
rect 5414 25542 5416 25594
rect 5170 25540 5176 25542
rect 5232 25540 5256 25542
rect 5312 25540 5336 25542
rect 5392 25540 5416 25542
rect 5472 25540 5478 25542
rect 5170 25531 5478 25540
rect 13611 25596 13919 25605
rect 13611 25594 13617 25596
rect 13673 25594 13697 25596
rect 13753 25594 13777 25596
rect 13833 25594 13857 25596
rect 13913 25594 13919 25596
rect 13673 25542 13675 25594
rect 13855 25542 13857 25594
rect 13611 25540 13617 25542
rect 13673 25540 13697 25542
rect 13753 25540 13777 25542
rect 13833 25540 13857 25542
rect 13913 25540 13919 25542
rect 13611 25531 13919 25540
rect 9390 25052 9698 25061
rect 9390 25050 9396 25052
rect 9452 25050 9476 25052
rect 9532 25050 9556 25052
rect 9612 25050 9636 25052
rect 9692 25050 9698 25052
rect 9452 24998 9454 25050
rect 9634 24998 9636 25050
rect 9390 24996 9396 24998
rect 9452 24996 9476 24998
rect 9532 24996 9556 24998
rect 9612 24996 9636 24998
rect 9692 24996 9698 24998
rect 9390 24987 9698 24996
rect 5170 24508 5478 24517
rect 5170 24506 5176 24508
rect 5232 24506 5256 24508
rect 5312 24506 5336 24508
rect 5392 24506 5416 24508
rect 5472 24506 5478 24508
rect 5232 24454 5234 24506
rect 5414 24454 5416 24506
rect 5170 24452 5176 24454
rect 5232 24452 5256 24454
rect 5312 24452 5336 24454
rect 5392 24452 5416 24454
rect 5472 24452 5478 24454
rect 5170 24443 5478 24452
rect 13611 24508 13919 24517
rect 13611 24506 13617 24508
rect 13673 24506 13697 24508
rect 13753 24506 13777 24508
rect 13833 24506 13857 24508
rect 13913 24506 13919 24508
rect 13673 24454 13675 24506
rect 13855 24454 13857 24506
rect 13611 24452 13617 24454
rect 13673 24452 13697 24454
rect 13753 24452 13777 24454
rect 13833 24452 13857 24454
rect 13913 24452 13919 24454
rect 13611 24443 13919 24452
rect 9390 23964 9698 23973
rect 9390 23962 9396 23964
rect 9452 23962 9476 23964
rect 9532 23962 9556 23964
rect 9612 23962 9636 23964
rect 9692 23962 9698 23964
rect 9452 23910 9454 23962
rect 9634 23910 9636 23962
rect 9390 23908 9396 23910
rect 9452 23908 9476 23910
rect 9532 23908 9556 23910
rect 9612 23908 9636 23910
rect 9692 23908 9698 23910
rect 9390 23899 9698 23908
rect 5170 23420 5478 23429
rect 5170 23418 5176 23420
rect 5232 23418 5256 23420
rect 5312 23418 5336 23420
rect 5392 23418 5416 23420
rect 5472 23418 5478 23420
rect 5232 23366 5234 23418
rect 5414 23366 5416 23418
rect 5170 23364 5176 23366
rect 5232 23364 5256 23366
rect 5312 23364 5336 23366
rect 5392 23364 5416 23366
rect 5472 23364 5478 23366
rect 5170 23355 5478 23364
rect 13611 23420 13919 23429
rect 13611 23418 13617 23420
rect 13673 23418 13697 23420
rect 13753 23418 13777 23420
rect 13833 23418 13857 23420
rect 13913 23418 13919 23420
rect 13673 23366 13675 23418
rect 13855 23366 13857 23418
rect 13611 23364 13617 23366
rect 13673 23364 13697 23366
rect 13753 23364 13777 23366
rect 13833 23364 13857 23366
rect 13913 23364 13919 23366
rect 13611 23355 13919 23364
rect 9390 22876 9698 22885
rect 9390 22874 9396 22876
rect 9452 22874 9476 22876
rect 9532 22874 9556 22876
rect 9612 22874 9636 22876
rect 9692 22874 9698 22876
rect 9452 22822 9454 22874
rect 9634 22822 9636 22874
rect 9390 22820 9396 22822
rect 9452 22820 9476 22822
rect 9532 22820 9556 22822
rect 9612 22820 9636 22822
rect 9692 22820 9698 22822
rect 9390 22811 9698 22820
rect 5170 22332 5478 22341
rect 5170 22330 5176 22332
rect 5232 22330 5256 22332
rect 5312 22330 5336 22332
rect 5392 22330 5416 22332
rect 5472 22330 5478 22332
rect 5232 22278 5234 22330
rect 5414 22278 5416 22330
rect 5170 22276 5176 22278
rect 5232 22276 5256 22278
rect 5312 22276 5336 22278
rect 5392 22276 5416 22278
rect 5472 22276 5478 22278
rect 5170 22267 5478 22276
rect 13611 22332 13919 22341
rect 13611 22330 13617 22332
rect 13673 22330 13697 22332
rect 13753 22330 13777 22332
rect 13833 22330 13857 22332
rect 13913 22330 13919 22332
rect 13673 22278 13675 22330
rect 13855 22278 13857 22330
rect 13611 22276 13617 22278
rect 13673 22276 13697 22278
rect 13753 22276 13777 22278
rect 13833 22276 13857 22278
rect 13913 22276 13919 22278
rect 13611 22267 13919 22276
rect 16132 22094 16160 39238
rect 17132 32292 17184 32298
rect 17132 32234 17184 32240
rect 17144 31822 17172 32234
rect 17316 32224 17368 32230
rect 17316 32166 17368 32172
rect 17328 31822 17356 32166
rect 16672 31816 16724 31822
rect 16672 31758 16724 31764
rect 17132 31816 17184 31822
rect 17132 31758 17184 31764
rect 17316 31816 17368 31822
rect 17316 31758 17368 31764
rect 16684 31686 16712 31758
rect 16672 31680 16724 31686
rect 16672 31622 16724 31628
rect 16684 31278 16712 31622
rect 16764 31340 16816 31346
rect 16764 31282 16816 31288
rect 16672 31272 16724 31278
rect 16672 31214 16724 31220
rect 16684 30190 16712 31214
rect 16776 30938 16804 31282
rect 17604 31090 17632 39238
rect 17831 39196 18139 39205
rect 17831 39194 17837 39196
rect 17893 39194 17917 39196
rect 17973 39194 17997 39196
rect 18053 39194 18077 39196
rect 18133 39194 18139 39196
rect 17893 39142 17895 39194
rect 18075 39142 18077 39194
rect 17831 39140 17837 39142
rect 17893 39140 17917 39142
rect 17973 39140 17997 39142
rect 18053 39140 18077 39142
rect 18133 39140 18139 39142
rect 17831 39131 18139 39140
rect 26272 39196 26580 39205
rect 26272 39194 26278 39196
rect 26334 39194 26358 39196
rect 26414 39194 26438 39196
rect 26494 39194 26518 39196
rect 26574 39194 26580 39196
rect 26334 39142 26336 39194
rect 26516 39142 26518 39194
rect 26272 39140 26278 39142
rect 26334 39140 26358 39142
rect 26414 39140 26438 39142
rect 26494 39140 26518 39142
rect 26574 39140 26580 39142
rect 26272 39131 26580 39140
rect 22052 38652 22360 38661
rect 22052 38650 22058 38652
rect 22114 38650 22138 38652
rect 22194 38650 22218 38652
rect 22274 38650 22298 38652
rect 22354 38650 22360 38652
rect 22114 38598 22116 38650
rect 22296 38598 22298 38650
rect 22052 38596 22058 38598
rect 22114 38596 22138 38598
rect 22194 38596 22218 38598
rect 22274 38596 22298 38598
rect 22354 38596 22360 38598
rect 22052 38587 22360 38596
rect 30493 38652 30801 38661
rect 30493 38650 30499 38652
rect 30555 38650 30579 38652
rect 30635 38650 30659 38652
rect 30715 38650 30739 38652
rect 30795 38650 30801 38652
rect 30555 38598 30557 38650
rect 30737 38598 30739 38650
rect 30493 38596 30499 38598
rect 30555 38596 30579 38598
rect 30635 38596 30659 38598
rect 30715 38596 30739 38598
rect 30795 38596 30801 38598
rect 30493 38587 30801 38596
rect 17831 38108 18139 38117
rect 17831 38106 17837 38108
rect 17893 38106 17917 38108
rect 17973 38106 17997 38108
rect 18053 38106 18077 38108
rect 18133 38106 18139 38108
rect 17893 38054 17895 38106
rect 18075 38054 18077 38106
rect 17831 38052 17837 38054
rect 17893 38052 17917 38054
rect 17973 38052 17997 38054
rect 18053 38052 18077 38054
rect 18133 38052 18139 38054
rect 17831 38043 18139 38052
rect 26272 38108 26580 38117
rect 26272 38106 26278 38108
rect 26334 38106 26358 38108
rect 26414 38106 26438 38108
rect 26494 38106 26518 38108
rect 26574 38106 26580 38108
rect 26334 38054 26336 38106
rect 26516 38054 26518 38106
rect 26272 38052 26278 38054
rect 26334 38052 26358 38054
rect 26414 38052 26438 38054
rect 26494 38052 26518 38054
rect 26574 38052 26580 38054
rect 26272 38043 26580 38052
rect 22052 37564 22360 37573
rect 22052 37562 22058 37564
rect 22114 37562 22138 37564
rect 22194 37562 22218 37564
rect 22274 37562 22298 37564
rect 22354 37562 22360 37564
rect 22114 37510 22116 37562
rect 22296 37510 22298 37562
rect 22052 37508 22058 37510
rect 22114 37508 22138 37510
rect 22194 37508 22218 37510
rect 22274 37508 22298 37510
rect 22354 37508 22360 37510
rect 22052 37499 22360 37508
rect 30493 37564 30801 37573
rect 30493 37562 30499 37564
rect 30555 37562 30579 37564
rect 30635 37562 30659 37564
rect 30715 37562 30739 37564
rect 30795 37562 30801 37564
rect 30555 37510 30557 37562
rect 30737 37510 30739 37562
rect 30493 37508 30499 37510
rect 30555 37508 30579 37510
rect 30635 37508 30659 37510
rect 30715 37508 30739 37510
rect 30795 37508 30801 37510
rect 30493 37499 30801 37508
rect 17831 37020 18139 37029
rect 17831 37018 17837 37020
rect 17893 37018 17917 37020
rect 17973 37018 17997 37020
rect 18053 37018 18077 37020
rect 18133 37018 18139 37020
rect 17893 36966 17895 37018
rect 18075 36966 18077 37018
rect 17831 36964 17837 36966
rect 17893 36964 17917 36966
rect 17973 36964 17997 36966
rect 18053 36964 18077 36966
rect 18133 36964 18139 36966
rect 17831 36955 18139 36964
rect 26272 37020 26580 37029
rect 26272 37018 26278 37020
rect 26334 37018 26358 37020
rect 26414 37018 26438 37020
rect 26494 37018 26518 37020
rect 26574 37018 26580 37020
rect 26334 36966 26336 37018
rect 26516 36966 26518 37018
rect 26272 36964 26278 36966
rect 26334 36964 26358 36966
rect 26414 36964 26438 36966
rect 26494 36964 26518 36966
rect 26574 36964 26580 36966
rect 26272 36955 26580 36964
rect 22052 36476 22360 36485
rect 22052 36474 22058 36476
rect 22114 36474 22138 36476
rect 22194 36474 22218 36476
rect 22274 36474 22298 36476
rect 22354 36474 22360 36476
rect 22114 36422 22116 36474
rect 22296 36422 22298 36474
rect 22052 36420 22058 36422
rect 22114 36420 22138 36422
rect 22194 36420 22218 36422
rect 22274 36420 22298 36422
rect 22354 36420 22360 36422
rect 22052 36411 22360 36420
rect 30493 36476 30801 36485
rect 30493 36474 30499 36476
rect 30555 36474 30579 36476
rect 30635 36474 30659 36476
rect 30715 36474 30739 36476
rect 30795 36474 30801 36476
rect 30555 36422 30557 36474
rect 30737 36422 30739 36474
rect 30493 36420 30499 36422
rect 30555 36420 30579 36422
rect 30635 36420 30659 36422
rect 30715 36420 30739 36422
rect 30795 36420 30801 36422
rect 30493 36411 30801 36420
rect 17831 35932 18139 35941
rect 17831 35930 17837 35932
rect 17893 35930 17917 35932
rect 17973 35930 17997 35932
rect 18053 35930 18077 35932
rect 18133 35930 18139 35932
rect 17893 35878 17895 35930
rect 18075 35878 18077 35930
rect 17831 35876 17837 35878
rect 17893 35876 17917 35878
rect 17973 35876 17997 35878
rect 18053 35876 18077 35878
rect 18133 35876 18139 35878
rect 17831 35867 18139 35876
rect 26272 35932 26580 35941
rect 26272 35930 26278 35932
rect 26334 35930 26358 35932
rect 26414 35930 26438 35932
rect 26494 35930 26518 35932
rect 26574 35930 26580 35932
rect 26334 35878 26336 35930
rect 26516 35878 26518 35930
rect 26272 35876 26278 35878
rect 26334 35876 26358 35878
rect 26414 35876 26438 35878
rect 26494 35876 26518 35878
rect 26574 35876 26580 35878
rect 26272 35867 26580 35876
rect 22052 35388 22360 35397
rect 22052 35386 22058 35388
rect 22114 35386 22138 35388
rect 22194 35386 22218 35388
rect 22274 35386 22298 35388
rect 22354 35386 22360 35388
rect 22114 35334 22116 35386
rect 22296 35334 22298 35386
rect 22052 35332 22058 35334
rect 22114 35332 22138 35334
rect 22194 35332 22218 35334
rect 22274 35332 22298 35334
rect 22354 35332 22360 35334
rect 22052 35323 22360 35332
rect 30493 35388 30801 35397
rect 30493 35386 30499 35388
rect 30555 35386 30579 35388
rect 30635 35386 30659 35388
rect 30715 35386 30739 35388
rect 30795 35386 30801 35388
rect 30555 35334 30557 35386
rect 30737 35334 30739 35386
rect 30493 35332 30499 35334
rect 30555 35332 30579 35334
rect 30635 35332 30659 35334
rect 30715 35332 30739 35334
rect 30795 35332 30801 35334
rect 30493 35323 30801 35332
rect 17831 34844 18139 34853
rect 17831 34842 17837 34844
rect 17893 34842 17917 34844
rect 17973 34842 17997 34844
rect 18053 34842 18077 34844
rect 18133 34842 18139 34844
rect 17893 34790 17895 34842
rect 18075 34790 18077 34842
rect 17831 34788 17837 34790
rect 17893 34788 17917 34790
rect 17973 34788 17997 34790
rect 18053 34788 18077 34790
rect 18133 34788 18139 34790
rect 17831 34779 18139 34788
rect 26272 34844 26580 34853
rect 26272 34842 26278 34844
rect 26334 34842 26358 34844
rect 26414 34842 26438 34844
rect 26494 34842 26518 34844
rect 26574 34842 26580 34844
rect 26334 34790 26336 34842
rect 26516 34790 26518 34842
rect 26272 34788 26278 34790
rect 26334 34788 26358 34790
rect 26414 34788 26438 34790
rect 26494 34788 26518 34790
rect 26574 34788 26580 34790
rect 26272 34779 26580 34788
rect 22052 34300 22360 34309
rect 22052 34298 22058 34300
rect 22114 34298 22138 34300
rect 22194 34298 22218 34300
rect 22274 34298 22298 34300
rect 22354 34298 22360 34300
rect 22114 34246 22116 34298
rect 22296 34246 22298 34298
rect 22052 34244 22058 34246
rect 22114 34244 22138 34246
rect 22194 34244 22218 34246
rect 22274 34244 22298 34246
rect 22354 34244 22360 34246
rect 22052 34235 22360 34244
rect 30493 34300 30801 34309
rect 30493 34298 30499 34300
rect 30555 34298 30579 34300
rect 30635 34298 30659 34300
rect 30715 34298 30739 34300
rect 30795 34298 30801 34300
rect 30555 34246 30557 34298
rect 30737 34246 30739 34298
rect 30493 34244 30499 34246
rect 30555 34244 30579 34246
rect 30635 34244 30659 34246
rect 30715 34244 30739 34246
rect 30795 34244 30801 34246
rect 30493 34235 30801 34244
rect 25964 33992 26016 33998
rect 25964 33934 26016 33940
rect 17831 33756 18139 33765
rect 17831 33754 17837 33756
rect 17893 33754 17917 33756
rect 17973 33754 17997 33756
rect 18053 33754 18077 33756
rect 18133 33754 18139 33756
rect 17893 33702 17895 33754
rect 18075 33702 18077 33754
rect 17831 33700 17837 33702
rect 17893 33700 17917 33702
rect 17973 33700 17997 33702
rect 18053 33700 18077 33702
rect 18133 33700 18139 33702
rect 17831 33691 18139 33700
rect 23940 33516 23992 33522
rect 23940 33458 23992 33464
rect 25504 33516 25556 33522
rect 25504 33458 25556 33464
rect 23848 33448 23900 33454
rect 23848 33390 23900 33396
rect 23480 33312 23532 33318
rect 23480 33254 23532 33260
rect 22052 33212 22360 33221
rect 22052 33210 22058 33212
rect 22114 33210 22138 33212
rect 22194 33210 22218 33212
rect 22274 33210 22298 33212
rect 22354 33210 22360 33212
rect 22114 33158 22116 33210
rect 22296 33158 22298 33210
rect 22052 33156 22058 33158
rect 22114 33156 22138 33158
rect 22194 33156 22218 33158
rect 22274 33156 22298 33158
rect 22354 33156 22360 33158
rect 22052 33147 22360 33156
rect 23388 32972 23440 32978
rect 23388 32914 23440 32920
rect 17831 32668 18139 32677
rect 17831 32666 17837 32668
rect 17893 32666 17917 32668
rect 17973 32666 17997 32668
rect 18053 32666 18077 32668
rect 18133 32666 18139 32668
rect 17893 32614 17895 32666
rect 18075 32614 18077 32666
rect 17831 32612 17837 32614
rect 17893 32612 17917 32614
rect 17973 32612 17997 32614
rect 18053 32612 18077 32614
rect 18133 32612 18139 32614
rect 17831 32603 18139 32612
rect 23400 32434 23428 32914
rect 23492 32910 23520 33254
rect 23860 32994 23888 33390
rect 23952 33114 23980 33458
rect 24492 33312 24544 33318
rect 24492 33254 24544 33260
rect 23940 33108 23992 33114
rect 23940 33050 23992 33056
rect 23860 32966 23980 32994
rect 23952 32910 23980 32966
rect 24504 32910 24532 33254
rect 23480 32904 23532 32910
rect 23480 32846 23532 32852
rect 23940 32904 23992 32910
rect 23940 32846 23992 32852
rect 24308 32904 24360 32910
rect 24308 32846 24360 32852
rect 24492 32904 24544 32910
rect 24492 32846 24544 32852
rect 18328 32428 18380 32434
rect 18328 32370 18380 32376
rect 18696 32428 18748 32434
rect 18696 32370 18748 32376
rect 20536 32428 20588 32434
rect 20536 32370 20588 32376
rect 20996 32428 21048 32434
rect 20996 32370 21048 32376
rect 21732 32428 21784 32434
rect 21732 32370 21784 32376
rect 23388 32428 23440 32434
rect 23388 32370 23440 32376
rect 18144 32360 18196 32366
rect 18144 32302 18196 32308
rect 17776 32224 17828 32230
rect 17776 32166 17828 32172
rect 17788 31754 17816 32166
rect 18156 32026 18184 32302
rect 18144 32020 18196 32026
rect 18144 31962 18196 31968
rect 17696 31726 17816 31754
rect 18156 31754 18184 31962
rect 18156 31726 18276 31754
rect 17696 31414 17724 31726
rect 17831 31580 18139 31589
rect 17831 31578 17837 31580
rect 17893 31578 17917 31580
rect 17973 31578 17997 31580
rect 18053 31578 18077 31580
rect 18133 31578 18139 31580
rect 17893 31526 17895 31578
rect 18075 31526 18077 31578
rect 17831 31524 17837 31526
rect 17893 31524 17917 31526
rect 17973 31524 17997 31526
rect 18053 31524 18077 31526
rect 18133 31524 18139 31526
rect 17831 31515 18139 31524
rect 18248 31482 18276 31726
rect 18236 31476 18288 31482
rect 18236 31418 18288 31424
rect 17684 31408 17736 31414
rect 17684 31350 17736 31356
rect 17328 31062 17632 31090
rect 16764 30932 16816 30938
rect 16764 30874 16816 30880
rect 17132 30728 17184 30734
rect 17132 30670 17184 30676
rect 16764 30252 16816 30258
rect 16764 30194 16816 30200
rect 16672 30184 16724 30190
rect 16672 30126 16724 30132
rect 16396 30048 16448 30054
rect 16396 29990 16448 29996
rect 16488 30048 16540 30054
rect 16488 29990 16540 29996
rect 16408 29102 16436 29990
rect 16500 29850 16528 29990
rect 16488 29844 16540 29850
rect 16488 29786 16540 29792
rect 16396 29096 16448 29102
rect 16396 29038 16448 29044
rect 16684 28762 16712 30126
rect 16776 29850 16804 30194
rect 17040 30048 17092 30054
rect 17144 30002 17172 30670
rect 17092 29996 17172 30002
rect 17040 29990 17172 29996
rect 17052 29974 17172 29990
rect 17144 29850 17172 29974
rect 16764 29844 16816 29850
rect 16764 29786 16816 29792
rect 17132 29844 17184 29850
rect 17132 29786 17184 29792
rect 17328 29050 17356 31062
rect 17696 30938 17724 31350
rect 18340 31278 18368 32370
rect 18708 32026 18736 32370
rect 19800 32292 19852 32298
rect 19800 32234 19852 32240
rect 20444 32292 20496 32298
rect 20444 32234 20496 32240
rect 19812 32026 19840 32234
rect 20456 32026 20484 32234
rect 18696 32020 18748 32026
rect 18696 31962 18748 31968
rect 19800 32020 19852 32026
rect 19800 31962 19852 31968
rect 20444 32020 20496 32026
rect 20444 31962 20496 31968
rect 18512 31816 18564 31822
rect 18512 31758 18564 31764
rect 18972 31816 19024 31822
rect 18972 31758 19024 31764
rect 20168 31816 20220 31822
rect 20168 31758 20220 31764
rect 18420 31340 18472 31346
rect 18420 31282 18472 31288
rect 18328 31272 18380 31278
rect 18328 31214 18380 31220
rect 17960 31136 18012 31142
rect 17960 31078 18012 31084
rect 17592 30932 17644 30938
rect 17592 30874 17644 30880
rect 17684 30932 17736 30938
rect 17684 30874 17736 30880
rect 17500 30592 17552 30598
rect 17420 30540 17500 30546
rect 17420 30534 17552 30540
rect 17420 30518 17540 30534
rect 17420 29510 17448 30518
rect 17604 30394 17632 30874
rect 17972 30666 18000 31078
rect 18432 30938 18460 31282
rect 18420 30932 18472 30938
rect 18420 30874 18472 30880
rect 17960 30660 18012 30666
rect 17960 30602 18012 30608
rect 18236 30592 18288 30598
rect 18236 30534 18288 30540
rect 17831 30492 18139 30501
rect 17831 30490 17837 30492
rect 17893 30490 17917 30492
rect 17973 30490 17997 30492
rect 18053 30490 18077 30492
rect 18133 30490 18139 30492
rect 17893 30438 17895 30490
rect 18075 30438 18077 30490
rect 17831 30436 17837 30438
rect 17893 30436 17917 30438
rect 17973 30436 17997 30438
rect 18053 30436 18077 30438
rect 18133 30436 18139 30438
rect 17831 30427 18139 30436
rect 17592 30388 17644 30394
rect 17592 30330 17644 30336
rect 17604 29714 17632 30330
rect 18248 30326 18276 30534
rect 18236 30320 18288 30326
rect 18236 30262 18288 30268
rect 18328 30252 18380 30258
rect 18328 30194 18380 30200
rect 18340 29850 18368 30194
rect 18328 29844 18380 29850
rect 18328 29786 18380 29792
rect 17592 29708 17644 29714
rect 17592 29650 17644 29656
rect 17408 29504 17460 29510
rect 17408 29446 17460 29452
rect 17420 29238 17448 29446
rect 17831 29404 18139 29413
rect 17831 29402 17837 29404
rect 17893 29402 17917 29404
rect 17973 29402 17997 29404
rect 18053 29402 18077 29404
rect 18133 29402 18139 29404
rect 17893 29350 17895 29402
rect 18075 29350 18077 29402
rect 17831 29348 17837 29350
rect 17893 29348 17917 29350
rect 17973 29348 17997 29350
rect 18053 29348 18077 29350
rect 18133 29348 18139 29350
rect 17831 29339 18139 29348
rect 17408 29232 17460 29238
rect 17408 29174 17460 29180
rect 17776 29164 17828 29170
rect 17776 29106 17828 29112
rect 17328 29022 17448 29050
rect 17040 28960 17092 28966
rect 17040 28902 17092 28908
rect 16672 28756 16724 28762
rect 16672 28698 16724 28704
rect 16856 28484 16908 28490
rect 16856 28426 16908 28432
rect 16868 28218 16896 28426
rect 16856 28212 16908 28218
rect 16856 28154 16908 28160
rect 17052 28082 17080 28902
rect 17040 28076 17092 28082
rect 17040 28018 17092 28024
rect 16672 27464 16724 27470
rect 16672 27406 16724 27412
rect 16684 26314 16712 27406
rect 16856 27124 16908 27130
rect 16856 27066 16908 27072
rect 16868 26382 16896 27066
rect 17316 26988 17368 26994
rect 17316 26930 17368 26936
rect 16948 26784 17000 26790
rect 16948 26726 17000 26732
rect 16856 26376 16908 26382
rect 16856 26318 16908 26324
rect 16672 26308 16724 26314
rect 16672 26250 16724 26256
rect 16960 25294 16988 26726
rect 17132 25900 17184 25906
rect 17132 25842 17184 25848
rect 17144 25498 17172 25842
rect 17328 25838 17356 26930
rect 17420 26246 17448 29022
rect 17788 28762 17816 29106
rect 18432 29102 18460 30874
rect 18524 30870 18552 31758
rect 18984 31482 19012 31758
rect 19800 31748 19852 31754
rect 19800 31690 19852 31696
rect 19524 31680 19576 31686
rect 19524 31622 19576 31628
rect 19708 31680 19760 31686
rect 19708 31622 19760 31628
rect 18880 31476 18932 31482
rect 18880 31418 18932 31424
rect 18972 31476 19024 31482
rect 18972 31418 19024 31424
rect 18892 30870 18920 31418
rect 19536 31142 19564 31622
rect 19720 31346 19748 31622
rect 19708 31340 19760 31346
rect 19708 31282 19760 31288
rect 19156 31136 19208 31142
rect 19156 31078 19208 31084
rect 19524 31136 19576 31142
rect 19524 31078 19576 31084
rect 18512 30864 18564 30870
rect 18512 30806 18564 30812
rect 18880 30864 18932 30870
rect 18880 30806 18932 30812
rect 19168 30818 19196 31078
rect 18524 30274 18552 30806
rect 18892 30734 18920 30806
rect 19064 30796 19116 30802
rect 19064 30738 19116 30744
rect 19168 30790 19380 30818
rect 18696 30728 18748 30734
rect 18694 30696 18696 30705
rect 18880 30728 18932 30734
rect 18748 30696 18750 30705
rect 18880 30670 18932 30676
rect 18694 30631 18750 30640
rect 19076 30394 19104 30738
rect 19064 30388 19116 30394
rect 19064 30330 19116 30336
rect 18524 30246 18644 30274
rect 19168 30258 19196 30790
rect 19352 30734 19380 30790
rect 19536 30734 19564 31078
rect 19812 30870 19840 31690
rect 20180 31346 20208 31758
rect 20260 31680 20312 31686
rect 20260 31622 20312 31628
rect 20352 31680 20404 31686
rect 20352 31622 20404 31628
rect 20272 31346 20300 31622
rect 20168 31340 20220 31346
rect 20168 31282 20220 31288
rect 20260 31340 20312 31346
rect 20260 31282 20312 31288
rect 19984 31136 20036 31142
rect 19984 31078 20036 31084
rect 19800 30864 19852 30870
rect 19800 30806 19852 30812
rect 19996 30802 20024 31078
rect 19984 30796 20036 30802
rect 19984 30738 20036 30744
rect 19340 30728 19392 30734
rect 19246 30696 19302 30705
rect 19340 30670 19392 30676
rect 19524 30728 19576 30734
rect 19524 30670 19576 30676
rect 19246 30631 19302 30640
rect 19260 30598 19288 30631
rect 19248 30592 19300 30598
rect 19248 30534 19300 30540
rect 19536 30326 19564 30670
rect 19524 30320 19576 30326
rect 19524 30262 19576 30268
rect 18616 29730 18644 30246
rect 19156 30252 19208 30258
rect 19156 30194 19208 30200
rect 19248 30252 19300 30258
rect 19248 30194 19300 30200
rect 19156 30048 19208 30054
rect 19156 29990 19208 29996
rect 19168 29850 19196 29990
rect 19260 29850 19288 30194
rect 20076 30048 20128 30054
rect 20076 29990 20128 29996
rect 19156 29844 19208 29850
rect 19156 29786 19208 29792
rect 19248 29844 19300 29850
rect 19248 29786 19300 29792
rect 18524 29702 18644 29730
rect 19892 29776 19944 29782
rect 19892 29718 19944 29724
rect 18420 29096 18472 29102
rect 18420 29038 18472 29044
rect 17776 28756 17828 28762
rect 17776 28698 17828 28704
rect 18328 28756 18380 28762
rect 18328 28698 18380 28704
rect 18236 28552 18288 28558
rect 18236 28494 18288 28500
rect 17500 28416 17552 28422
rect 17500 28358 17552 28364
rect 17512 28082 17540 28358
rect 17831 28316 18139 28325
rect 17831 28314 17837 28316
rect 17893 28314 17917 28316
rect 17973 28314 17997 28316
rect 18053 28314 18077 28316
rect 18133 28314 18139 28316
rect 17893 28262 17895 28314
rect 18075 28262 18077 28314
rect 17831 28260 17837 28262
rect 17893 28260 17917 28262
rect 17973 28260 17997 28262
rect 18053 28260 18077 28262
rect 18133 28260 18139 28262
rect 17831 28251 18139 28260
rect 17500 28076 17552 28082
rect 17500 28018 17552 28024
rect 18144 28076 18196 28082
rect 18144 28018 18196 28024
rect 17512 27334 17540 28018
rect 17960 28008 18012 28014
rect 17960 27950 18012 27956
rect 17972 27674 18000 27950
rect 18052 27872 18104 27878
rect 18052 27814 18104 27820
rect 17960 27668 18012 27674
rect 17960 27610 18012 27616
rect 17972 27470 18000 27610
rect 18064 27606 18092 27814
rect 18156 27674 18184 28018
rect 18144 27668 18196 27674
rect 18144 27610 18196 27616
rect 18052 27600 18104 27606
rect 18052 27542 18104 27548
rect 17960 27464 18012 27470
rect 17960 27406 18012 27412
rect 17500 27328 17552 27334
rect 17500 27270 17552 27276
rect 17512 26858 17540 27270
rect 17831 27228 18139 27237
rect 17831 27226 17837 27228
rect 17893 27226 17917 27228
rect 17973 27226 17997 27228
rect 18053 27226 18077 27228
rect 18133 27226 18139 27228
rect 17893 27174 17895 27226
rect 18075 27174 18077 27226
rect 17831 27172 17837 27174
rect 17893 27172 17917 27174
rect 17973 27172 17997 27174
rect 18053 27172 18077 27174
rect 18133 27172 18139 27174
rect 17831 27163 18139 27172
rect 18248 27130 18276 28494
rect 18340 28082 18368 28698
rect 18420 28484 18472 28490
rect 18420 28426 18472 28432
rect 18432 28218 18460 28426
rect 18420 28212 18472 28218
rect 18420 28154 18472 28160
rect 18328 28076 18380 28082
rect 18328 28018 18380 28024
rect 18420 27396 18472 27402
rect 18420 27338 18472 27344
rect 18236 27124 18288 27130
rect 18236 27066 18288 27072
rect 18432 26994 18460 27338
rect 17684 26988 17736 26994
rect 17604 26948 17684 26976
rect 17500 26852 17552 26858
rect 17500 26794 17552 26800
rect 17408 26240 17460 26246
rect 17408 26182 17460 26188
rect 17512 26042 17540 26794
rect 17604 26382 17632 26948
rect 17684 26930 17736 26936
rect 17868 26988 17920 26994
rect 17868 26930 17920 26936
rect 18420 26988 18472 26994
rect 18420 26930 18472 26936
rect 17880 26586 17908 26930
rect 18236 26920 18288 26926
rect 18236 26862 18288 26868
rect 17684 26580 17736 26586
rect 17684 26522 17736 26528
rect 17868 26580 17920 26586
rect 17868 26522 17920 26528
rect 17592 26376 17644 26382
rect 17592 26318 17644 26324
rect 17500 26036 17552 26042
rect 17500 25978 17552 25984
rect 17316 25832 17368 25838
rect 17604 25820 17632 26318
rect 17696 25922 17724 26522
rect 17831 26140 18139 26149
rect 17831 26138 17837 26140
rect 17893 26138 17917 26140
rect 17973 26138 17997 26140
rect 18053 26138 18077 26140
rect 18133 26138 18139 26140
rect 17893 26086 17895 26138
rect 18075 26086 18077 26138
rect 17831 26084 17837 26086
rect 17893 26084 17917 26086
rect 17973 26084 17997 26086
rect 18053 26084 18077 26086
rect 18133 26084 18139 26086
rect 17831 26075 18139 26084
rect 17776 25968 17828 25974
rect 17696 25916 17776 25922
rect 17696 25910 17828 25916
rect 17696 25894 17816 25910
rect 17960 25900 18012 25906
rect 17880 25860 17960 25888
rect 17880 25820 17908 25860
rect 17960 25842 18012 25848
rect 17604 25792 17908 25820
rect 17316 25774 17368 25780
rect 17224 25696 17276 25702
rect 17224 25638 17276 25644
rect 17132 25492 17184 25498
rect 17132 25434 17184 25440
rect 16948 25288 17000 25294
rect 17000 25236 17080 25242
rect 16948 25230 17080 25236
rect 16960 25214 17080 25230
rect 16948 25152 17000 25158
rect 16948 25094 17000 25100
rect 16960 24886 16988 25094
rect 16948 24880 17000 24886
rect 16948 24822 17000 24828
rect 16948 24608 17000 24614
rect 16948 24550 17000 24556
rect 16960 24274 16988 24550
rect 16948 24268 17000 24274
rect 16948 24210 17000 24216
rect 17052 23118 17080 25214
rect 17144 24954 17172 25434
rect 17236 25158 17264 25638
rect 18248 25498 18276 26862
rect 18524 26790 18552 29702
rect 18604 29640 18656 29646
rect 18604 29582 18656 29588
rect 18696 29640 18748 29646
rect 18696 29582 18748 29588
rect 18880 29640 18932 29646
rect 18880 29582 18932 29588
rect 18616 29306 18644 29582
rect 18604 29300 18656 29306
rect 18604 29242 18656 29248
rect 18616 28422 18644 29242
rect 18708 28558 18736 29582
rect 18892 28762 18920 29582
rect 19904 29238 19932 29718
rect 20088 29714 20116 29990
rect 20076 29708 20128 29714
rect 20076 29650 20128 29656
rect 19892 29232 19944 29238
rect 19892 29174 19944 29180
rect 20088 29170 20116 29650
rect 20180 29578 20208 31282
rect 20364 31210 20392 31622
rect 20444 31408 20496 31414
rect 20444 31350 20496 31356
rect 20352 31204 20404 31210
rect 20352 31146 20404 31152
rect 20456 31142 20484 31350
rect 20548 31260 20576 32370
rect 20720 32360 20772 32366
rect 20720 32302 20772 32308
rect 20628 32224 20680 32230
rect 20628 32166 20680 32172
rect 20640 31958 20668 32166
rect 20628 31952 20680 31958
rect 20628 31894 20680 31900
rect 20640 31482 20668 31894
rect 20628 31476 20680 31482
rect 20628 31418 20680 31424
rect 20732 31414 20760 32302
rect 21008 32026 21036 32370
rect 21180 32224 21232 32230
rect 21180 32166 21232 32172
rect 21192 32026 21220 32166
rect 21744 32026 21772 32370
rect 21824 32224 21876 32230
rect 21824 32166 21876 32172
rect 21916 32224 21968 32230
rect 21916 32166 21968 32172
rect 20996 32020 21048 32026
rect 20996 31962 21048 31968
rect 21180 32020 21232 32026
rect 21180 31962 21232 31968
rect 21732 32020 21784 32026
rect 21732 31962 21784 31968
rect 20904 31816 20956 31822
rect 20904 31758 20956 31764
rect 20812 31680 20864 31686
rect 20812 31622 20864 31628
rect 20720 31408 20772 31414
rect 20720 31350 20772 31356
rect 20720 31272 20772 31278
rect 20548 31232 20720 31260
rect 20720 31214 20772 31220
rect 20444 31136 20496 31142
rect 20444 31078 20496 31084
rect 20260 30796 20312 30802
rect 20260 30738 20312 30744
rect 20272 30394 20300 30738
rect 20260 30388 20312 30394
rect 20260 30330 20312 30336
rect 20824 30258 20852 31622
rect 20916 30410 20944 31758
rect 21008 31482 21036 31962
rect 21836 31958 21864 32166
rect 21824 31952 21876 31958
rect 21824 31894 21876 31900
rect 21928 31822 21956 32166
rect 22052 32124 22360 32133
rect 22052 32122 22058 32124
rect 22114 32122 22138 32124
rect 22194 32122 22218 32124
rect 22274 32122 22298 32124
rect 22354 32122 22360 32124
rect 22114 32070 22116 32122
rect 22296 32070 22298 32122
rect 22052 32068 22058 32070
rect 22114 32068 22138 32070
rect 22194 32068 22218 32070
rect 22274 32068 22298 32070
rect 22354 32068 22360 32070
rect 22052 32059 22360 32068
rect 21456 31816 21508 31822
rect 21376 31764 21456 31770
rect 21376 31758 21508 31764
rect 21548 31816 21600 31822
rect 21548 31758 21600 31764
rect 21824 31816 21876 31822
rect 21824 31758 21876 31764
rect 21916 31816 21968 31822
rect 21916 31758 21968 31764
rect 21376 31754 21496 31758
rect 21192 31742 21496 31754
rect 21192 31726 21404 31742
rect 20996 31476 21048 31482
rect 20996 31418 21048 31424
rect 20916 30382 21128 30410
rect 20260 30252 20312 30258
rect 20260 30194 20312 30200
rect 20444 30252 20496 30258
rect 20812 30252 20864 30258
rect 20444 30194 20496 30200
rect 20732 30212 20812 30240
rect 20168 29572 20220 29578
rect 20168 29514 20220 29520
rect 20272 29170 20300 30194
rect 20352 30116 20404 30122
rect 20352 30058 20404 30064
rect 20364 29714 20392 30058
rect 20352 29708 20404 29714
rect 20352 29650 20404 29656
rect 20352 29504 20404 29510
rect 20352 29446 20404 29452
rect 20364 29209 20392 29446
rect 20456 29306 20484 30194
rect 20536 30184 20588 30190
rect 20536 30126 20588 30132
rect 20548 29782 20576 30126
rect 20628 30116 20680 30122
rect 20628 30058 20680 30064
rect 20536 29776 20588 29782
rect 20536 29718 20588 29724
rect 20640 29306 20668 30058
rect 20444 29300 20496 29306
rect 20444 29242 20496 29248
rect 20628 29300 20680 29306
rect 20628 29242 20680 29248
rect 20350 29200 20406 29209
rect 20076 29164 20128 29170
rect 20076 29106 20128 29112
rect 20260 29164 20312 29170
rect 20732 29186 20760 30212
rect 20812 30194 20864 30200
rect 20904 30252 20956 30258
rect 20904 30194 20956 30200
rect 20916 29850 20944 30194
rect 20996 30184 21048 30190
rect 20996 30126 21048 30132
rect 20904 29844 20956 29850
rect 20904 29786 20956 29792
rect 20812 29640 20864 29646
rect 20812 29582 20864 29588
rect 20350 29135 20406 29144
rect 20640 29158 20760 29186
rect 20260 29106 20312 29112
rect 18880 28756 18932 28762
rect 18880 28698 18932 28704
rect 18696 28552 18748 28558
rect 18696 28494 18748 28500
rect 18604 28416 18656 28422
rect 18604 28358 18656 28364
rect 18708 28014 18736 28494
rect 18972 28076 19024 28082
rect 18972 28018 19024 28024
rect 19340 28076 19392 28082
rect 19340 28018 19392 28024
rect 18696 28008 18748 28014
rect 18696 27950 18748 27956
rect 18880 27532 18932 27538
rect 18880 27474 18932 27480
rect 18512 26784 18564 26790
rect 18512 26726 18564 26732
rect 18512 26580 18564 26586
rect 18512 26522 18564 26528
rect 18524 26314 18552 26522
rect 18892 26518 18920 27474
rect 18984 27334 19012 28018
rect 19352 27334 19380 28018
rect 20088 28014 20116 29106
rect 20272 29034 20300 29106
rect 20260 29028 20312 29034
rect 20260 28970 20312 28976
rect 20640 28642 20668 29158
rect 20720 29096 20772 29102
rect 20720 29038 20772 29044
rect 20732 28762 20760 29038
rect 20824 29034 20852 29582
rect 21008 29306 21036 30126
rect 20996 29300 21048 29306
rect 20996 29242 21048 29248
rect 20902 29200 20958 29209
rect 21100 29186 21128 30382
rect 21192 30258 21220 31726
rect 21560 31346 21588 31758
rect 21548 31340 21600 31346
rect 21548 31282 21600 31288
rect 21836 31278 21864 31758
rect 21916 31680 21968 31686
rect 21916 31622 21968 31628
rect 21928 31414 21956 31622
rect 23400 31482 23428 32370
rect 23952 31822 23980 32846
rect 24320 32026 24348 32846
rect 25516 32230 25544 33458
rect 25596 33108 25648 33114
rect 25596 33050 25648 33056
rect 25608 32502 25636 33050
rect 25976 32858 26004 33934
rect 26884 33924 26936 33930
rect 26884 33866 26936 33872
rect 26148 33856 26200 33862
rect 26148 33798 26200 33804
rect 26792 33856 26844 33862
rect 26792 33798 26844 33804
rect 26160 33454 26188 33798
rect 26272 33756 26580 33765
rect 26272 33754 26278 33756
rect 26334 33754 26358 33756
rect 26414 33754 26438 33756
rect 26494 33754 26518 33756
rect 26574 33754 26580 33756
rect 26334 33702 26336 33754
rect 26516 33702 26518 33754
rect 26272 33700 26278 33702
rect 26334 33700 26358 33702
rect 26414 33700 26438 33702
rect 26494 33700 26518 33702
rect 26574 33700 26580 33702
rect 26272 33691 26580 33700
rect 26804 33658 26832 33798
rect 26792 33652 26844 33658
rect 26792 33594 26844 33600
rect 26148 33448 26200 33454
rect 26148 33390 26200 33396
rect 26608 33448 26660 33454
rect 26608 33390 26660 33396
rect 26240 33380 26292 33386
rect 26240 33322 26292 33328
rect 26252 33130 26280 33322
rect 26332 33312 26384 33318
rect 26332 33254 26384 33260
rect 26160 33102 26280 33130
rect 26160 33046 26188 33102
rect 26148 33040 26200 33046
rect 26344 32994 26372 33254
rect 26148 32982 26200 32988
rect 26252 32966 26372 32994
rect 26252 32910 26280 32966
rect 26240 32904 26292 32910
rect 25700 32830 26004 32858
rect 25700 32774 25728 32830
rect 25688 32768 25740 32774
rect 25688 32710 25740 32716
rect 25872 32768 25924 32774
rect 25872 32710 25924 32716
rect 25596 32496 25648 32502
rect 25596 32438 25648 32444
rect 25504 32224 25556 32230
rect 25504 32166 25556 32172
rect 24308 32020 24360 32026
rect 24308 31962 24360 31968
rect 23940 31816 23992 31822
rect 23940 31758 23992 31764
rect 23388 31476 23440 31482
rect 23388 31418 23440 31424
rect 21916 31408 21968 31414
rect 21916 31350 21968 31356
rect 23296 31340 23348 31346
rect 23296 31282 23348 31288
rect 21272 31272 21324 31278
rect 21272 31214 21324 31220
rect 21824 31272 21876 31278
rect 21824 31214 21876 31220
rect 21180 30252 21232 30258
rect 21180 30194 21232 30200
rect 21008 29170 21128 29186
rect 20902 29135 20958 29144
rect 20996 29164 21128 29170
rect 20916 29102 20944 29135
rect 21048 29158 21128 29164
rect 21192 29730 21220 30194
rect 21284 30054 21312 31214
rect 22052 31036 22360 31045
rect 22052 31034 22058 31036
rect 22114 31034 22138 31036
rect 22194 31034 22218 31036
rect 22274 31034 22298 31036
rect 22354 31034 22360 31036
rect 22114 30982 22116 31034
rect 22296 30982 22298 31034
rect 22052 30980 22058 30982
rect 22114 30980 22138 30982
rect 22194 30980 22218 30982
rect 22274 30980 22298 30982
rect 22354 30980 22360 30982
rect 22052 30971 22360 30980
rect 22652 30660 22704 30666
rect 22652 30602 22704 30608
rect 21548 30116 21600 30122
rect 21548 30058 21600 30064
rect 21272 30048 21324 30054
rect 21272 29990 21324 29996
rect 21284 29850 21312 29990
rect 21560 29850 21588 30058
rect 22052 29948 22360 29957
rect 22052 29946 22058 29948
rect 22114 29946 22138 29948
rect 22194 29946 22218 29948
rect 22274 29946 22298 29948
rect 22354 29946 22360 29948
rect 22114 29894 22116 29946
rect 22296 29894 22298 29946
rect 22052 29892 22058 29894
rect 22114 29892 22138 29894
rect 22194 29892 22218 29894
rect 22274 29892 22298 29894
rect 22354 29892 22360 29894
rect 22052 29883 22360 29892
rect 22664 29850 22692 30602
rect 23112 30592 23164 30598
rect 23112 30534 23164 30540
rect 23204 30592 23256 30598
rect 23204 30534 23256 30540
rect 23124 30394 23152 30534
rect 23112 30388 23164 30394
rect 23112 30330 23164 30336
rect 21272 29844 21324 29850
rect 21272 29786 21324 29792
rect 21548 29844 21600 29850
rect 21548 29786 21600 29792
rect 22652 29844 22704 29850
rect 22652 29786 22704 29792
rect 23216 29782 23244 30534
rect 23204 29776 23256 29782
rect 21192 29702 21588 29730
rect 23204 29718 23256 29724
rect 20996 29106 21048 29112
rect 20904 29096 20956 29102
rect 20904 29038 20956 29044
rect 20812 29028 20864 29034
rect 20812 28970 20864 28976
rect 20720 28756 20772 28762
rect 20720 28698 20772 28704
rect 20640 28614 20760 28642
rect 20628 28552 20680 28558
rect 20628 28494 20680 28500
rect 20076 28008 20128 28014
rect 20076 27950 20128 27956
rect 18972 27328 19024 27334
rect 18972 27270 19024 27276
rect 19340 27328 19392 27334
rect 19340 27270 19392 27276
rect 19432 27328 19484 27334
rect 19432 27270 19484 27276
rect 18984 27062 19012 27270
rect 19352 27130 19380 27270
rect 19340 27124 19392 27130
rect 19340 27066 19392 27072
rect 19444 27062 19472 27270
rect 18972 27056 19024 27062
rect 18972 26998 19024 27004
rect 19432 27056 19484 27062
rect 19432 26998 19484 27004
rect 20088 26926 20116 27950
rect 20260 27940 20312 27946
rect 20260 27882 20312 27888
rect 20272 27470 20300 27882
rect 20640 27606 20668 28494
rect 20628 27600 20680 27606
rect 20628 27542 20680 27548
rect 20260 27464 20312 27470
rect 20260 27406 20312 27412
rect 20442 27432 20498 27441
rect 20442 27367 20444 27376
rect 20496 27367 20498 27376
rect 20444 27338 20496 27344
rect 20352 27328 20404 27334
rect 20352 27270 20404 27276
rect 20364 27062 20392 27270
rect 20352 27056 20404 27062
rect 20352 26998 20404 27004
rect 20536 26988 20588 26994
rect 20536 26930 20588 26936
rect 19708 26920 19760 26926
rect 20076 26920 20128 26926
rect 19708 26862 19760 26868
rect 20074 26888 20076 26897
rect 20128 26888 20130 26897
rect 19432 26784 19484 26790
rect 19432 26726 19484 26732
rect 18880 26512 18932 26518
rect 18880 26454 18932 26460
rect 18512 26308 18564 26314
rect 18512 26250 18564 26256
rect 18420 25764 18472 25770
rect 18420 25706 18472 25712
rect 18328 25696 18380 25702
rect 18328 25638 18380 25644
rect 18340 25498 18368 25638
rect 18236 25492 18288 25498
rect 18236 25434 18288 25440
rect 18328 25492 18380 25498
rect 18328 25434 18380 25440
rect 17316 25424 17368 25430
rect 17316 25366 17368 25372
rect 17224 25152 17276 25158
rect 17224 25094 17276 25100
rect 17132 24948 17184 24954
rect 17132 24890 17184 24896
rect 17328 24206 17356 25366
rect 18236 25152 18288 25158
rect 18236 25094 18288 25100
rect 17831 25052 18139 25061
rect 17831 25050 17837 25052
rect 17893 25050 17917 25052
rect 17973 25050 17997 25052
rect 18053 25050 18077 25052
rect 18133 25050 18139 25052
rect 17893 24998 17895 25050
rect 18075 24998 18077 25050
rect 17831 24996 17837 24998
rect 17893 24996 17917 24998
rect 17973 24996 17997 24998
rect 18053 24996 18077 24998
rect 18133 24996 18139 24998
rect 17831 24987 18139 24996
rect 18248 24954 18276 25094
rect 18432 24954 18460 25706
rect 18236 24948 18288 24954
rect 18236 24890 18288 24896
rect 18420 24948 18472 24954
rect 18420 24890 18472 24896
rect 18236 24744 18288 24750
rect 18236 24686 18288 24692
rect 18248 24274 18276 24686
rect 18432 24410 18460 24890
rect 18524 24750 18552 26250
rect 18696 25696 18748 25702
rect 18696 25638 18748 25644
rect 18708 25498 18736 25638
rect 18696 25492 18748 25498
rect 18696 25434 18748 25440
rect 18512 24744 18564 24750
rect 18512 24686 18564 24692
rect 18420 24404 18472 24410
rect 18420 24346 18472 24352
rect 18892 24274 18920 26454
rect 19444 26382 19472 26726
rect 19720 26586 19748 26862
rect 20074 26823 20130 26832
rect 20088 26586 20116 26823
rect 19708 26580 19760 26586
rect 19708 26522 19760 26528
rect 20076 26580 20128 26586
rect 20076 26522 20128 26528
rect 20548 26382 20576 26930
rect 19432 26376 19484 26382
rect 19432 26318 19484 26324
rect 20536 26376 20588 26382
rect 20640 26353 20668 27542
rect 20732 27010 20760 28614
rect 20810 27432 20866 27441
rect 20810 27367 20866 27376
rect 20824 27334 20852 27367
rect 20812 27328 20864 27334
rect 20812 27270 20864 27276
rect 20916 27130 20944 29038
rect 21008 27538 21036 29106
rect 21088 28484 21140 28490
rect 21192 28472 21220 29702
rect 21456 29640 21508 29646
rect 21456 29582 21508 29588
rect 21468 28762 21496 29582
rect 21560 29102 21588 29702
rect 22836 29640 22888 29646
rect 22836 29582 22888 29588
rect 22848 29306 22876 29582
rect 22836 29300 22888 29306
rect 22836 29242 22888 29248
rect 23020 29164 23072 29170
rect 23020 29106 23072 29112
rect 21548 29096 21600 29102
rect 21548 29038 21600 29044
rect 21548 28960 21600 28966
rect 21548 28902 21600 28908
rect 21456 28756 21508 28762
rect 21456 28698 21508 28704
rect 21468 28558 21496 28698
rect 21560 28558 21588 28902
rect 22052 28860 22360 28869
rect 22052 28858 22058 28860
rect 22114 28858 22138 28860
rect 22194 28858 22218 28860
rect 22274 28858 22298 28860
rect 22354 28858 22360 28860
rect 22114 28806 22116 28858
rect 22296 28806 22298 28858
rect 22052 28804 22058 28806
rect 22114 28804 22138 28806
rect 22194 28804 22218 28806
rect 22274 28804 22298 28806
rect 22354 28804 22360 28806
rect 22052 28795 22360 28804
rect 23032 28558 23060 29106
rect 21456 28552 21508 28558
rect 21456 28494 21508 28500
rect 21548 28552 21600 28558
rect 21548 28494 21600 28500
rect 23020 28552 23072 28558
rect 23020 28494 23072 28500
rect 21140 28444 21220 28472
rect 21088 28426 21140 28432
rect 21100 27674 21128 28426
rect 22928 28076 22980 28082
rect 22928 28018 22980 28024
rect 22052 27772 22360 27781
rect 22052 27770 22058 27772
rect 22114 27770 22138 27772
rect 22194 27770 22218 27772
rect 22274 27770 22298 27772
rect 22354 27770 22360 27772
rect 22114 27718 22116 27770
rect 22296 27718 22298 27770
rect 22052 27716 22058 27718
rect 22114 27716 22138 27718
rect 22194 27716 22218 27718
rect 22274 27716 22298 27718
rect 22354 27716 22360 27718
rect 22052 27707 22360 27716
rect 22940 27674 22968 28018
rect 21088 27668 21140 27674
rect 21088 27610 21140 27616
rect 21824 27668 21876 27674
rect 21824 27610 21876 27616
rect 22928 27668 22980 27674
rect 22928 27610 22980 27616
rect 20996 27532 21048 27538
rect 20996 27474 21048 27480
rect 20904 27124 20956 27130
rect 20904 27066 20956 27072
rect 20810 27024 20866 27033
rect 20732 26982 20810 27010
rect 20810 26959 20866 26968
rect 20720 26920 20772 26926
rect 20720 26862 20772 26868
rect 20732 26790 20760 26862
rect 20720 26784 20772 26790
rect 20720 26726 20772 26732
rect 20732 26450 20760 26726
rect 20824 26518 20852 26959
rect 20904 26580 20956 26586
rect 20904 26522 20956 26528
rect 20812 26512 20864 26518
rect 20916 26489 20944 26522
rect 20812 26454 20864 26460
rect 20902 26480 20958 26489
rect 20720 26444 20772 26450
rect 20902 26415 20958 26424
rect 20720 26386 20772 26392
rect 20904 26376 20956 26382
rect 20536 26318 20588 26324
rect 20626 26344 20682 26353
rect 20260 26308 20312 26314
rect 20260 26250 20312 26256
rect 19156 25900 19208 25906
rect 19156 25842 19208 25848
rect 19984 25900 20036 25906
rect 19984 25842 20036 25848
rect 19168 25770 19196 25842
rect 19892 25832 19944 25838
rect 19892 25774 19944 25780
rect 19156 25764 19208 25770
rect 19156 25706 19208 25712
rect 19800 25696 19852 25702
rect 19800 25638 19852 25644
rect 19812 25498 19840 25638
rect 19904 25498 19932 25774
rect 19996 25498 20024 25842
rect 19800 25492 19852 25498
rect 19800 25434 19852 25440
rect 19892 25492 19944 25498
rect 19892 25434 19944 25440
rect 19984 25492 20036 25498
rect 19984 25434 20036 25440
rect 19340 25424 19392 25430
rect 19340 25366 19392 25372
rect 19248 24812 19300 24818
rect 19248 24754 19300 24760
rect 19260 24410 19288 24754
rect 19248 24404 19300 24410
rect 19248 24346 19300 24352
rect 18236 24268 18288 24274
rect 18236 24210 18288 24216
rect 18880 24268 18932 24274
rect 18880 24210 18932 24216
rect 17316 24200 17368 24206
rect 17316 24142 17368 24148
rect 17831 23964 18139 23973
rect 17831 23962 17837 23964
rect 17893 23962 17917 23964
rect 17973 23962 17997 23964
rect 18053 23962 18077 23964
rect 18133 23962 18139 23964
rect 17893 23910 17895 23962
rect 18075 23910 18077 23962
rect 17831 23908 17837 23910
rect 17893 23908 17917 23910
rect 17973 23908 17997 23910
rect 18053 23908 18077 23910
rect 18133 23908 18139 23910
rect 17831 23899 18139 23908
rect 17040 23112 17092 23118
rect 17040 23054 17092 23060
rect 18328 23112 18380 23118
rect 18328 23054 18380 23060
rect 16948 22568 17000 22574
rect 16948 22510 17000 22516
rect 16040 22066 16160 22094
rect 16960 22094 16988 22510
rect 17052 22250 17080 23054
rect 17408 22976 17460 22982
rect 17408 22918 17460 22924
rect 17420 22778 17448 22918
rect 17831 22876 18139 22885
rect 17831 22874 17837 22876
rect 17893 22874 17917 22876
rect 17973 22874 17997 22876
rect 18053 22874 18077 22876
rect 18133 22874 18139 22876
rect 17893 22822 17895 22874
rect 18075 22822 18077 22874
rect 17831 22820 17837 22822
rect 17893 22820 17917 22822
rect 17973 22820 17997 22822
rect 18053 22820 18077 22822
rect 18133 22820 18139 22822
rect 17831 22811 18139 22820
rect 18340 22778 18368 23054
rect 17408 22772 17460 22778
rect 17408 22714 17460 22720
rect 18328 22772 18380 22778
rect 18328 22714 18380 22720
rect 18788 22636 18840 22642
rect 18788 22578 18840 22584
rect 18604 22500 18656 22506
rect 18604 22442 18656 22448
rect 17052 22234 17264 22250
rect 17052 22228 17276 22234
rect 17052 22222 17224 22228
rect 17224 22170 17276 22176
rect 16960 22066 17172 22094
rect 9390 21788 9698 21797
rect 9390 21786 9396 21788
rect 9452 21786 9476 21788
rect 9532 21786 9556 21788
rect 9612 21786 9636 21788
rect 9692 21786 9698 21788
rect 9452 21734 9454 21786
rect 9634 21734 9636 21786
rect 9390 21732 9396 21734
rect 9452 21732 9476 21734
rect 9532 21732 9556 21734
rect 9612 21732 9636 21734
rect 9692 21732 9698 21734
rect 9390 21723 9698 21732
rect 5170 21244 5478 21253
rect 5170 21242 5176 21244
rect 5232 21242 5256 21244
rect 5312 21242 5336 21244
rect 5392 21242 5416 21244
rect 5472 21242 5478 21244
rect 5232 21190 5234 21242
rect 5414 21190 5416 21242
rect 5170 21188 5176 21190
rect 5232 21188 5256 21190
rect 5312 21188 5336 21190
rect 5392 21188 5416 21190
rect 5472 21188 5478 21190
rect 5170 21179 5478 21188
rect 13611 21244 13919 21253
rect 13611 21242 13617 21244
rect 13673 21242 13697 21244
rect 13753 21242 13777 21244
rect 13833 21242 13857 21244
rect 13913 21242 13919 21244
rect 13673 21190 13675 21242
rect 13855 21190 13857 21242
rect 13611 21188 13617 21190
rect 13673 21188 13697 21190
rect 13753 21188 13777 21190
rect 13833 21188 13857 21190
rect 13913 21188 13919 21190
rect 13611 21179 13919 21188
rect 9390 20700 9698 20709
rect 9390 20698 9396 20700
rect 9452 20698 9476 20700
rect 9532 20698 9556 20700
rect 9612 20698 9636 20700
rect 9692 20698 9698 20700
rect 9452 20646 9454 20698
rect 9634 20646 9636 20698
rect 9390 20644 9396 20646
rect 9452 20644 9476 20646
rect 9532 20644 9556 20646
rect 9612 20644 9636 20646
rect 9692 20644 9698 20646
rect 9390 20635 9698 20644
rect 5170 20156 5478 20165
rect 5170 20154 5176 20156
rect 5232 20154 5256 20156
rect 5312 20154 5336 20156
rect 5392 20154 5416 20156
rect 5472 20154 5478 20156
rect 5232 20102 5234 20154
rect 5414 20102 5416 20154
rect 5170 20100 5176 20102
rect 5232 20100 5256 20102
rect 5312 20100 5336 20102
rect 5392 20100 5416 20102
rect 5472 20100 5478 20102
rect 5170 20091 5478 20100
rect 13611 20156 13919 20165
rect 13611 20154 13617 20156
rect 13673 20154 13697 20156
rect 13753 20154 13777 20156
rect 13833 20154 13857 20156
rect 13913 20154 13919 20156
rect 13673 20102 13675 20154
rect 13855 20102 13857 20154
rect 13611 20100 13617 20102
rect 13673 20100 13697 20102
rect 13753 20100 13777 20102
rect 13833 20100 13857 20102
rect 13913 20100 13919 20102
rect 13611 20091 13919 20100
rect 940 19848 992 19854
rect 938 19816 940 19825
rect 992 19816 994 19825
rect 938 19751 994 19760
rect 9390 19612 9698 19621
rect 9390 19610 9396 19612
rect 9452 19610 9476 19612
rect 9532 19610 9556 19612
rect 9612 19610 9636 19612
rect 9692 19610 9698 19612
rect 9452 19558 9454 19610
rect 9634 19558 9636 19610
rect 9390 19556 9396 19558
rect 9452 19556 9476 19558
rect 9532 19556 9556 19558
rect 9612 19556 9636 19558
rect 9692 19556 9698 19558
rect 9390 19547 9698 19556
rect 5170 19068 5478 19077
rect 5170 19066 5176 19068
rect 5232 19066 5256 19068
rect 5312 19066 5336 19068
rect 5392 19066 5416 19068
rect 5472 19066 5478 19068
rect 5232 19014 5234 19066
rect 5414 19014 5416 19066
rect 5170 19012 5176 19014
rect 5232 19012 5256 19014
rect 5312 19012 5336 19014
rect 5392 19012 5416 19014
rect 5472 19012 5478 19014
rect 5170 19003 5478 19012
rect 13611 19068 13919 19077
rect 13611 19066 13617 19068
rect 13673 19066 13697 19068
rect 13753 19066 13777 19068
rect 13833 19066 13857 19068
rect 13913 19066 13919 19068
rect 13673 19014 13675 19066
rect 13855 19014 13857 19066
rect 13611 19012 13617 19014
rect 13673 19012 13697 19014
rect 13753 19012 13777 19014
rect 13833 19012 13857 19014
rect 13913 19012 13919 19014
rect 13611 19003 13919 19012
rect 9390 18524 9698 18533
rect 9390 18522 9396 18524
rect 9452 18522 9476 18524
rect 9532 18522 9556 18524
rect 9612 18522 9636 18524
rect 9692 18522 9698 18524
rect 9452 18470 9454 18522
rect 9634 18470 9636 18522
rect 9390 18468 9396 18470
rect 9452 18468 9476 18470
rect 9532 18468 9556 18470
rect 9612 18468 9636 18470
rect 9692 18468 9698 18470
rect 9390 18459 9698 18468
rect 5170 17980 5478 17989
rect 5170 17978 5176 17980
rect 5232 17978 5256 17980
rect 5312 17978 5336 17980
rect 5392 17978 5416 17980
rect 5472 17978 5478 17980
rect 5232 17926 5234 17978
rect 5414 17926 5416 17978
rect 5170 17924 5176 17926
rect 5232 17924 5256 17926
rect 5312 17924 5336 17926
rect 5392 17924 5416 17926
rect 5472 17924 5478 17926
rect 5170 17915 5478 17924
rect 13611 17980 13919 17989
rect 13611 17978 13617 17980
rect 13673 17978 13697 17980
rect 13753 17978 13777 17980
rect 13833 17978 13857 17980
rect 13913 17978 13919 17980
rect 13673 17926 13675 17978
rect 13855 17926 13857 17978
rect 13611 17924 13617 17926
rect 13673 17924 13697 17926
rect 13753 17924 13777 17926
rect 13833 17924 13857 17926
rect 13913 17924 13919 17926
rect 13611 17915 13919 17924
rect 15568 17672 15620 17678
rect 15568 17614 15620 17620
rect 9390 17436 9698 17445
rect 9390 17434 9396 17436
rect 9452 17434 9476 17436
rect 9532 17434 9556 17436
rect 9612 17434 9636 17436
rect 9692 17434 9698 17436
rect 9452 17382 9454 17434
rect 9634 17382 9636 17434
rect 9390 17380 9396 17382
rect 9452 17380 9476 17382
rect 9532 17380 9556 17382
rect 9612 17380 9636 17382
rect 9692 17380 9698 17382
rect 9390 17371 9698 17380
rect 15580 17338 15608 17614
rect 15568 17332 15620 17338
rect 15568 17274 15620 17280
rect 16040 17270 16068 22066
rect 17144 22030 17172 22066
rect 17132 22024 17184 22030
rect 17132 21966 17184 21972
rect 17144 20602 17172 21966
rect 17236 21622 17264 22170
rect 18616 22030 18644 22442
rect 18800 22030 18828 22578
rect 18892 22574 18920 24210
rect 19352 24206 19380 25366
rect 20272 25362 20300 26250
rect 20260 25356 20312 25362
rect 20260 25298 20312 25304
rect 19524 25288 19576 25294
rect 19524 25230 19576 25236
rect 20444 25288 20496 25294
rect 20444 25230 20496 25236
rect 19536 24954 19564 25230
rect 20260 25220 20312 25226
rect 20260 25162 20312 25168
rect 19524 24948 19576 24954
rect 19524 24890 19576 24896
rect 19536 24274 19564 24890
rect 19524 24268 19576 24274
rect 19524 24210 19576 24216
rect 19340 24200 19392 24206
rect 19340 24142 19392 24148
rect 20168 24064 20220 24070
rect 20168 24006 20220 24012
rect 20180 23866 20208 24006
rect 20168 23860 20220 23866
rect 20168 23802 20220 23808
rect 19800 23044 19852 23050
rect 19800 22986 19852 22992
rect 19064 22976 19116 22982
rect 19064 22918 19116 22924
rect 19076 22642 19104 22918
rect 19812 22778 19840 22986
rect 19984 22976 20036 22982
rect 19984 22918 20036 22924
rect 19800 22772 19852 22778
rect 19800 22714 19852 22720
rect 19064 22636 19116 22642
rect 19064 22578 19116 22584
rect 18880 22568 18932 22574
rect 18880 22510 18932 22516
rect 18604 22024 18656 22030
rect 18604 21966 18656 21972
rect 18788 22024 18840 22030
rect 18788 21966 18840 21972
rect 18328 21956 18380 21962
rect 18328 21898 18380 21904
rect 17684 21888 17736 21894
rect 17684 21830 17736 21836
rect 17696 21690 17724 21830
rect 17831 21788 18139 21797
rect 17831 21786 17837 21788
rect 17893 21786 17917 21788
rect 17973 21786 17997 21788
rect 18053 21786 18077 21788
rect 18133 21786 18139 21788
rect 17893 21734 17895 21786
rect 18075 21734 18077 21786
rect 17831 21732 17837 21734
rect 17893 21732 17917 21734
rect 17973 21732 17997 21734
rect 18053 21732 18077 21734
rect 18133 21732 18139 21734
rect 17831 21723 18139 21732
rect 18340 21690 18368 21898
rect 18512 21888 18564 21894
rect 18512 21830 18564 21836
rect 17684 21684 17736 21690
rect 17684 21626 17736 21632
rect 18328 21684 18380 21690
rect 18328 21626 18380 21632
rect 18524 21622 18552 21830
rect 17224 21616 17276 21622
rect 17224 21558 17276 21564
rect 18512 21616 18564 21622
rect 18512 21558 18564 21564
rect 18616 21570 18644 21966
rect 18800 21894 18828 21966
rect 18788 21888 18840 21894
rect 18788 21830 18840 21836
rect 18616 21554 18736 21570
rect 18616 21548 18748 21554
rect 18616 21542 18696 21548
rect 18696 21490 18748 21496
rect 18052 21344 18104 21350
rect 18052 21286 18104 21292
rect 18064 20942 18092 21286
rect 18892 21010 18920 22510
rect 19996 22234 20024 22918
rect 19984 22228 20036 22234
rect 19984 22170 20036 22176
rect 18972 22024 19024 22030
rect 18972 21966 19024 21972
rect 18984 21622 19012 21966
rect 19432 21956 19484 21962
rect 19432 21898 19484 21904
rect 18972 21616 19024 21622
rect 18972 21558 19024 21564
rect 19444 21554 19472 21898
rect 19892 21888 19944 21894
rect 19892 21830 19944 21836
rect 19616 21684 19668 21690
rect 19616 21626 19668 21632
rect 19432 21548 19484 21554
rect 19432 21490 19484 21496
rect 19628 21350 19656 21626
rect 19904 21554 19932 21830
rect 19708 21548 19760 21554
rect 19708 21490 19760 21496
rect 19892 21548 19944 21554
rect 19892 21490 19944 21496
rect 19616 21344 19668 21350
rect 19616 21286 19668 21292
rect 18880 21004 18932 21010
rect 18880 20946 18932 20952
rect 17684 20936 17736 20942
rect 17684 20878 17736 20884
rect 18052 20936 18104 20942
rect 18052 20878 18104 20884
rect 17592 20868 17644 20874
rect 17592 20810 17644 20816
rect 17132 20596 17184 20602
rect 17132 20538 17184 20544
rect 17604 20466 17632 20810
rect 17592 20460 17644 20466
rect 17592 20402 17644 20408
rect 17696 20330 17724 20878
rect 18236 20800 18288 20806
rect 18236 20742 18288 20748
rect 18512 20800 18564 20806
rect 18512 20742 18564 20748
rect 17831 20700 18139 20709
rect 17831 20698 17837 20700
rect 17893 20698 17917 20700
rect 17973 20698 17997 20700
rect 18053 20698 18077 20700
rect 18133 20698 18139 20700
rect 17893 20646 17895 20698
rect 18075 20646 18077 20698
rect 17831 20644 17837 20646
rect 17893 20644 17917 20646
rect 17973 20644 17997 20646
rect 18053 20644 18077 20646
rect 18133 20644 18139 20646
rect 17831 20635 18139 20644
rect 18248 20602 18276 20742
rect 17776 20596 17828 20602
rect 17776 20538 17828 20544
rect 18236 20596 18288 20602
rect 18236 20538 18288 20544
rect 17788 20380 17816 20538
rect 17960 20392 18012 20398
rect 17788 20352 17960 20380
rect 17684 20324 17736 20330
rect 17684 20266 17736 20272
rect 17696 20058 17724 20266
rect 17684 20052 17736 20058
rect 17684 19994 17736 20000
rect 17684 19848 17736 19854
rect 17788 19836 17816 20352
rect 17960 20334 18012 20340
rect 18144 20256 18196 20262
rect 18144 20198 18196 20204
rect 18156 20058 18184 20198
rect 18144 20052 18196 20058
rect 18144 19994 18196 20000
rect 17736 19808 17816 19836
rect 17684 19790 17736 19796
rect 18524 19786 18552 20742
rect 19628 20602 19656 21286
rect 19720 20602 19748 21490
rect 19800 21480 19852 21486
rect 19800 21422 19852 21428
rect 19812 21146 19840 21422
rect 19800 21140 19852 21146
rect 19800 21082 19852 21088
rect 19616 20596 19668 20602
rect 19616 20538 19668 20544
rect 19708 20596 19760 20602
rect 19708 20538 19760 20544
rect 19708 20460 19760 20466
rect 19708 20402 19760 20408
rect 19340 20256 19392 20262
rect 19340 20198 19392 20204
rect 19432 20256 19484 20262
rect 19432 20198 19484 20204
rect 19352 20058 19380 20198
rect 19340 20052 19392 20058
rect 19340 19994 19392 20000
rect 18512 19780 18564 19786
rect 18512 19722 18564 19728
rect 18696 19780 18748 19786
rect 18696 19722 18748 19728
rect 18236 19712 18288 19718
rect 18236 19654 18288 19660
rect 18328 19712 18380 19718
rect 18328 19654 18380 19660
rect 17831 19612 18139 19621
rect 17831 19610 17837 19612
rect 17893 19610 17917 19612
rect 17973 19610 17997 19612
rect 18053 19610 18077 19612
rect 18133 19610 18139 19612
rect 17893 19558 17895 19610
rect 18075 19558 18077 19610
rect 17831 19556 17837 19558
rect 17893 19556 17917 19558
rect 17973 19556 17997 19558
rect 18053 19556 18077 19558
rect 18133 19556 18139 19558
rect 17831 19547 18139 19556
rect 18248 19310 18276 19654
rect 18340 19378 18368 19654
rect 18708 19378 18736 19722
rect 19248 19712 19300 19718
rect 19248 19654 19300 19660
rect 19260 19514 19288 19654
rect 19444 19514 19472 20198
rect 19720 20058 19748 20402
rect 19708 20052 19760 20058
rect 19708 19994 19760 20000
rect 19800 19984 19852 19990
rect 19800 19926 19852 19932
rect 19248 19508 19300 19514
rect 19248 19450 19300 19456
rect 19432 19508 19484 19514
rect 19432 19450 19484 19456
rect 18328 19372 18380 19378
rect 18328 19314 18380 19320
rect 18696 19372 18748 19378
rect 18696 19314 18748 19320
rect 18972 19372 19024 19378
rect 18972 19314 19024 19320
rect 19708 19372 19760 19378
rect 19812 19360 19840 19926
rect 19760 19332 19840 19360
rect 19708 19314 19760 19320
rect 18236 19304 18288 19310
rect 18236 19246 18288 19252
rect 17132 19236 17184 19242
rect 17132 19178 17184 19184
rect 16212 18760 16264 18766
rect 16212 18702 16264 18708
rect 16224 17762 16252 18702
rect 17144 18290 17172 19178
rect 18236 19168 18288 19174
rect 18236 19110 18288 19116
rect 17224 18760 17276 18766
rect 17224 18702 17276 18708
rect 17236 18426 17264 18702
rect 17684 18624 17736 18630
rect 17684 18566 17736 18572
rect 17224 18420 17276 18426
rect 17224 18362 17276 18368
rect 17132 18284 17184 18290
rect 17132 18226 17184 18232
rect 17696 18222 17724 18566
rect 17831 18524 18139 18533
rect 17831 18522 17837 18524
rect 17893 18522 17917 18524
rect 17973 18522 17997 18524
rect 18053 18522 18077 18524
rect 18133 18522 18139 18524
rect 17893 18470 17895 18522
rect 18075 18470 18077 18522
rect 17831 18468 17837 18470
rect 17893 18468 17917 18470
rect 17973 18468 17997 18470
rect 18053 18468 18077 18470
rect 18133 18468 18139 18470
rect 17831 18459 18139 18468
rect 18248 18408 18276 19110
rect 18340 18970 18368 19314
rect 18984 18970 19012 19314
rect 19340 19304 19392 19310
rect 19340 19246 19392 19252
rect 19156 19168 19208 19174
rect 19156 19110 19208 19116
rect 18328 18964 18380 18970
rect 18328 18906 18380 18912
rect 18972 18964 19024 18970
rect 18972 18906 19024 18912
rect 18340 18426 18368 18906
rect 18984 18834 19012 18906
rect 18972 18828 19024 18834
rect 18972 18770 19024 18776
rect 19168 18766 19196 19110
rect 19352 18766 19380 19246
rect 19720 18970 19748 19314
rect 19708 18964 19760 18970
rect 19708 18906 19760 18912
rect 19156 18760 19208 18766
rect 19156 18702 19208 18708
rect 19340 18760 19392 18766
rect 19340 18702 19392 18708
rect 19616 18760 19668 18766
rect 19616 18702 19668 18708
rect 19800 18760 19852 18766
rect 19996 18714 20024 22170
rect 20272 21622 20300 25162
rect 20352 25152 20404 25158
rect 20352 25094 20404 25100
rect 20364 24682 20392 25094
rect 20456 24954 20484 25230
rect 20548 24954 20576 26318
rect 20904 26318 20956 26324
rect 20626 26279 20682 26288
rect 20444 24948 20496 24954
rect 20444 24890 20496 24896
rect 20536 24948 20588 24954
rect 20536 24890 20588 24896
rect 20352 24676 20404 24682
rect 20352 24618 20404 24624
rect 20640 24188 20668 26279
rect 20916 26042 20944 26318
rect 20904 26036 20956 26042
rect 20904 25978 20956 25984
rect 21008 25838 21036 27474
rect 21088 27464 21140 27470
rect 21088 27406 21140 27412
rect 21100 27130 21128 27406
rect 21088 27124 21140 27130
rect 21088 27066 21140 27072
rect 21272 27124 21324 27130
rect 21272 27066 21324 27072
rect 21284 27033 21312 27066
rect 21270 27024 21326 27033
rect 21180 26988 21232 26994
rect 21270 26959 21326 26968
rect 21364 26988 21416 26994
rect 21180 26930 21232 26936
rect 21364 26930 21416 26936
rect 21192 26790 21220 26930
rect 21272 26920 21324 26926
rect 21376 26897 21404 26930
rect 21272 26862 21324 26868
rect 21362 26888 21418 26897
rect 21088 26784 21140 26790
rect 21088 26726 21140 26732
rect 21180 26784 21232 26790
rect 21180 26726 21232 26732
rect 21100 26518 21128 26726
rect 21088 26512 21140 26518
rect 21088 26454 21140 26460
rect 21192 25974 21220 26726
rect 21284 26382 21312 26862
rect 21362 26823 21418 26832
rect 21732 26784 21784 26790
rect 21732 26726 21784 26732
rect 21744 26382 21772 26726
rect 21272 26376 21324 26382
rect 21364 26376 21416 26382
rect 21272 26318 21324 26324
rect 21362 26344 21364 26353
rect 21732 26376 21784 26382
rect 21416 26344 21418 26353
rect 21732 26318 21784 26324
rect 21836 26314 21864 27610
rect 22468 26988 22520 26994
rect 22468 26930 22520 26936
rect 22052 26684 22360 26693
rect 22052 26682 22058 26684
rect 22114 26682 22138 26684
rect 22194 26682 22218 26684
rect 22274 26682 22298 26684
rect 22354 26682 22360 26684
rect 22114 26630 22116 26682
rect 22296 26630 22298 26682
rect 22052 26628 22058 26630
rect 22114 26628 22138 26630
rect 22194 26628 22218 26630
rect 22274 26628 22298 26630
rect 22354 26628 22360 26630
rect 22052 26619 22360 26628
rect 22480 26586 22508 26930
rect 22836 26784 22888 26790
rect 22836 26726 22888 26732
rect 22468 26580 22520 26586
rect 22468 26522 22520 26528
rect 21916 26512 21968 26518
rect 21914 26480 21916 26489
rect 21968 26480 21970 26489
rect 21914 26415 21970 26424
rect 22848 26382 22876 26726
rect 22836 26376 22888 26382
rect 22836 26318 22888 26324
rect 21362 26279 21418 26288
rect 21824 26308 21876 26314
rect 22468 26308 22520 26314
rect 21876 26268 21956 26296
rect 21824 26250 21876 26256
rect 21272 26240 21324 26246
rect 21272 26182 21324 26188
rect 21180 25968 21232 25974
rect 21180 25910 21232 25916
rect 20996 25832 21048 25838
rect 20996 25774 21048 25780
rect 21284 25430 21312 26182
rect 21456 25900 21508 25906
rect 21456 25842 21508 25848
rect 20904 25424 20956 25430
rect 20904 25366 20956 25372
rect 20996 25424 21048 25430
rect 20996 25366 21048 25372
rect 21272 25424 21324 25430
rect 21272 25366 21324 25372
rect 20720 25152 20772 25158
rect 20720 25094 20772 25100
rect 20732 24750 20760 25094
rect 20720 24744 20772 24750
rect 20720 24686 20772 24692
rect 20916 24206 20944 25366
rect 21008 25226 21036 25366
rect 21468 25226 21496 25842
rect 21548 25832 21600 25838
rect 21548 25774 21600 25780
rect 20996 25220 21048 25226
rect 20996 25162 21048 25168
rect 21456 25220 21508 25226
rect 21456 25162 21508 25168
rect 20720 24200 20772 24206
rect 20640 24160 20720 24188
rect 20720 24142 20772 24148
rect 20904 24200 20956 24206
rect 20904 24142 20956 24148
rect 20732 23118 20760 24142
rect 21008 24070 21036 25162
rect 21272 25152 21324 25158
rect 21272 25094 21324 25100
rect 21284 24614 21312 25094
rect 21560 24818 21588 25774
rect 21824 25288 21876 25294
rect 21824 25230 21876 25236
rect 21548 24812 21600 24818
rect 21548 24754 21600 24760
rect 21088 24608 21140 24614
rect 21088 24550 21140 24556
rect 21272 24608 21324 24614
rect 21272 24550 21324 24556
rect 21100 24410 21128 24550
rect 21560 24410 21588 24754
rect 21088 24404 21140 24410
rect 21088 24346 21140 24352
rect 21548 24404 21600 24410
rect 21548 24346 21600 24352
rect 20996 24064 21048 24070
rect 20996 24006 21048 24012
rect 21456 24064 21508 24070
rect 21456 24006 21508 24012
rect 21468 23866 21496 24006
rect 21456 23860 21508 23866
rect 21456 23802 21508 23808
rect 20628 23112 20680 23118
rect 20628 23054 20680 23060
rect 20720 23112 20772 23118
rect 20720 23054 20772 23060
rect 20904 23112 20956 23118
rect 20904 23054 20956 23060
rect 21732 23112 21784 23118
rect 21732 23054 21784 23060
rect 20640 22234 20668 23054
rect 20812 22432 20864 22438
rect 20812 22374 20864 22380
rect 20628 22228 20680 22234
rect 20628 22170 20680 22176
rect 20352 21956 20404 21962
rect 20352 21898 20404 21904
rect 20364 21690 20392 21898
rect 20720 21888 20772 21894
rect 20720 21830 20772 21836
rect 20352 21684 20404 21690
rect 20352 21626 20404 21632
rect 20260 21616 20312 21622
rect 20260 21558 20312 21564
rect 20732 21486 20760 21830
rect 20720 21480 20772 21486
rect 20720 21422 20772 21428
rect 20260 21344 20312 21350
rect 20260 21286 20312 21292
rect 20444 21344 20496 21350
rect 20444 21286 20496 21292
rect 20272 20466 20300 21286
rect 20456 21146 20484 21286
rect 20444 21140 20496 21146
rect 20444 21082 20496 21088
rect 20732 21010 20760 21422
rect 20824 21350 20852 22374
rect 20812 21344 20864 21350
rect 20812 21286 20864 21292
rect 20720 21004 20772 21010
rect 20720 20946 20772 20952
rect 20260 20460 20312 20466
rect 20260 20402 20312 20408
rect 20076 19848 20128 19854
rect 20076 19790 20128 19796
rect 20088 19514 20116 19790
rect 20720 19712 20772 19718
rect 20720 19654 20772 19660
rect 20076 19508 20128 19514
rect 20076 19450 20128 19456
rect 20168 19372 20220 19378
rect 20168 19314 20220 19320
rect 20180 18970 20208 19314
rect 20168 18964 20220 18970
rect 20168 18906 20220 18912
rect 20536 18964 20588 18970
rect 20536 18906 20588 18912
rect 20548 18766 20576 18906
rect 20732 18766 20760 19654
rect 20824 18970 20852 21286
rect 20916 19446 20944 23054
rect 21744 22778 21772 23054
rect 21836 22982 21864 25230
rect 21928 24954 21956 26268
rect 22468 26250 22520 26256
rect 22052 25596 22360 25605
rect 22052 25594 22058 25596
rect 22114 25594 22138 25596
rect 22194 25594 22218 25596
rect 22274 25594 22298 25596
rect 22354 25594 22360 25596
rect 22114 25542 22116 25594
rect 22296 25542 22298 25594
rect 22052 25540 22058 25542
rect 22114 25540 22138 25542
rect 22194 25540 22218 25542
rect 22274 25540 22298 25542
rect 22354 25540 22360 25542
rect 22052 25531 22360 25540
rect 22480 25294 22508 26250
rect 22848 25906 22876 26318
rect 22744 25900 22796 25906
rect 22744 25842 22796 25848
rect 22836 25900 22888 25906
rect 22836 25842 22888 25848
rect 22756 25498 22784 25842
rect 22744 25492 22796 25498
rect 22744 25434 22796 25440
rect 22468 25288 22520 25294
rect 22468 25230 22520 25236
rect 22744 25220 22796 25226
rect 22744 25162 22796 25168
rect 21916 24948 21968 24954
rect 21916 24890 21968 24896
rect 21928 24342 21956 24890
rect 22560 24812 22612 24818
rect 22560 24754 22612 24760
rect 22052 24508 22360 24517
rect 22052 24506 22058 24508
rect 22114 24506 22138 24508
rect 22194 24506 22218 24508
rect 22274 24506 22298 24508
rect 22354 24506 22360 24508
rect 22114 24454 22116 24506
rect 22296 24454 22298 24506
rect 22052 24452 22058 24454
rect 22114 24452 22138 24454
rect 22194 24452 22218 24454
rect 22274 24452 22298 24454
rect 22354 24452 22360 24454
rect 22052 24443 22360 24452
rect 22572 24410 22600 24754
rect 22652 24608 22704 24614
rect 22652 24550 22704 24556
rect 22560 24404 22612 24410
rect 22560 24346 22612 24352
rect 22664 24342 22692 24550
rect 22756 24410 22784 25162
rect 22744 24404 22796 24410
rect 22744 24346 22796 24352
rect 21916 24336 21968 24342
rect 21916 24278 21968 24284
rect 22652 24336 22704 24342
rect 22652 24278 22704 24284
rect 22928 24200 22980 24206
rect 22928 24142 22980 24148
rect 22744 24064 22796 24070
rect 22744 24006 22796 24012
rect 22756 23866 22784 24006
rect 22744 23860 22796 23866
rect 22744 23802 22796 23808
rect 22940 23798 22968 24142
rect 22928 23792 22980 23798
rect 22928 23734 22980 23740
rect 22376 23724 22428 23730
rect 22376 23666 22428 23672
rect 22052 23420 22360 23429
rect 22052 23418 22058 23420
rect 22114 23418 22138 23420
rect 22194 23418 22218 23420
rect 22274 23418 22298 23420
rect 22354 23418 22360 23420
rect 22114 23366 22116 23418
rect 22296 23366 22298 23418
rect 22052 23364 22058 23366
rect 22114 23364 22138 23366
rect 22194 23364 22218 23366
rect 22274 23364 22298 23366
rect 22354 23364 22360 23366
rect 22052 23355 22360 23364
rect 22388 23322 22416 23666
rect 22928 23520 22980 23526
rect 22928 23462 22980 23468
rect 22376 23316 22428 23322
rect 22376 23258 22428 23264
rect 22376 23044 22428 23050
rect 22376 22986 22428 22992
rect 21824 22976 21876 22982
rect 21824 22918 21876 22924
rect 21732 22772 21784 22778
rect 21732 22714 21784 22720
rect 22388 22710 22416 22986
rect 22376 22704 22428 22710
rect 22376 22646 22428 22652
rect 22940 22642 22968 23462
rect 23032 22778 23060 28494
rect 23112 28416 23164 28422
rect 23112 28358 23164 28364
rect 23204 28416 23256 28422
rect 23204 28358 23256 28364
rect 23124 27470 23152 28358
rect 23112 27464 23164 27470
rect 23112 27406 23164 27412
rect 23216 26994 23244 28358
rect 23308 28082 23336 31282
rect 23400 30938 23428 31418
rect 23388 30932 23440 30938
rect 23388 30874 23440 30880
rect 23400 30394 23428 30874
rect 23664 30728 23716 30734
rect 23664 30670 23716 30676
rect 23848 30728 23900 30734
rect 23848 30670 23900 30676
rect 23480 30592 23532 30598
rect 23480 30534 23532 30540
rect 23572 30592 23624 30598
rect 23572 30534 23624 30540
rect 23388 30388 23440 30394
rect 23388 30330 23440 30336
rect 23388 30252 23440 30258
rect 23388 30194 23440 30200
rect 23400 29850 23428 30194
rect 23492 29850 23520 30534
rect 23388 29844 23440 29850
rect 23388 29786 23440 29792
rect 23480 29844 23532 29850
rect 23480 29786 23532 29792
rect 23492 29170 23520 29786
rect 23584 29646 23612 30534
rect 23676 29714 23704 30670
rect 23664 29708 23716 29714
rect 23664 29650 23716 29656
rect 23572 29640 23624 29646
rect 23572 29582 23624 29588
rect 23480 29164 23532 29170
rect 23480 29106 23532 29112
rect 23676 28762 23704 29650
rect 23860 29238 23888 30670
rect 23848 29232 23900 29238
rect 23848 29174 23900 29180
rect 23664 28756 23716 28762
rect 23664 28698 23716 28704
rect 23848 28416 23900 28422
rect 23848 28358 23900 28364
rect 23664 28212 23716 28218
rect 23664 28154 23716 28160
rect 23296 28076 23348 28082
rect 23296 28018 23348 28024
rect 23572 28076 23624 28082
rect 23572 28018 23624 28024
rect 23584 27130 23612 28018
rect 23676 27470 23704 28154
rect 23860 27614 23888 28358
rect 23768 27606 23888 27614
rect 23756 27600 23888 27606
rect 23808 27586 23888 27600
rect 23756 27542 23808 27548
rect 23664 27464 23716 27470
rect 23664 27406 23716 27412
rect 23768 27334 23796 27542
rect 23756 27328 23808 27334
rect 23756 27270 23808 27276
rect 23572 27124 23624 27130
rect 23572 27066 23624 27072
rect 23204 26988 23256 26994
rect 23204 26930 23256 26936
rect 23216 26858 23244 26930
rect 23204 26852 23256 26858
rect 23204 26794 23256 26800
rect 23768 26586 23796 27270
rect 23756 26580 23808 26586
rect 23756 26522 23808 26528
rect 23480 26308 23532 26314
rect 23480 26250 23532 26256
rect 23492 25838 23520 26250
rect 23572 26240 23624 26246
rect 23572 26182 23624 26188
rect 23584 25906 23612 26182
rect 23572 25900 23624 25906
rect 23572 25842 23624 25848
rect 23480 25832 23532 25838
rect 23480 25774 23532 25780
rect 23584 25702 23612 25842
rect 23572 25696 23624 25702
rect 23572 25638 23624 25644
rect 23584 25226 23612 25638
rect 23952 25362 23980 31758
rect 25516 31754 25544 32166
rect 25424 31726 25544 31754
rect 24492 31408 24544 31414
rect 24492 31350 24544 31356
rect 24504 30870 24532 31350
rect 24676 31136 24728 31142
rect 24676 31078 24728 31084
rect 24768 31136 24820 31142
rect 24768 31078 24820 31084
rect 24688 30938 24716 31078
rect 24676 30932 24728 30938
rect 24676 30874 24728 30880
rect 24492 30864 24544 30870
rect 24492 30806 24544 30812
rect 24780 30734 24808 31078
rect 25424 30734 25452 31726
rect 25504 31136 25556 31142
rect 25504 31078 25556 31084
rect 25516 30938 25544 31078
rect 25504 30932 25556 30938
rect 25504 30874 25556 30880
rect 24216 30728 24268 30734
rect 24216 30670 24268 30676
rect 24768 30728 24820 30734
rect 24768 30670 24820 30676
rect 25412 30728 25464 30734
rect 25412 30670 25464 30676
rect 25596 30728 25648 30734
rect 25596 30670 25648 30676
rect 24032 30252 24084 30258
rect 24032 30194 24084 30200
rect 24044 29850 24072 30194
rect 24228 29850 24256 30670
rect 24308 30660 24360 30666
rect 24308 30602 24360 30608
rect 24952 30660 25004 30666
rect 24952 30602 25004 30608
rect 24032 29844 24084 29850
rect 24032 29786 24084 29792
rect 24216 29844 24268 29850
rect 24216 29786 24268 29792
rect 24032 28484 24084 28490
rect 24032 28426 24084 28432
rect 24044 28218 24072 28426
rect 24032 28212 24084 28218
rect 24032 28154 24084 28160
rect 24032 28076 24084 28082
rect 24032 28018 24084 28024
rect 24044 27674 24072 28018
rect 24032 27668 24084 27674
rect 24032 27610 24084 27616
rect 24124 27396 24176 27402
rect 24124 27338 24176 27344
rect 24136 27062 24164 27338
rect 24124 27056 24176 27062
rect 24124 26998 24176 27004
rect 24216 26240 24268 26246
rect 24216 26182 24268 26188
rect 24228 25974 24256 26182
rect 24320 25974 24348 30602
rect 24964 30190 24992 30602
rect 25608 30258 25636 30670
rect 25700 30598 25728 32710
rect 25884 32570 25912 32710
rect 25976 32570 26004 32830
rect 26068 32852 26240 32858
rect 26068 32846 26292 32852
rect 26068 32830 26280 32846
rect 25780 32564 25832 32570
rect 25780 32506 25832 32512
rect 25872 32564 25924 32570
rect 25872 32506 25924 32512
rect 25964 32564 26016 32570
rect 25964 32506 26016 32512
rect 25792 32298 25820 32506
rect 25872 32360 25924 32366
rect 25872 32302 25924 32308
rect 25780 32292 25832 32298
rect 25780 32234 25832 32240
rect 25884 31890 25912 32302
rect 26068 31958 26096 32830
rect 26148 32768 26200 32774
rect 26148 32710 26200 32716
rect 26056 31952 26108 31958
rect 26056 31894 26108 31900
rect 26160 31890 26188 32710
rect 26272 32668 26580 32677
rect 26272 32666 26278 32668
rect 26334 32666 26358 32668
rect 26414 32666 26438 32668
rect 26494 32666 26518 32668
rect 26574 32666 26580 32668
rect 26334 32614 26336 32666
rect 26516 32614 26518 32666
rect 26272 32612 26278 32614
rect 26334 32612 26358 32614
rect 26414 32612 26438 32614
rect 26494 32612 26518 32614
rect 26574 32612 26580 32614
rect 26272 32603 26580 32612
rect 26620 32502 26648 33390
rect 26896 32502 26924 33866
rect 26976 33516 27028 33522
rect 26976 33458 27028 33464
rect 29552 33516 29604 33522
rect 29552 33458 29604 33464
rect 30196 33516 30248 33522
rect 30196 33458 30248 33464
rect 30288 33516 30340 33522
rect 30288 33458 30340 33464
rect 31024 33516 31076 33522
rect 31024 33458 31076 33464
rect 32220 33516 32272 33522
rect 32220 33458 32272 33464
rect 26988 33046 27016 33458
rect 27068 33448 27120 33454
rect 27068 33390 27120 33396
rect 27252 33448 27304 33454
rect 27252 33390 27304 33396
rect 28356 33448 28408 33454
rect 28356 33390 28408 33396
rect 26976 33040 27028 33046
rect 26976 32982 27028 32988
rect 26988 32570 27016 32982
rect 27080 32774 27108 33390
rect 27160 33312 27212 33318
rect 27160 33254 27212 33260
rect 27172 32978 27200 33254
rect 27264 33114 27292 33390
rect 27436 33380 27488 33386
rect 27436 33322 27488 33328
rect 27252 33108 27304 33114
rect 27252 33050 27304 33056
rect 27160 32972 27212 32978
rect 27160 32914 27212 32920
rect 27068 32768 27120 32774
rect 27068 32710 27120 32716
rect 26976 32564 27028 32570
rect 26976 32506 27028 32512
rect 26608 32496 26660 32502
rect 26608 32438 26660 32444
rect 26884 32496 26936 32502
rect 26884 32438 26936 32444
rect 26240 32360 26292 32366
rect 26240 32302 26292 32308
rect 25872 31884 25924 31890
rect 25872 31826 25924 31832
rect 26148 31884 26200 31890
rect 26148 31826 26200 31832
rect 26252 31668 26280 32302
rect 26700 32224 26752 32230
rect 26700 32166 26752 32172
rect 26712 31890 26740 32166
rect 26700 31884 26752 31890
rect 26700 31826 26752 31832
rect 26160 31640 26280 31668
rect 25780 30728 25832 30734
rect 25780 30670 25832 30676
rect 25688 30592 25740 30598
rect 25688 30534 25740 30540
rect 25700 30258 25728 30534
rect 25792 30394 25820 30670
rect 25780 30388 25832 30394
rect 25780 30330 25832 30336
rect 26160 30274 26188 31640
rect 26272 31580 26580 31589
rect 26272 31578 26278 31580
rect 26334 31578 26358 31580
rect 26414 31578 26438 31580
rect 26494 31578 26518 31580
rect 26574 31578 26580 31580
rect 26334 31526 26336 31578
rect 26516 31526 26518 31578
rect 26272 31524 26278 31526
rect 26334 31524 26358 31526
rect 26414 31524 26438 31526
rect 26494 31524 26518 31526
rect 26574 31524 26580 31526
rect 26272 31515 26580 31524
rect 26896 30802 26924 32438
rect 27080 32026 27108 32710
rect 27172 32570 27200 32914
rect 27344 32904 27396 32910
rect 27344 32846 27396 32852
rect 27160 32564 27212 32570
rect 27160 32506 27212 32512
rect 27356 32416 27384 32846
rect 27448 32570 27476 33322
rect 28368 32570 28396 33390
rect 29564 33114 29592 33458
rect 30012 33448 30064 33454
rect 30012 33390 30064 33396
rect 29920 33312 29972 33318
rect 29920 33254 29972 33260
rect 29552 33108 29604 33114
rect 29552 33050 29604 33056
rect 29932 32910 29960 33254
rect 29736 32904 29788 32910
rect 29736 32846 29788 32852
rect 29920 32904 29972 32910
rect 29920 32846 29972 32852
rect 28908 32768 28960 32774
rect 28908 32710 28960 32716
rect 29092 32768 29144 32774
rect 29092 32710 29144 32716
rect 27436 32564 27488 32570
rect 27436 32506 27488 32512
rect 28356 32564 28408 32570
rect 28356 32506 28408 32512
rect 27436 32428 27488 32434
rect 27356 32388 27436 32416
rect 27068 32020 27120 32026
rect 27068 31962 27120 31968
rect 27356 30938 27384 32388
rect 27436 32370 27488 32376
rect 27620 31884 27672 31890
rect 27620 31826 27672 31832
rect 27436 31340 27488 31346
rect 27436 31282 27488 31288
rect 27344 30932 27396 30938
rect 27344 30874 27396 30880
rect 26884 30796 26936 30802
rect 26884 30738 26936 30744
rect 26608 30728 26660 30734
rect 26608 30670 26660 30676
rect 26272 30492 26580 30501
rect 26272 30490 26278 30492
rect 26334 30490 26358 30492
rect 26414 30490 26438 30492
rect 26494 30490 26518 30492
rect 26574 30490 26580 30492
rect 26334 30438 26336 30490
rect 26516 30438 26518 30490
rect 26272 30436 26278 30438
rect 26334 30436 26358 30438
rect 26414 30436 26438 30438
rect 26494 30436 26518 30438
rect 26574 30436 26580 30438
rect 26272 30427 26580 30436
rect 26620 30394 26648 30670
rect 26896 30598 26924 30738
rect 27448 30734 27476 31282
rect 27436 30728 27488 30734
rect 27436 30670 27488 30676
rect 27528 30728 27580 30734
rect 27528 30670 27580 30676
rect 26884 30592 26936 30598
rect 26884 30534 26936 30540
rect 27540 30394 27568 30670
rect 26608 30388 26660 30394
rect 26608 30330 26660 30336
rect 27528 30388 27580 30394
rect 27528 30330 27580 30336
rect 26160 30258 26372 30274
rect 26620 30258 26648 30330
rect 27540 30258 27568 30330
rect 27632 30258 27660 31826
rect 28920 31822 28948 32710
rect 29104 32434 29132 32710
rect 29460 32496 29512 32502
rect 29460 32438 29512 32444
rect 29092 32428 29144 32434
rect 29092 32370 29144 32376
rect 29472 32298 29500 32438
rect 29460 32292 29512 32298
rect 29460 32234 29512 32240
rect 29472 31890 29500 32234
rect 29748 32026 29776 32846
rect 29932 32570 29960 32846
rect 30024 32774 30052 33390
rect 30104 33312 30156 33318
rect 30104 33254 30156 33260
rect 30012 32768 30064 32774
rect 30012 32710 30064 32716
rect 29920 32564 29972 32570
rect 29920 32506 29972 32512
rect 30024 32434 30052 32710
rect 30116 32570 30144 33254
rect 30104 32564 30156 32570
rect 30104 32506 30156 32512
rect 30208 32502 30236 33458
rect 30300 32842 30328 33458
rect 30380 33312 30432 33318
rect 30380 33254 30432 33260
rect 30840 33312 30892 33318
rect 30840 33254 30892 33260
rect 30288 32836 30340 32842
rect 30288 32778 30340 32784
rect 30196 32496 30248 32502
rect 30196 32438 30248 32444
rect 30012 32428 30064 32434
rect 30012 32370 30064 32376
rect 29736 32020 29788 32026
rect 29736 31962 29788 31968
rect 30024 31890 30052 32370
rect 29460 31884 29512 31890
rect 29460 31826 29512 31832
rect 30012 31884 30064 31890
rect 30012 31826 30064 31832
rect 28908 31816 28960 31822
rect 28908 31758 28960 31764
rect 30288 31680 30340 31686
rect 30288 31622 30340 31628
rect 30300 31482 30328 31622
rect 30288 31476 30340 31482
rect 30288 31418 30340 31424
rect 28816 31340 28868 31346
rect 28816 31282 28868 31288
rect 27988 31136 28040 31142
rect 27988 31078 28040 31084
rect 28080 31136 28132 31142
rect 28080 31078 28132 31084
rect 28000 30870 28028 31078
rect 27988 30864 28040 30870
rect 27988 30806 28040 30812
rect 27712 30728 27764 30734
rect 27712 30670 27764 30676
rect 27804 30728 27856 30734
rect 27804 30670 27856 30676
rect 25136 30252 25188 30258
rect 25136 30194 25188 30200
rect 25320 30252 25372 30258
rect 25320 30194 25372 30200
rect 25596 30252 25648 30258
rect 25596 30194 25648 30200
rect 25688 30252 25740 30258
rect 26160 30252 26384 30258
rect 26160 30246 26332 30252
rect 25688 30194 25740 30200
rect 26332 30194 26384 30200
rect 26608 30252 26660 30258
rect 26608 30194 26660 30200
rect 27528 30252 27580 30258
rect 27528 30194 27580 30200
rect 27620 30252 27672 30258
rect 27620 30194 27672 30200
rect 24952 30184 25004 30190
rect 24952 30126 25004 30132
rect 24676 30048 24728 30054
rect 24676 29990 24728 29996
rect 24688 29850 24716 29990
rect 24964 29850 24992 30126
rect 25148 29850 25176 30194
rect 25332 29850 25360 30194
rect 24676 29844 24728 29850
rect 24676 29786 24728 29792
rect 24952 29844 25004 29850
rect 24952 29786 25004 29792
rect 25136 29844 25188 29850
rect 25136 29786 25188 29792
rect 25320 29844 25372 29850
rect 25320 29786 25372 29792
rect 25504 29572 25556 29578
rect 25504 29514 25556 29520
rect 25044 29164 25096 29170
rect 25044 29106 25096 29112
rect 25056 28694 25084 29106
rect 25136 28960 25188 28966
rect 25136 28902 25188 28908
rect 25148 28694 25176 28902
rect 25044 28688 25096 28694
rect 25044 28630 25096 28636
rect 25136 28688 25188 28694
rect 25136 28630 25188 28636
rect 25056 28218 25084 28630
rect 25516 28626 25544 29514
rect 25504 28620 25556 28626
rect 25504 28562 25556 28568
rect 25136 28552 25188 28558
rect 25136 28494 25188 28500
rect 25320 28552 25372 28558
rect 25320 28494 25372 28500
rect 25044 28212 25096 28218
rect 25044 28154 25096 28160
rect 25056 27674 25084 28154
rect 25148 27674 25176 28494
rect 25044 27668 25096 27674
rect 25044 27610 25096 27616
rect 25136 27668 25188 27674
rect 25136 27610 25188 27616
rect 25332 27470 25360 28494
rect 25504 28484 25556 28490
rect 25504 28426 25556 28432
rect 25516 28218 25544 28426
rect 25504 28212 25556 28218
rect 25504 28154 25556 28160
rect 25412 28008 25464 28014
rect 25412 27950 25464 27956
rect 25320 27464 25372 27470
rect 25320 27406 25372 27412
rect 24768 27396 24820 27402
rect 24768 27338 24820 27344
rect 24952 27396 25004 27402
rect 24952 27338 25004 27344
rect 24780 27130 24808 27338
rect 24768 27124 24820 27130
rect 24768 27066 24820 27072
rect 24492 27056 24544 27062
rect 24492 26998 24544 27004
rect 24216 25968 24268 25974
rect 24216 25910 24268 25916
rect 24308 25968 24360 25974
rect 24308 25910 24360 25916
rect 23940 25356 23992 25362
rect 23940 25298 23992 25304
rect 23572 25220 23624 25226
rect 23572 25162 23624 25168
rect 23756 25152 23808 25158
rect 23756 25094 23808 25100
rect 23768 24954 23796 25094
rect 23756 24948 23808 24954
rect 23756 24890 23808 24896
rect 23112 24608 23164 24614
rect 23112 24550 23164 24556
rect 23204 24608 23256 24614
rect 23204 24550 23256 24556
rect 24308 24608 24360 24614
rect 24308 24550 24360 24556
rect 23124 24410 23152 24550
rect 23112 24404 23164 24410
rect 23112 24346 23164 24352
rect 23112 24064 23164 24070
rect 23112 24006 23164 24012
rect 23124 23322 23152 24006
rect 23216 23866 23244 24550
rect 24320 24410 24348 24550
rect 24308 24404 24360 24410
rect 24308 24346 24360 24352
rect 23572 24200 23624 24206
rect 23572 24142 23624 24148
rect 23848 24200 23900 24206
rect 23848 24142 23900 24148
rect 23584 23866 23612 24142
rect 23204 23860 23256 23866
rect 23204 23802 23256 23808
rect 23572 23860 23624 23866
rect 23572 23802 23624 23808
rect 23388 23588 23440 23594
rect 23388 23530 23440 23536
rect 23296 23520 23348 23526
rect 23296 23462 23348 23468
rect 23112 23316 23164 23322
rect 23112 23258 23164 23264
rect 23308 23118 23336 23462
rect 23296 23112 23348 23118
rect 23296 23054 23348 23060
rect 23400 22794 23428 23530
rect 23584 23322 23612 23802
rect 23664 23656 23716 23662
rect 23664 23598 23716 23604
rect 23676 23338 23704 23598
rect 23572 23316 23624 23322
rect 23676 23310 23796 23338
rect 23572 23258 23624 23264
rect 23768 23254 23796 23310
rect 23756 23248 23808 23254
rect 23756 23190 23808 23196
rect 23768 23118 23796 23190
rect 23860 23186 23888 24142
rect 24124 24064 24176 24070
rect 24124 24006 24176 24012
rect 23848 23180 23900 23186
rect 23848 23122 23900 23128
rect 24136 23118 24164 24006
rect 24504 23730 24532 26998
rect 24964 26994 24992 27338
rect 24768 26988 24820 26994
rect 24768 26930 24820 26936
rect 24952 26988 25004 26994
rect 24952 26930 25004 26936
rect 25320 26988 25372 26994
rect 25320 26930 25372 26936
rect 24584 26580 24636 26586
rect 24584 26522 24636 26528
rect 24596 26042 24624 26522
rect 24780 26314 24808 26930
rect 25332 26586 25360 26930
rect 25320 26580 25372 26586
rect 25320 26522 25372 26528
rect 24768 26308 24820 26314
rect 24768 26250 24820 26256
rect 24952 26240 25004 26246
rect 24952 26182 25004 26188
rect 24584 26036 24636 26042
rect 24584 25978 24636 25984
rect 24676 25900 24728 25906
rect 24676 25842 24728 25848
rect 24688 25498 24716 25842
rect 24860 25696 24912 25702
rect 24964 25684 24992 26182
rect 25044 25968 25096 25974
rect 25044 25910 25096 25916
rect 24912 25656 24992 25684
rect 24860 25638 24912 25644
rect 24676 25492 24728 25498
rect 24676 25434 24728 25440
rect 24964 25430 24992 25656
rect 24952 25424 25004 25430
rect 24952 25366 25004 25372
rect 25056 24954 25084 25910
rect 25424 25906 25452 27950
rect 25516 27470 25544 28154
rect 25504 27464 25556 27470
rect 25504 27406 25556 27412
rect 25504 26988 25556 26994
rect 25504 26930 25556 26936
rect 25516 26586 25544 26930
rect 25504 26580 25556 26586
rect 25504 26522 25556 26528
rect 25608 26353 25636 30194
rect 26620 29850 26648 30194
rect 26884 30184 26936 30190
rect 26884 30126 26936 30132
rect 26700 30048 26752 30054
rect 26700 29990 26752 29996
rect 26608 29844 26660 29850
rect 26608 29786 26660 29792
rect 26712 29646 26740 29990
rect 25688 29640 25740 29646
rect 25688 29582 25740 29588
rect 25780 29640 25832 29646
rect 25780 29582 25832 29588
rect 26700 29640 26752 29646
rect 26700 29582 26752 29588
rect 25700 28558 25728 29582
rect 25792 28762 25820 29582
rect 26272 29404 26580 29413
rect 26272 29402 26278 29404
rect 26334 29402 26358 29404
rect 26414 29402 26438 29404
rect 26494 29402 26518 29404
rect 26574 29402 26580 29404
rect 26334 29350 26336 29402
rect 26516 29350 26518 29402
rect 26272 29348 26278 29350
rect 26334 29348 26358 29350
rect 26414 29348 26438 29350
rect 26494 29348 26518 29350
rect 26574 29348 26580 29350
rect 26272 29339 26580 29348
rect 26896 29306 26924 30126
rect 27436 30048 27488 30054
rect 27436 29990 27488 29996
rect 27448 29646 27476 29990
rect 27436 29640 27488 29646
rect 27436 29582 27488 29588
rect 26884 29300 26936 29306
rect 26884 29242 26936 29248
rect 26896 28994 26924 29242
rect 26896 28966 27016 28994
rect 25780 28756 25832 28762
rect 25780 28698 25832 28704
rect 25688 28552 25740 28558
rect 25688 28494 25740 28500
rect 26272 28316 26580 28325
rect 26272 28314 26278 28316
rect 26334 28314 26358 28316
rect 26414 28314 26438 28316
rect 26494 28314 26518 28316
rect 26574 28314 26580 28316
rect 26334 28262 26336 28314
rect 26516 28262 26518 28314
rect 26272 28260 26278 28262
rect 26334 28260 26358 28262
rect 26414 28260 26438 28262
rect 26494 28260 26518 28262
rect 26574 28260 26580 28262
rect 26272 28251 26580 28260
rect 25964 28076 26016 28082
rect 25964 28018 26016 28024
rect 25976 27674 26004 28018
rect 25964 27668 26016 27674
rect 25964 27610 26016 27616
rect 26988 27470 27016 28966
rect 27632 28948 27660 30194
rect 27724 29850 27752 30670
rect 27816 30258 27844 30670
rect 27896 30592 27948 30598
rect 27896 30534 27948 30540
rect 27908 30258 27936 30534
rect 28092 30258 28120 31078
rect 28172 30796 28224 30802
rect 28172 30738 28224 30744
rect 28184 30598 28212 30738
rect 28828 30734 28856 31282
rect 30392 31210 30420 33254
rect 30493 33212 30801 33221
rect 30493 33210 30499 33212
rect 30555 33210 30579 33212
rect 30635 33210 30659 33212
rect 30715 33210 30739 33212
rect 30795 33210 30801 33212
rect 30555 33158 30557 33210
rect 30737 33158 30739 33210
rect 30493 33156 30499 33158
rect 30555 33156 30579 33158
rect 30635 33156 30659 33158
rect 30715 33156 30739 33158
rect 30795 33156 30801 33158
rect 30493 33147 30801 33156
rect 30852 32502 30880 33254
rect 30840 32496 30892 32502
rect 30840 32438 30892 32444
rect 30493 32124 30801 32133
rect 30493 32122 30499 32124
rect 30555 32122 30579 32124
rect 30635 32122 30659 32124
rect 30715 32122 30739 32124
rect 30795 32122 30801 32124
rect 30555 32070 30557 32122
rect 30737 32070 30739 32122
rect 30493 32068 30499 32070
rect 30555 32068 30579 32070
rect 30635 32068 30659 32070
rect 30715 32068 30739 32070
rect 30795 32068 30801 32070
rect 30493 32059 30801 32068
rect 31036 32026 31064 33458
rect 31300 33380 31352 33386
rect 31300 33322 31352 33328
rect 31312 32910 31340 33322
rect 31208 32904 31260 32910
rect 31208 32846 31260 32852
rect 31300 32904 31352 32910
rect 31300 32846 31352 32852
rect 31220 32434 31248 32846
rect 31208 32428 31260 32434
rect 31260 32388 31340 32416
rect 31208 32370 31260 32376
rect 31116 32224 31168 32230
rect 31116 32166 31168 32172
rect 31024 32020 31076 32026
rect 31024 31962 31076 31968
rect 31128 31414 31156 32166
rect 31208 31816 31260 31822
rect 31208 31758 31260 31764
rect 31116 31408 31168 31414
rect 31116 31350 31168 31356
rect 30748 31340 30800 31346
rect 30748 31282 30800 31288
rect 30760 31226 30788 31282
rect 30380 31204 30432 31210
rect 30760 31198 30880 31226
rect 30380 31146 30432 31152
rect 29828 31136 29880 31142
rect 29828 31078 29880 31084
rect 30104 31136 30156 31142
rect 30104 31078 30156 31084
rect 29840 30734 29868 31078
rect 28816 30728 28868 30734
rect 28816 30670 28868 30676
rect 29552 30728 29604 30734
rect 29552 30670 29604 30676
rect 29828 30728 29880 30734
rect 29828 30670 29880 30676
rect 28172 30592 28224 30598
rect 28172 30534 28224 30540
rect 28540 30592 28592 30598
rect 28540 30534 28592 30540
rect 28552 30258 28580 30534
rect 27804 30252 27856 30258
rect 27804 30194 27856 30200
rect 27896 30252 27948 30258
rect 27896 30194 27948 30200
rect 28080 30252 28132 30258
rect 28080 30194 28132 30200
rect 28540 30252 28592 30258
rect 28540 30194 28592 30200
rect 27712 29844 27764 29850
rect 27712 29786 27764 29792
rect 27816 29510 27844 30194
rect 27908 29850 27936 30194
rect 28264 30184 28316 30190
rect 28264 30126 28316 30132
rect 27988 30116 28040 30122
rect 27988 30058 28040 30064
rect 28000 29850 28028 30058
rect 28172 30048 28224 30054
rect 28172 29990 28224 29996
rect 28184 29850 28212 29990
rect 27896 29844 27948 29850
rect 27896 29786 27948 29792
rect 27988 29844 28040 29850
rect 27988 29786 28040 29792
rect 28172 29844 28224 29850
rect 28172 29786 28224 29792
rect 27804 29504 27856 29510
rect 27804 29446 27856 29452
rect 27632 28920 27844 28948
rect 27712 28620 27764 28626
rect 27712 28562 27764 28568
rect 27344 28552 27396 28558
rect 27344 28494 27396 28500
rect 27160 28416 27212 28422
rect 27160 28358 27212 28364
rect 27172 28082 27200 28358
rect 27160 28076 27212 28082
rect 27160 28018 27212 28024
rect 25780 27464 25832 27470
rect 25780 27406 25832 27412
rect 26884 27464 26936 27470
rect 26884 27406 26936 27412
rect 26976 27464 27028 27470
rect 26976 27406 27028 27412
rect 25792 27130 25820 27406
rect 26272 27228 26580 27237
rect 26272 27226 26278 27228
rect 26334 27226 26358 27228
rect 26414 27226 26438 27228
rect 26494 27226 26518 27228
rect 26574 27226 26580 27228
rect 26334 27174 26336 27226
rect 26516 27174 26518 27226
rect 26272 27172 26278 27174
rect 26334 27172 26358 27174
rect 26414 27172 26438 27174
rect 26494 27172 26518 27174
rect 26574 27172 26580 27174
rect 26272 27163 26580 27172
rect 25780 27124 25832 27130
rect 25780 27066 25832 27072
rect 26896 26518 26924 27406
rect 26988 26586 27016 27406
rect 27356 26926 27384 28494
rect 27528 28416 27580 28422
rect 27528 28358 27580 28364
rect 27620 28416 27672 28422
rect 27620 28358 27672 28364
rect 27540 28218 27568 28358
rect 27528 28212 27580 28218
rect 27528 28154 27580 28160
rect 27632 28014 27660 28358
rect 27724 28218 27752 28562
rect 27712 28212 27764 28218
rect 27712 28154 27764 28160
rect 27620 28008 27672 28014
rect 27620 27950 27672 27956
rect 27436 27940 27488 27946
rect 27436 27882 27488 27888
rect 27448 27470 27476 27882
rect 27436 27464 27488 27470
rect 27436 27406 27488 27412
rect 27344 26920 27396 26926
rect 27344 26862 27396 26868
rect 26976 26580 27028 26586
rect 26976 26522 27028 26528
rect 27436 26580 27488 26586
rect 27436 26522 27488 26528
rect 26884 26512 26936 26518
rect 26884 26454 26936 26460
rect 27252 26444 27304 26450
rect 27252 26386 27304 26392
rect 26148 26376 26200 26382
rect 25594 26344 25650 26353
rect 26148 26318 26200 26324
rect 26240 26376 26292 26382
rect 26240 26318 26292 26324
rect 25594 26279 25650 26288
rect 25412 25900 25464 25906
rect 25412 25842 25464 25848
rect 25424 25294 25452 25842
rect 25412 25288 25464 25294
rect 25412 25230 25464 25236
rect 25504 25220 25556 25226
rect 25504 25162 25556 25168
rect 25044 24948 25096 24954
rect 25044 24890 25096 24896
rect 24952 24812 25004 24818
rect 24952 24754 25004 24760
rect 24676 24200 24728 24206
rect 24728 24148 24900 24154
rect 24676 24142 24900 24148
rect 24688 24126 24900 24142
rect 24400 23724 24452 23730
rect 24400 23666 24452 23672
rect 24492 23724 24544 23730
rect 24492 23666 24544 23672
rect 24412 23322 24440 23666
rect 24400 23316 24452 23322
rect 24400 23258 24452 23264
rect 23756 23112 23808 23118
rect 23756 23054 23808 23060
rect 24124 23112 24176 23118
rect 24124 23054 24176 23060
rect 23124 22778 23428 22794
rect 23020 22772 23072 22778
rect 23020 22714 23072 22720
rect 23124 22772 23440 22778
rect 23124 22766 23388 22772
rect 21364 22636 21416 22642
rect 21364 22578 21416 22584
rect 22100 22636 22152 22642
rect 22100 22578 22152 22584
rect 22928 22636 22980 22642
rect 22928 22578 22980 22584
rect 21376 22234 21404 22578
rect 21456 22432 21508 22438
rect 21456 22374 21508 22380
rect 21824 22432 21876 22438
rect 22112 22420 22140 22578
rect 22112 22392 22600 22420
rect 21824 22374 21876 22380
rect 21364 22228 21416 22234
rect 21364 22170 21416 22176
rect 21468 22094 21496 22374
rect 21468 22066 21680 22094
rect 21548 21888 21600 21894
rect 21548 21830 21600 21836
rect 20996 21548 21048 21554
rect 20996 21490 21048 21496
rect 21180 21548 21232 21554
rect 21180 21490 21232 21496
rect 20904 19440 20956 19446
rect 20904 19382 20956 19388
rect 20812 18964 20864 18970
rect 20812 18906 20864 18912
rect 19800 18702 19852 18708
rect 19628 18426 19656 18702
rect 18156 18380 18276 18408
rect 18328 18420 18380 18426
rect 17684 18216 17736 18222
rect 17684 18158 17736 18164
rect 17500 18080 17552 18086
rect 17500 18022 17552 18028
rect 17512 17882 17540 18022
rect 18156 17882 18184 18380
rect 18328 18362 18380 18368
rect 19616 18420 19668 18426
rect 19616 18362 19668 18368
rect 19812 18358 19840 18702
rect 19904 18686 20024 18714
rect 20536 18760 20588 18766
rect 20536 18702 20588 18708
rect 20720 18760 20772 18766
rect 20720 18702 20772 18708
rect 19340 18352 19392 18358
rect 19340 18294 19392 18300
rect 19800 18352 19852 18358
rect 19800 18294 19852 18300
rect 18236 18284 18288 18290
rect 18236 18226 18288 18232
rect 18788 18284 18840 18290
rect 18788 18226 18840 18232
rect 17500 17876 17552 17882
rect 17500 17818 17552 17824
rect 18144 17876 18196 17882
rect 18144 17818 18196 17824
rect 16132 17746 16252 17762
rect 16120 17740 16252 17746
rect 16172 17734 16252 17740
rect 16120 17682 16172 17688
rect 16120 17604 16172 17610
rect 16120 17546 16172 17552
rect 16132 17338 16160 17546
rect 16120 17332 16172 17338
rect 16120 17274 16172 17280
rect 16028 17264 16080 17270
rect 16028 17206 16080 17212
rect 5170 16892 5478 16901
rect 5170 16890 5176 16892
rect 5232 16890 5256 16892
rect 5312 16890 5336 16892
rect 5392 16890 5416 16892
rect 5472 16890 5478 16892
rect 5232 16838 5234 16890
rect 5414 16838 5416 16890
rect 5170 16836 5176 16838
rect 5232 16836 5256 16838
rect 5312 16836 5336 16838
rect 5392 16836 5416 16838
rect 5472 16836 5478 16838
rect 5170 16827 5478 16836
rect 13611 16892 13919 16901
rect 13611 16890 13617 16892
rect 13673 16890 13697 16892
rect 13753 16890 13777 16892
rect 13833 16890 13857 16892
rect 13913 16890 13919 16892
rect 13673 16838 13675 16890
rect 13855 16838 13857 16890
rect 13611 16836 13617 16838
rect 13673 16836 13697 16838
rect 13753 16836 13777 16838
rect 13833 16836 13857 16838
rect 13913 16836 13919 16838
rect 13611 16827 13919 16836
rect 9390 16348 9698 16357
rect 9390 16346 9396 16348
rect 9452 16346 9476 16348
rect 9532 16346 9556 16348
rect 9612 16346 9636 16348
rect 9692 16346 9698 16348
rect 9452 16294 9454 16346
rect 9634 16294 9636 16346
rect 9390 16292 9396 16294
rect 9452 16292 9476 16294
rect 9532 16292 9556 16294
rect 9612 16292 9636 16294
rect 9692 16292 9698 16294
rect 9390 16283 9698 16292
rect 5170 15804 5478 15813
rect 5170 15802 5176 15804
rect 5232 15802 5256 15804
rect 5312 15802 5336 15804
rect 5392 15802 5416 15804
rect 5472 15802 5478 15804
rect 5232 15750 5234 15802
rect 5414 15750 5416 15802
rect 5170 15748 5176 15750
rect 5232 15748 5256 15750
rect 5312 15748 5336 15750
rect 5392 15748 5416 15750
rect 5472 15748 5478 15750
rect 5170 15739 5478 15748
rect 13611 15804 13919 15813
rect 13611 15802 13617 15804
rect 13673 15802 13697 15804
rect 13753 15802 13777 15804
rect 13833 15802 13857 15804
rect 13913 15802 13919 15804
rect 13673 15750 13675 15802
rect 13855 15750 13857 15802
rect 13611 15748 13617 15750
rect 13673 15748 13697 15750
rect 13753 15748 13777 15750
rect 13833 15748 13857 15750
rect 13913 15748 13919 15750
rect 13611 15739 13919 15748
rect 9390 15260 9698 15269
rect 9390 15258 9396 15260
rect 9452 15258 9476 15260
rect 9532 15258 9556 15260
rect 9612 15258 9636 15260
rect 9692 15258 9698 15260
rect 9452 15206 9454 15258
rect 9634 15206 9636 15258
rect 9390 15204 9396 15206
rect 9452 15204 9476 15206
rect 9532 15204 9556 15206
rect 9612 15204 9636 15206
rect 9692 15204 9698 15206
rect 9390 15195 9698 15204
rect 5170 14716 5478 14725
rect 5170 14714 5176 14716
rect 5232 14714 5256 14716
rect 5312 14714 5336 14716
rect 5392 14714 5416 14716
rect 5472 14714 5478 14716
rect 5232 14662 5234 14714
rect 5414 14662 5416 14714
rect 5170 14660 5176 14662
rect 5232 14660 5256 14662
rect 5312 14660 5336 14662
rect 5392 14660 5416 14662
rect 5472 14660 5478 14662
rect 5170 14651 5478 14660
rect 13611 14716 13919 14725
rect 13611 14714 13617 14716
rect 13673 14714 13697 14716
rect 13753 14714 13777 14716
rect 13833 14714 13857 14716
rect 13913 14714 13919 14716
rect 13673 14662 13675 14714
rect 13855 14662 13857 14714
rect 13611 14660 13617 14662
rect 13673 14660 13697 14662
rect 13753 14660 13777 14662
rect 13833 14660 13857 14662
rect 13913 14660 13919 14662
rect 13611 14651 13919 14660
rect 1676 14340 1728 14346
rect 1676 14282 1728 14288
rect 1400 10056 1452 10062
rect 1400 9998 1452 10004
rect 1412 9625 1440 9998
rect 1398 9616 1454 9625
rect 1398 9551 1454 9560
rect 1688 2514 1716 14282
rect 9390 14172 9698 14181
rect 9390 14170 9396 14172
rect 9452 14170 9476 14172
rect 9532 14170 9556 14172
rect 9612 14170 9636 14172
rect 9692 14170 9698 14172
rect 9452 14118 9454 14170
rect 9634 14118 9636 14170
rect 9390 14116 9396 14118
rect 9452 14116 9476 14118
rect 9532 14116 9556 14118
rect 9612 14116 9636 14118
rect 9692 14116 9698 14118
rect 9390 14107 9698 14116
rect 5170 13628 5478 13637
rect 5170 13626 5176 13628
rect 5232 13626 5256 13628
rect 5312 13626 5336 13628
rect 5392 13626 5416 13628
rect 5472 13626 5478 13628
rect 5232 13574 5234 13626
rect 5414 13574 5416 13626
rect 5170 13572 5176 13574
rect 5232 13572 5256 13574
rect 5312 13572 5336 13574
rect 5392 13572 5416 13574
rect 5472 13572 5478 13574
rect 5170 13563 5478 13572
rect 13611 13628 13919 13637
rect 13611 13626 13617 13628
rect 13673 13626 13697 13628
rect 13753 13626 13777 13628
rect 13833 13626 13857 13628
rect 13913 13626 13919 13628
rect 13673 13574 13675 13626
rect 13855 13574 13857 13626
rect 13611 13572 13617 13574
rect 13673 13572 13697 13574
rect 13753 13572 13777 13574
rect 13833 13572 13857 13574
rect 13913 13572 13919 13574
rect 13611 13563 13919 13572
rect 9390 13084 9698 13093
rect 9390 13082 9396 13084
rect 9452 13082 9476 13084
rect 9532 13082 9556 13084
rect 9612 13082 9636 13084
rect 9692 13082 9698 13084
rect 9452 13030 9454 13082
rect 9634 13030 9636 13082
rect 9390 13028 9396 13030
rect 9452 13028 9476 13030
rect 9532 13028 9556 13030
rect 9612 13028 9636 13030
rect 9692 13028 9698 13030
rect 9390 13019 9698 13028
rect 5170 12540 5478 12549
rect 5170 12538 5176 12540
rect 5232 12538 5256 12540
rect 5312 12538 5336 12540
rect 5392 12538 5416 12540
rect 5472 12538 5478 12540
rect 5232 12486 5234 12538
rect 5414 12486 5416 12538
rect 5170 12484 5176 12486
rect 5232 12484 5256 12486
rect 5312 12484 5336 12486
rect 5392 12484 5416 12486
rect 5472 12484 5478 12486
rect 5170 12475 5478 12484
rect 13611 12540 13919 12549
rect 13611 12538 13617 12540
rect 13673 12538 13697 12540
rect 13753 12538 13777 12540
rect 13833 12538 13857 12540
rect 13913 12538 13919 12540
rect 13673 12486 13675 12538
rect 13855 12486 13857 12538
rect 13611 12484 13617 12486
rect 13673 12484 13697 12486
rect 13753 12484 13777 12486
rect 13833 12484 13857 12486
rect 13913 12484 13919 12486
rect 13611 12475 13919 12484
rect 16040 12238 16068 17206
rect 16224 17202 16252 17734
rect 18248 17542 18276 18226
rect 18420 18080 18472 18086
rect 18420 18022 18472 18028
rect 18512 18080 18564 18086
rect 18512 18022 18564 18028
rect 18432 17542 18460 18022
rect 17132 17536 17184 17542
rect 17132 17478 17184 17484
rect 18236 17536 18288 17542
rect 18236 17478 18288 17484
rect 18420 17536 18472 17542
rect 18420 17478 18472 17484
rect 17144 17338 17172 17478
rect 17831 17436 18139 17445
rect 17831 17434 17837 17436
rect 17893 17434 17917 17436
rect 17973 17434 17997 17436
rect 18053 17434 18077 17436
rect 18133 17434 18139 17436
rect 17893 17382 17895 17434
rect 18075 17382 18077 17434
rect 17831 17380 17837 17382
rect 17893 17380 17917 17382
rect 17973 17380 17997 17382
rect 18053 17380 18077 17382
rect 18133 17380 18139 17382
rect 17831 17371 18139 17380
rect 18248 17338 18276 17478
rect 17132 17332 17184 17338
rect 17132 17274 17184 17280
rect 18236 17332 18288 17338
rect 18236 17274 18288 17280
rect 18432 17202 18460 17478
rect 18524 17270 18552 18022
rect 18800 17338 18828 18226
rect 19352 17882 19380 18294
rect 19340 17876 19392 17882
rect 19340 17818 19392 17824
rect 19708 17536 19760 17542
rect 19708 17478 19760 17484
rect 18788 17332 18840 17338
rect 18788 17274 18840 17280
rect 18512 17264 18564 17270
rect 18512 17206 18564 17212
rect 19720 17202 19748 17478
rect 16212 17196 16264 17202
rect 16212 17138 16264 17144
rect 18420 17196 18472 17202
rect 18420 17138 18472 17144
rect 19432 17196 19484 17202
rect 19432 17138 19484 17144
rect 19708 17196 19760 17202
rect 19708 17138 19760 17144
rect 16224 16658 16252 17138
rect 18236 16992 18288 16998
rect 18236 16934 18288 16940
rect 16212 16652 16264 16658
rect 16212 16594 16264 16600
rect 17684 16448 17736 16454
rect 17684 16390 17736 16396
rect 17696 16250 17724 16390
rect 17831 16348 18139 16357
rect 17831 16346 17837 16348
rect 17893 16346 17917 16348
rect 17973 16346 17997 16348
rect 18053 16346 18077 16348
rect 18133 16346 18139 16348
rect 17893 16294 17895 16346
rect 18075 16294 18077 16346
rect 17831 16292 17837 16294
rect 17893 16292 17917 16294
rect 17973 16292 17997 16294
rect 18053 16292 18077 16294
rect 18133 16292 18139 16294
rect 17831 16283 18139 16292
rect 17684 16244 17736 16250
rect 17684 16186 17736 16192
rect 18248 16114 18276 16934
rect 18236 16108 18288 16114
rect 18236 16050 18288 16056
rect 18432 15978 18460 17138
rect 18972 17128 19024 17134
rect 18972 17070 19024 17076
rect 18984 16794 19012 17070
rect 19340 16992 19392 16998
rect 19340 16934 19392 16940
rect 19352 16794 19380 16934
rect 18972 16788 19024 16794
rect 18972 16730 19024 16736
rect 19340 16788 19392 16794
rect 19340 16730 19392 16736
rect 18512 16584 18564 16590
rect 18512 16526 18564 16532
rect 18524 16046 18552 16526
rect 18984 16250 19012 16730
rect 19444 16454 19472 17138
rect 19708 16992 19760 16998
rect 19708 16934 19760 16940
rect 19720 16658 19748 16934
rect 19904 16794 19932 18686
rect 19984 18624 20036 18630
rect 19984 18566 20036 18572
rect 19996 18426 20024 18566
rect 19984 18420 20036 18426
rect 19984 18362 20036 18368
rect 20260 17672 20312 17678
rect 20260 17614 20312 17620
rect 20076 17536 20128 17542
rect 20076 17478 20128 17484
rect 20168 17536 20220 17542
rect 20168 17478 20220 17484
rect 19984 17332 20036 17338
rect 19984 17274 20036 17280
rect 19892 16788 19944 16794
rect 19892 16730 19944 16736
rect 19708 16652 19760 16658
rect 19708 16594 19760 16600
rect 19708 16516 19760 16522
rect 19708 16458 19760 16464
rect 19432 16448 19484 16454
rect 19432 16390 19484 16396
rect 19444 16250 19472 16390
rect 18972 16244 19024 16250
rect 18972 16186 19024 16192
rect 19432 16244 19484 16250
rect 19432 16186 19484 16192
rect 18512 16040 18564 16046
rect 18512 15982 18564 15988
rect 18420 15972 18472 15978
rect 18420 15914 18472 15920
rect 17831 15260 18139 15269
rect 17831 15258 17837 15260
rect 17893 15258 17917 15260
rect 17973 15258 17997 15260
rect 18053 15258 18077 15260
rect 18133 15258 18139 15260
rect 17893 15206 17895 15258
rect 18075 15206 18077 15258
rect 17831 15204 17837 15206
rect 17893 15204 17917 15206
rect 17973 15204 17997 15206
rect 18053 15204 18077 15206
rect 18133 15204 18139 15206
rect 17831 15195 18139 15204
rect 17831 14172 18139 14181
rect 17831 14170 17837 14172
rect 17893 14170 17917 14172
rect 17973 14170 17997 14172
rect 18053 14170 18077 14172
rect 18133 14170 18139 14172
rect 17893 14118 17895 14170
rect 18075 14118 18077 14170
rect 17831 14116 17837 14118
rect 17893 14116 17917 14118
rect 17973 14116 17997 14118
rect 18053 14116 18077 14118
rect 18133 14116 18139 14118
rect 17831 14107 18139 14116
rect 17831 13084 18139 13093
rect 17831 13082 17837 13084
rect 17893 13082 17917 13084
rect 17973 13082 17997 13084
rect 18053 13082 18077 13084
rect 18133 13082 18139 13084
rect 17893 13030 17895 13082
rect 18075 13030 18077 13082
rect 17831 13028 17837 13030
rect 17893 13028 17917 13030
rect 17973 13028 17997 13030
rect 18053 13028 18077 13030
rect 18133 13028 18139 13030
rect 17831 13019 18139 13028
rect 16028 12232 16080 12238
rect 16028 12174 16080 12180
rect 9390 11996 9698 12005
rect 9390 11994 9396 11996
rect 9452 11994 9476 11996
rect 9532 11994 9556 11996
rect 9612 11994 9636 11996
rect 9692 11994 9698 11996
rect 9452 11942 9454 11994
rect 9634 11942 9636 11994
rect 9390 11940 9396 11942
rect 9452 11940 9476 11942
rect 9532 11940 9556 11942
rect 9612 11940 9636 11942
rect 9692 11940 9698 11942
rect 9390 11931 9698 11940
rect 17831 11996 18139 12005
rect 17831 11994 17837 11996
rect 17893 11994 17917 11996
rect 17973 11994 17997 11996
rect 18053 11994 18077 11996
rect 18133 11994 18139 11996
rect 17893 11942 17895 11994
rect 18075 11942 18077 11994
rect 17831 11940 17837 11942
rect 17893 11940 17917 11942
rect 17973 11940 17997 11942
rect 18053 11940 18077 11942
rect 18133 11940 18139 11942
rect 17831 11931 18139 11940
rect 5170 11452 5478 11461
rect 5170 11450 5176 11452
rect 5232 11450 5256 11452
rect 5312 11450 5336 11452
rect 5392 11450 5416 11452
rect 5472 11450 5478 11452
rect 5232 11398 5234 11450
rect 5414 11398 5416 11450
rect 5170 11396 5176 11398
rect 5232 11396 5256 11398
rect 5312 11396 5336 11398
rect 5392 11396 5416 11398
rect 5472 11396 5478 11398
rect 5170 11387 5478 11396
rect 13611 11452 13919 11461
rect 13611 11450 13617 11452
rect 13673 11450 13697 11452
rect 13753 11450 13777 11452
rect 13833 11450 13857 11452
rect 13913 11450 13919 11452
rect 13673 11398 13675 11450
rect 13855 11398 13857 11450
rect 13611 11396 13617 11398
rect 13673 11396 13697 11398
rect 13753 11396 13777 11398
rect 13833 11396 13857 11398
rect 13913 11396 13919 11398
rect 13611 11387 13919 11396
rect 9390 10908 9698 10917
rect 9390 10906 9396 10908
rect 9452 10906 9476 10908
rect 9532 10906 9556 10908
rect 9612 10906 9636 10908
rect 9692 10906 9698 10908
rect 9452 10854 9454 10906
rect 9634 10854 9636 10906
rect 9390 10852 9396 10854
rect 9452 10852 9476 10854
rect 9532 10852 9556 10854
rect 9612 10852 9636 10854
rect 9692 10852 9698 10854
rect 9390 10843 9698 10852
rect 17831 10908 18139 10917
rect 17831 10906 17837 10908
rect 17893 10906 17917 10908
rect 17973 10906 17997 10908
rect 18053 10906 18077 10908
rect 18133 10906 18139 10908
rect 17893 10854 17895 10906
rect 18075 10854 18077 10906
rect 17831 10852 17837 10854
rect 17893 10852 17917 10854
rect 17973 10852 17997 10854
rect 18053 10852 18077 10854
rect 18133 10852 18139 10854
rect 17831 10843 18139 10852
rect 5170 10364 5478 10373
rect 5170 10362 5176 10364
rect 5232 10362 5256 10364
rect 5312 10362 5336 10364
rect 5392 10362 5416 10364
rect 5472 10362 5478 10364
rect 5232 10310 5234 10362
rect 5414 10310 5416 10362
rect 5170 10308 5176 10310
rect 5232 10308 5256 10310
rect 5312 10308 5336 10310
rect 5392 10308 5416 10310
rect 5472 10308 5478 10310
rect 5170 10299 5478 10308
rect 13611 10364 13919 10373
rect 13611 10362 13617 10364
rect 13673 10362 13697 10364
rect 13753 10362 13777 10364
rect 13833 10362 13857 10364
rect 13913 10362 13919 10364
rect 13673 10310 13675 10362
rect 13855 10310 13857 10362
rect 13611 10308 13617 10310
rect 13673 10308 13697 10310
rect 13753 10308 13777 10310
rect 13833 10308 13857 10310
rect 13913 10308 13919 10310
rect 13611 10299 13919 10308
rect 9390 9820 9698 9829
rect 9390 9818 9396 9820
rect 9452 9818 9476 9820
rect 9532 9818 9556 9820
rect 9612 9818 9636 9820
rect 9692 9818 9698 9820
rect 9452 9766 9454 9818
rect 9634 9766 9636 9818
rect 9390 9764 9396 9766
rect 9452 9764 9476 9766
rect 9532 9764 9556 9766
rect 9612 9764 9636 9766
rect 9692 9764 9698 9766
rect 9390 9755 9698 9764
rect 17831 9820 18139 9829
rect 17831 9818 17837 9820
rect 17893 9818 17917 9820
rect 17973 9818 17997 9820
rect 18053 9818 18077 9820
rect 18133 9818 18139 9820
rect 17893 9766 17895 9818
rect 18075 9766 18077 9818
rect 17831 9764 17837 9766
rect 17893 9764 17917 9766
rect 17973 9764 17997 9766
rect 18053 9764 18077 9766
rect 18133 9764 18139 9766
rect 17831 9755 18139 9764
rect 5170 9276 5478 9285
rect 5170 9274 5176 9276
rect 5232 9274 5256 9276
rect 5312 9274 5336 9276
rect 5392 9274 5416 9276
rect 5472 9274 5478 9276
rect 5232 9222 5234 9274
rect 5414 9222 5416 9274
rect 5170 9220 5176 9222
rect 5232 9220 5256 9222
rect 5312 9220 5336 9222
rect 5392 9220 5416 9222
rect 5472 9220 5478 9222
rect 5170 9211 5478 9220
rect 13611 9276 13919 9285
rect 13611 9274 13617 9276
rect 13673 9274 13697 9276
rect 13753 9274 13777 9276
rect 13833 9274 13857 9276
rect 13913 9274 13919 9276
rect 13673 9222 13675 9274
rect 13855 9222 13857 9274
rect 13611 9220 13617 9222
rect 13673 9220 13697 9222
rect 13753 9220 13777 9222
rect 13833 9220 13857 9222
rect 13913 9220 13919 9222
rect 13611 9211 13919 9220
rect 9390 8732 9698 8741
rect 9390 8730 9396 8732
rect 9452 8730 9476 8732
rect 9532 8730 9556 8732
rect 9612 8730 9636 8732
rect 9692 8730 9698 8732
rect 9452 8678 9454 8730
rect 9634 8678 9636 8730
rect 9390 8676 9396 8678
rect 9452 8676 9476 8678
rect 9532 8676 9556 8678
rect 9612 8676 9636 8678
rect 9692 8676 9698 8678
rect 9390 8667 9698 8676
rect 17831 8732 18139 8741
rect 17831 8730 17837 8732
rect 17893 8730 17917 8732
rect 17973 8730 17997 8732
rect 18053 8730 18077 8732
rect 18133 8730 18139 8732
rect 17893 8678 17895 8730
rect 18075 8678 18077 8730
rect 17831 8676 17837 8678
rect 17893 8676 17917 8678
rect 17973 8676 17997 8678
rect 18053 8676 18077 8678
rect 18133 8676 18139 8678
rect 17831 8667 18139 8676
rect 5170 8188 5478 8197
rect 5170 8186 5176 8188
rect 5232 8186 5256 8188
rect 5312 8186 5336 8188
rect 5392 8186 5416 8188
rect 5472 8186 5478 8188
rect 5232 8134 5234 8186
rect 5414 8134 5416 8186
rect 5170 8132 5176 8134
rect 5232 8132 5256 8134
rect 5312 8132 5336 8134
rect 5392 8132 5416 8134
rect 5472 8132 5478 8134
rect 5170 8123 5478 8132
rect 13611 8188 13919 8197
rect 13611 8186 13617 8188
rect 13673 8186 13697 8188
rect 13753 8186 13777 8188
rect 13833 8186 13857 8188
rect 13913 8186 13919 8188
rect 13673 8134 13675 8186
rect 13855 8134 13857 8186
rect 13611 8132 13617 8134
rect 13673 8132 13697 8134
rect 13753 8132 13777 8134
rect 13833 8132 13857 8134
rect 13913 8132 13919 8134
rect 13611 8123 13919 8132
rect 9390 7644 9698 7653
rect 9390 7642 9396 7644
rect 9452 7642 9476 7644
rect 9532 7642 9556 7644
rect 9612 7642 9636 7644
rect 9692 7642 9698 7644
rect 9452 7590 9454 7642
rect 9634 7590 9636 7642
rect 9390 7588 9396 7590
rect 9452 7588 9476 7590
rect 9532 7588 9556 7590
rect 9612 7588 9636 7590
rect 9692 7588 9698 7590
rect 9390 7579 9698 7588
rect 17831 7644 18139 7653
rect 17831 7642 17837 7644
rect 17893 7642 17917 7644
rect 17973 7642 17997 7644
rect 18053 7642 18077 7644
rect 18133 7642 18139 7644
rect 17893 7590 17895 7642
rect 18075 7590 18077 7642
rect 17831 7588 17837 7590
rect 17893 7588 17917 7590
rect 17973 7588 17997 7590
rect 18053 7588 18077 7590
rect 18133 7588 18139 7590
rect 17831 7579 18139 7588
rect 5170 7100 5478 7109
rect 5170 7098 5176 7100
rect 5232 7098 5256 7100
rect 5312 7098 5336 7100
rect 5392 7098 5416 7100
rect 5472 7098 5478 7100
rect 5232 7046 5234 7098
rect 5414 7046 5416 7098
rect 5170 7044 5176 7046
rect 5232 7044 5256 7046
rect 5312 7044 5336 7046
rect 5392 7044 5416 7046
rect 5472 7044 5478 7046
rect 5170 7035 5478 7044
rect 13611 7100 13919 7109
rect 13611 7098 13617 7100
rect 13673 7098 13697 7100
rect 13753 7098 13777 7100
rect 13833 7098 13857 7100
rect 13913 7098 13919 7100
rect 13673 7046 13675 7098
rect 13855 7046 13857 7098
rect 13611 7044 13617 7046
rect 13673 7044 13697 7046
rect 13753 7044 13777 7046
rect 13833 7044 13857 7046
rect 13913 7044 13919 7046
rect 13611 7035 13919 7044
rect 19720 6914 19748 16458
rect 19892 16448 19944 16454
rect 19892 16390 19944 16396
rect 19904 16182 19932 16390
rect 19892 16176 19944 16182
rect 19892 16118 19944 16124
rect 19996 15042 20024 17274
rect 20088 17202 20116 17478
rect 20076 17196 20128 17202
rect 20076 17138 20128 17144
rect 20180 16454 20208 17478
rect 20272 17338 20300 17614
rect 20352 17536 20404 17542
rect 20352 17478 20404 17484
rect 20364 17338 20392 17478
rect 20260 17332 20312 17338
rect 20260 17274 20312 17280
rect 20352 17332 20404 17338
rect 20352 17274 20404 17280
rect 20548 17202 20576 18702
rect 20720 18624 20772 18630
rect 20720 18566 20772 18572
rect 20732 18426 20760 18566
rect 20720 18420 20772 18426
rect 20720 18362 20772 18368
rect 20720 18284 20772 18290
rect 20720 18226 20772 18232
rect 20628 17672 20680 17678
rect 20732 17626 20760 18226
rect 20824 18154 20852 18906
rect 21008 18714 21036 21490
rect 21192 20806 21220 21490
rect 21560 21486 21588 21830
rect 21652 21690 21680 22066
rect 21836 22030 21864 22374
rect 22052 22332 22360 22341
rect 22052 22330 22058 22332
rect 22114 22330 22138 22332
rect 22194 22330 22218 22332
rect 22274 22330 22298 22332
rect 22354 22330 22360 22332
rect 22114 22278 22116 22330
rect 22296 22278 22298 22330
rect 22052 22276 22058 22278
rect 22114 22276 22138 22278
rect 22194 22276 22218 22278
rect 22274 22276 22298 22278
rect 22354 22276 22360 22278
rect 22052 22267 22360 22276
rect 21824 22024 21876 22030
rect 21824 21966 21876 21972
rect 22572 21894 22600 22392
rect 23124 22234 23152 22766
rect 23388 22714 23440 22720
rect 23388 22636 23440 22642
rect 23388 22578 23440 22584
rect 23112 22228 23164 22234
rect 23112 22170 23164 22176
rect 21916 21888 21968 21894
rect 21916 21830 21968 21836
rect 22560 21888 22612 21894
rect 22560 21830 22612 21836
rect 21640 21684 21692 21690
rect 21640 21626 21692 21632
rect 21928 21622 21956 21830
rect 22376 21684 22428 21690
rect 22376 21626 22428 21632
rect 21916 21616 21968 21622
rect 21916 21558 21968 21564
rect 21928 21486 21956 21558
rect 21548 21480 21600 21486
rect 21548 21422 21600 21428
rect 21916 21480 21968 21486
rect 21916 21422 21968 21428
rect 21928 21146 21956 21422
rect 22052 21244 22360 21253
rect 22052 21242 22058 21244
rect 22114 21242 22138 21244
rect 22194 21242 22218 21244
rect 22274 21242 22298 21244
rect 22354 21242 22360 21244
rect 22114 21190 22116 21242
rect 22296 21190 22298 21242
rect 22052 21188 22058 21190
rect 22114 21188 22138 21190
rect 22194 21188 22218 21190
rect 22274 21188 22298 21190
rect 22354 21188 22360 21190
rect 22052 21179 22360 21188
rect 21916 21140 21968 21146
rect 21916 21082 21968 21088
rect 21180 20800 21232 20806
rect 21180 20742 21232 20748
rect 21548 20800 21600 20806
rect 21548 20742 21600 20748
rect 21180 19848 21232 19854
rect 21180 19790 21232 19796
rect 21088 19372 21140 19378
rect 21088 19314 21140 19320
rect 21100 18834 21128 19314
rect 21088 18828 21140 18834
rect 21088 18770 21140 18776
rect 21008 18686 21128 18714
rect 20812 18148 20864 18154
rect 20812 18090 20864 18096
rect 20680 17620 20760 17626
rect 20628 17614 20760 17620
rect 20812 17672 20864 17678
rect 20812 17614 20864 17620
rect 20996 17672 21048 17678
rect 20996 17614 21048 17620
rect 20640 17598 20760 17614
rect 20824 17338 20852 17614
rect 20904 17604 20956 17610
rect 20904 17546 20956 17552
rect 20812 17332 20864 17338
rect 20812 17274 20864 17280
rect 20444 17196 20496 17202
rect 20444 17138 20496 17144
rect 20536 17196 20588 17202
rect 20536 17138 20588 17144
rect 20456 16590 20484 17138
rect 20916 16726 20944 17546
rect 21008 16794 21036 17614
rect 21100 16998 21128 18686
rect 21192 18630 21220 19790
rect 21364 19712 21416 19718
rect 21364 19654 21416 19660
rect 21376 19514 21404 19654
rect 21364 19508 21416 19514
rect 21364 19450 21416 19456
rect 21456 19372 21508 19378
rect 21456 19314 21508 19320
rect 21364 19304 21416 19310
rect 21364 19246 21416 19252
rect 21376 18816 21404 19246
rect 21468 18970 21496 19314
rect 21456 18964 21508 18970
rect 21456 18906 21508 18912
rect 21560 18834 21588 20742
rect 22052 20156 22360 20165
rect 22052 20154 22058 20156
rect 22114 20154 22138 20156
rect 22194 20154 22218 20156
rect 22274 20154 22298 20156
rect 22354 20154 22360 20156
rect 22114 20102 22116 20154
rect 22296 20102 22298 20154
rect 22052 20100 22058 20102
rect 22114 20100 22138 20102
rect 22194 20100 22218 20102
rect 22274 20100 22298 20102
rect 22354 20100 22360 20102
rect 22052 20091 22360 20100
rect 21916 19984 21968 19990
rect 21916 19926 21968 19932
rect 21732 19712 21784 19718
rect 21732 19654 21784 19660
rect 21744 18970 21772 19654
rect 21928 19514 21956 19926
rect 22192 19916 22244 19922
rect 22192 19858 22244 19864
rect 21916 19508 21968 19514
rect 21916 19450 21968 19456
rect 21824 19440 21876 19446
rect 21824 19382 21876 19388
rect 21732 18964 21784 18970
rect 21732 18906 21784 18912
rect 21456 18828 21508 18834
rect 21376 18788 21456 18816
rect 21456 18770 21508 18776
rect 21548 18828 21600 18834
rect 21548 18770 21600 18776
rect 21180 18624 21232 18630
rect 21180 18566 21232 18572
rect 21468 17746 21496 18770
rect 21560 18290 21588 18770
rect 21836 18766 21864 19382
rect 22204 19242 22232 19858
rect 22388 19854 22416 21626
rect 22572 21554 22600 21830
rect 22560 21548 22612 21554
rect 22560 21490 22612 21496
rect 23020 21548 23072 21554
rect 23020 21490 23072 21496
rect 22572 21010 22600 21490
rect 22836 21344 22888 21350
rect 22836 21286 22888 21292
rect 22560 21004 22612 21010
rect 22560 20946 22612 20952
rect 22468 20528 22520 20534
rect 22468 20470 22520 20476
rect 22480 20058 22508 20470
rect 22652 20460 22704 20466
rect 22652 20402 22704 20408
rect 22468 20052 22520 20058
rect 22468 19994 22520 20000
rect 22376 19848 22428 19854
rect 22376 19790 22428 19796
rect 22388 19378 22416 19790
rect 22376 19372 22428 19378
rect 22376 19314 22428 19320
rect 22192 19236 22244 19242
rect 22192 19178 22244 19184
rect 22468 19168 22520 19174
rect 22468 19110 22520 19116
rect 22560 19168 22612 19174
rect 22560 19110 22612 19116
rect 22052 19068 22360 19077
rect 22052 19066 22058 19068
rect 22114 19066 22138 19068
rect 22194 19066 22218 19068
rect 22274 19066 22298 19068
rect 22354 19066 22360 19068
rect 22114 19014 22116 19066
rect 22296 19014 22298 19066
rect 22052 19012 22058 19014
rect 22114 19012 22138 19014
rect 22194 19012 22218 19014
rect 22274 19012 22298 19014
rect 22354 19012 22360 19014
rect 22052 19003 22360 19012
rect 21824 18760 21876 18766
rect 21824 18702 21876 18708
rect 21640 18624 21692 18630
rect 21640 18566 21692 18572
rect 21916 18624 21968 18630
rect 21916 18566 21968 18572
rect 21652 18426 21680 18566
rect 21640 18420 21692 18426
rect 21640 18362 21692 18368
rect 21548 18284 21600 18290
rect 21600 18244 21680 18272
rect 21548 18226 21600 18232
rect 21456 17740 21508 17746
rect 21456 17682 21508 17688
rect 21456 17536 21508 17542
rect 21456 17478 21508 17484
rect 21088 16992 21140 16998
rect 21088 16934 21140 16940
rect 20996 16788 21048 16794
rect 20996 16730 21048 16736
rect 20904 16720 20956 16726
rect 20904 16662 20956 16668
rect 20444 16584 20496 16590
rect 20444 16526 20496 16532
rect 20628 16584 20680 16590
rect 20628 16526 20680 16532
rect 20168 16448 20220 16454
rect 20168 16390 20220 16396
rect 20180 15978 20208 16390
rect 20640 16046 20668 16526
rect 20916 16402 20944 16662
rect 21468 16590 21496 17478
rect 21652 17134 21680 18244
rect 21928 17678 21956 18566
rect 22480 18290 22508 19110
rect 22572 18834 22600 19110
rect 22560 18828 22612 18834
rect 22560 18770 22612 18776
rect 22376 18284 22428 18290
rect 22376 18226 22428 18232
rect 22468 18284 22520 18290
rect 22468 18226 22520 18232
rect 22052 17980 22360 17989
rect 22052 17978 22058 17980
rect 22114 17978 22138 17980
rect 22194 17978 22218 17980
rect 22274 17978 22298 17980
rect 22354 17978 22360 17980
rect 22114 17926 22116 17978
rect 22296 17926 22298 17978
rect 22052 17924 22058 17926
rect 22114 17924 22138 17926
rect 22194 17924 22218 17926
rect 22274 17924 22298 17926
rect 22354 17924 22360 17926
rect 22052 17915 22360 17924
rect 22100 17876 22152 17882
rect 22100 17818 22152 17824
rect 21732 17672 21784 17678
rect 21732 17614 21784 17620
rect 21916 17672 21968 17678
rect 21916 17614 21968 17620
rect 21640 17128 21692 17134
rect 21640 17070 21692 17076
rect 21744 16998 21772 17614
rect 21824 17536 21876 17542
rect 21824 17478 21876 17484
rect 21836 17202 21864 17478
rect 21824 17196 21876 17202
rect 21824 17138 21876 17144
rect 21928 17082 21956 17614
rect 21836 17054 21956 17082
rect 21732 16992 21784 16998
rect 21732 16934 21784 16940
rect 21744 16794 21772 16934
rect 21836 16794 21864 17054
rect 22112 16980 22140 17818
rect 22388 17678 22416 18226
rect 22480 17814 22508 18226
rect 22572 17882 22600 18770
rect 22664 18766 22692 20402
rect 22744 20256 22796 20262
rect 22744 20198 22796 20204
rect 22756 20058 22784 20198
rect 22744 20052 22796 20058
rect 22744 19994 22796 20000
rect 22848 19922 22876 21286
rect 23032 21146 23060 21490
rect 23124 21486 23152 22170
rect 23400 21894 23428 22578
rect 23664 22568 23716 22574
rect 23664 22510 23716 22516
rect 23388 21888 23440 21894
rect 23388 21830 23440 21836
rect 23112 21480 23164 21486
rect 23112 21422 23164 21428
rect 23020 21140 23072 21146
rect 23020 21082 23072 21088
rect 23032 20602 23060 21082
rect 23020 20596 23072 20602
rect 23020 20538 23072 20544
rect 22836 19916 22888 19922
rect 22836 19858 22888 19864
rect 22928 19712 22980 19718
rect 22928 19654 22980 19660
rect 22744 19372 22796 19378
rect 22744 19314 22796 19320
rect 22652 18760 22704 18766
rect 22652 18702 22704 18708
rect 22756 18612 22784 19314
rect 22940 18970 22968 19654
rect 23032 19446 23060 20538
rect 23204 20460 23256 20466
rect 23204 20402 23256 20408
rect 23112 20256 23164 20262
rect 23112 20198 23164 20204
rect 23124 19854 23152 20198
rect 23216 20058 23244 20402
rect 23204 20052 23256 20058
rect 23204 19994 23256 20000
rect 23112 19848 23164 19854
rect 23112 19790 23164 19796
rect 23020 19440 23072 19446
rect 23020 19382 23072 19388
rect 23400 19378 23428 21830
rect 23676 20466 23704 22510
rect 24308 22432 24360 22438
rect 24308 22374 24360 22380
rect 24320 22030 24348 22374
rect 24308 22024 24360 22030
rect 24308 21966 24360 21972
rect 24400 21888 24452 21894
rect 24400 21830 24452 21836
rect 24412 21622 24440 21830
rect 24400 21616 24452 21622
rect 24400 21558 24452 21564
rect 23940 21548 23992 21554
rect 23940 21490 23992 21496
rect 23952 21078 23980 21490
rect 24504 21434 24532 23666
rect 24872 23662 24900 24126
rect 24860 23656 24912 23662
rect 24860 23598 24912 23604
rect 24860 23044 24912 23050
rect 24860 22986 24912 22992
rect 24768 22568 24820 22574
rect 24768 22510 24820 22516
rect 24780 21690 24808 22510
rect 24768 21684 24820 21690
rect 24768 21626 24820 21632
rect 24412 21406 24532 21434
rect 24780 21418 24808 21626
rect 24768 21412 24820 21418
rect 23940 21072 23992 21078
rect 23940 21014 23992 21020
rect 23952 20942 23980 21014
rect 24032 21004 24084 21010
rect 24308 21004 24360 21010
rect 24084 20964 24308 20992
rect 24032 20946 24084 20952
rect 24308 20946 24360 20952
rect 23940 20936 23992 20942
rect 23940 20878 23992 20884
rect 23480 20460 23532 20466
rect 23480 20402 23532 20408
rect 23664 20460 23716 20466
rect 23664 20402 23716 20408
rect 23388 19372 23440 19378
rect 23388 19314 23440 19320
rect 22928 18964 22980 18970
rect 22928 18906 22980 18912
rect 23492 18766 23520 20402
rect 23676 19258 23704 20402
rect 23848 19372 23900 19378
rect 23848 19314 23900 19320
rect 23584 19230 23704 19258
rect 23584 18970 23612 19230
rect 23664 19168 23716 19174
rect 23664 19110 23716 19116
rect 23572 18964 23624 18970
rect 23572 18906 23624 18912
rect 23676 18766 23704 19110
rect 23860 18970 23888 19314
rect 23848 18964 23900 18970
rect 23848 18906 23900 18912
rect 23480 18760 23532 18766
rect 23480 18702 23532 18708
rect 23664 18760 23716 18766
rect 23664 18702 23716 18708
rect 22664 18584 22784 18612
rect 22560 17876 22612 17882
rect 22560 17818 22612 17824
rect 22468 17808 22520 17814
rect 22468 17750 22520 17756
rect 22376 17672 22428 17678
rect 22376 17614 22428 17620
rect 22284 17536 22336 17542
rect 22388 17524 22416 17614
rect 22336 17496 22416 17524
rect 22284 17478 22336 17484
rect 22296 17202 22324 17478
rect 22480 17354 22508 17750
rect 22388 17326 22508 17354
rect 22388 17202 22416 17326
rect 22284 17196 22336 17202
rect 22284 17138 22336 17144
rect 22376 17196 22428 17202
rect 22376 17138 22428 17144
rect 22468 17196 22520 17202
rect 22468 17138 22520 17144
rect 22376 17060 22428 17066
rect 22376 17002 22428 17008
rect 21928 16952 22140 16980
rect 21732 16788 21784 16794
rect 21732 16730 21784 16736
rect 21824 16788 21876 16794
rect 21824 16730 21876 16736
rect 21456 16584 21508 16590
rect 21456 16526 21508 16532
rect 21928 16522 21956 16952
rect 22052 16892 22360 16901
rect 22052 16890 22058 16892
rect 22114 16890 22138 16892
rect 22194 16890 22218 16892
rect 22274 16890 22298 16892
rect 22354 16890 22360 16892
rect 22114 16838 22116 16890
rect 22296 16838 22298 16890
rect 22052 16836 22058 16838
rect 22114 16836 22138 16838
rect 22194 16836 22218 16838
rect 22274 16836 22298 16838
rect 22354 16836 22360 16838
rect 22052 16827 22360 16836
rect 22388 16794 22416 17002
rect 22480 16794 22508 17138
rect 22376 16788 22428 16794
rect 22376 16730 22428 16736
rect 22468 16788 22520 16794
rect 22468 16730 22520 16736
rect 22572 16658 22600 17818
rect 22560 16652 22612 16658
rect 22560 16594 22612 16600
rect 21916 16516 21968 16522
rect 21916 16458 21968 16464
rect 21088 16448 21140 16454
rect 20916 16396 21088 16402
rect 20916 16390 21140 16396
rect 20916 16374 21128 16390
rect 20628 16040 20680 16046
rect 20628 15982 20680 15988
rect 20168 15972 20220 15978
rect 20168 15914 20220 15920
rect 20640 15162 20668 15982
rect 22052 15804 22360 15813
rect 22052 15802 22058 15804
rect 22114 15802 22138 15804
rect 22194 15802 22218 15804
rect 22274 15802 22298 15804
rect 22354 15802 22360 15804
rect 22114 15750 22116 15802
rect 22296 15750 22298 15802
rect 22052 15748 22058 15750
rect 22114 15748 22138 15750
rect 22194 15748 22218 15750
rect 22274 15748 22298 15750
rect 22354 15748 22360 15750
rect 22052 15739 22360 15748
rect 20628 15156 20680 15162
rect 20628 15098 20680 15104
rect 22664 15094 22692 18584
rect 22744 18080 22796 18086
rect 22744 18022 22796 18028
rect 22756 17882 22784 18022
rect 22744 17876 22796 17882
rect 22744 17818 22796 17824
rect 23112 17876 23164 17882
rect 23112 17818 23164 17824
rect 22928 17672 22980 17678
rect 22928 17614 22980 17620
rect 22744 17536 22796 17542
rect 22744 17478 22796 17484
rect 22756 17338 22784 17478
rect 22744 17332 22796 17338
rect 22744 17274 22796 17280
rect 22836 17332 22888 17338
rect 22836 17274 22888 17280
rect 22848 17202 22876 17274
rect 22836 17196 22888 17202
rect 22836 17138 22888 17144
rect 22940 17066 22968 17614
rect 23020 17196 23072 17202
rect 23020 17138 23072 17144
rect 22928 17060 22980 17066
rect 22928 17002 22980 17008
rect 22836 16992 22888 16998
rect 22836 16934 22888 16940
rect 22848 16590 22876 16934
rect 22940 16590 22968 17002
rect 23032 16794 23060 17138
rect 23020 16788 23072 16794
rect 23020 16730 23072 16736
rect 23124 16590 23152 17818
rect 23296 17808 23348 17814
rect 23296 17750 23348 17756
rect 23308 17678 23336 17750
rect 23204 17672 23256 17678
rect 23204 17614 23256 17620
rect 23296 17672 23348 17678
rect 23492 17660 23520 18702
rect 23676 18630 23704 18702
rect 23940 18692 23992 18698
rect 23940 18634 23992 18640
rect 23664 18624 23716 18630
rect 23664 18566 23716 18572
rect 23572 17672 23624 17678
rect 23492 17632 23572 17660
rect 23296 17614 23348 17620
rect 23572 17614 23624 17620
rect 23216 16794 23244 17614
rect 23584 17270 23612 17614
rect 23572 17264 23624 17270
rect 23572 17206 23624 17212
rect 23388 17196 23440 17202
rect 23388 17138 23440 17144
rect 23204 16788 23256 16794
rect 23256 16748 23336 16776
rect 23204 16730 23256 16736
rect 23308 16590 23336 16748
rect 22836 16584 22888 16590
rect 22836 16526 22888 16532
rect 22928 16584 22980 16590
rect 22928 16526 22980 16532
rect 23112 16584 23164 16590
rect 23112 16526 23164 16532
rect 23296 16584 23348 16590
rect 23296 16526 23348 16532
rect 23400 16522 23428 17138
rect 23676 16658 23704 18566
rect 23952 17882 23980 18634
rect 23940 17876 23992 17882
rect 23940 17818 23992 17824
rect 24308 17672 24360 17678
rect 24308 17614 24360 17620
rect 23664 16652 23716 16658
rect 23664 16594 23716 16600
rect 23388 16516 23440 16522
rect 23388 16458 23440 16464
rect 24320 15434 24348 17614
rect 24412 17338 24440 21406
rect 24768 21354 24820 21360
rect 24492 21344 24544 21350
rect 24492 21286 24544 21292
rect 24504 20890 24532 21286
rect 24504 20862 24624 20890
rect 24596 20806 24624 20862
rect 24584 20800 24636 20806
rect 24584 20742 24636 20748
rect 24872 19514 24900 22986
rect 24964 22778 24992 24754
rect 25136 24608 25188 24614
rect 25136 24550 25188 24556
rect 25148 23866 25176 24550
rect 25412 24064 25464 24070
rect 25412 24006 25464 24012
rect 25136 23860 25188 23866
rect 25136 23802 25188 23808
rect 25424 23798 25452 24006
rect 25412 23792 25464 23798
rect 25412 23734 25464 23740
rect 25424 23118 25452 23734
rect 25516 23322 25544 25162
rect 25608 23866 25636 26279
rect 25688 26240 25740 26246
rect 25688 26182 25740 26188
rect 25700 25906 25728 26182
rect 26160 25974 26188 26318
rect 26252 26246 26280 26318
rect 26240 26240 26292 26246
rect 26240 26182 26292 26188
rect 26700 26240 26752 26246
rect 26700 26182 26752 26188
rect 26272 26140 26580 26149
rect 26272 26138 26278 26140
rect 26334 26138 26358 26140
rect 26414 26138 26438 26140
rect 26494 26138 26518 26140
rect 26574 26138 26580 26140
rect 26334 26086 26336 26138
rect 26516 26086 26518 26138
rect 26272 26084 26278 26086
rect 26334 26084 26358 26086
rect 26414 26084 26438 26086
rect 26494 26084 26518 26086
rect 26574 26084 26580 26086
rect 26272 26075 26580 26084
rect 26712 26042 26740 26182
rect 26700 26036 26752 26042
rect 26700 25978 26752 25984
rect 26148 25968 26200 25974
rect 26148 25910 26200 25916
rect 25688 25900 25740 25906
rect 25688 25842 25740 25848
rect 26700 25900 26752 25906
rect 26700 25842 26752 25848
rect 25700 25430 25728 25842
rect 25872 25696 25924 25702
rect 25872 25638 25924 25644
rect 26056 25696 26108 25702
rect 26056 25638 26108 25644
rect 25884 25498 25912 25638
rect 25872 25492 25924 25498
rect 25872 25434 25924 25440
rect 25688 25424 25740 25430
rect 25688 25366 25740 25372
rect 25964 25220 26016 25226
rect 25964 25162 26016 25168
rect 25976 24954 26004 25162
rect 25964 24948 26016 24954
rect 25964 24890 26016 24896
rect 26068 24818 26096 25638
rect 26712 25498 26740 25842
rect 27264 25702 27292 26386
rect 27448 26382 27476 26522
rect 27344 26376 27396 26382
rect 27344 26318 27396 26324
rect 27436 26376 27488 26382
rect 27436 26318 27488 26324
rect 27356 26042 27384 26318
rect 27344 26036 27396 26042
rect 27344 25978 27396 25984
rect 27448 25838 27476 26318
rect 27632 26042 27660 27950
rect 27724 27878 27752 28154
rect 27712 27872 27764 27878
rect 27712 27814 27764 27820
rect 27724 27402 27752 27814
rect 27816 27588 27844 28920
rect 27908 28762 27936 29786
rect 28276 29306 28304 30126
rect 28540 30116 28592 30122
rect 28540 30058 28592 30064
rect 28632 30116 28684 30122
rect 28632 30058 28684 30064
rect 28448 30048 28500 30054
rect 28448 29990 28500 29996
rect 28264 29300 28316 29306
rect 28264 29242 28316 29248
rect 28460 29186 28488 29990
rect 28276 29170 28488 29186
rect 28264 29164 28488 29170
rect 28316 29158 28488 29164
rect 28264 29106 28316 29112
rect 27896 28756 27948 28762
rect 27896 28698 27948 28704
rect 27896 28416 27948 28422
rect 27896 28358 27948 28364
rect 28080 28416 28132 28422
rect 28080 28358 28132 28364
rect 27908 28014 27936 28358
rect 27896 28008 27948 28014
rect 27896 27950 27948 27956
rect 27988 27940 28040 27946
rect 27988 27882 28040 27888
rect 27896 27600 27948 27606
rect 27816 27560 27896 27588
rect 27712 27396 27764 27402
rect 27712 27338 27764 27344
rect 27816 26450 27844 27560
rect 27896 27542 27948 27548
rect 27896 27464 27948 27470
rect 28000 27452 28028 27882
rect 28092 27674 28120 28358
rect 28080 27668 28132 27674
rect 28080 27610 28132 27616
rect 28276 27470 28304 29106
rect 28552 29034 28580 30058
rect 28644 29850 28672 30058
rect 28632 29844 28684 29850
rect 28632 29786 28684 29792
rect 28632 29504 28684 29510
rect 28632 29446 28684 29452
rect 28644 29170 28672 29446
rect 28632 29164 28684 29170
rect 28632 29106 28684 29112
rect 28540 29028 28592 29034
rect 28540 28970 28592 28976
rect 28828 28218 28856 30670
rect 29564 29714 29592 30670
rect 30012 30592 30064 30598
rect 30012 30534 30064 30540
rect 30024 30258 30052 30534
rect 30116 30394 30144 31078
rect 30493 31036 30801 31045
rect 30493 31034 30499 31036
rect 30555 31034 30579 31036
rect 30635 31034 30659 31036
rect 30715 31034 30739 31036
rect 30795 31034 30801 31036
rect 30555 30982 30557 31034
rect 30737 30982 30739 31034
rect 30493 30980 30499 30982
rect 30555 30980 30579 30982
rect 30635 30980 30659 30982
rect 30715 30980 30739 30982
rect 30795 30980 30801 30982
rect 30493 30971 30801 30980
rect 30656 30592 30708 30598
rect 30656 30534 30708 30540
rect 30104 30388 30156 30394
rect 30104 30330 30156 30336
rect 30668 30258 30696 30534
rect 30012 30252 30064 30258
rect 30012 30194 30064 30200
rect 30656 30252 30708 30258
rect 30656 30194 30708 30200
rect 29828 30048 29880 30054
rect 29828 29990 29880 29996
rect 29552 29708 29604 29714
rect 29552 29650 29604 29656
rect 29840 29646 29868 29990
rect 30493 29948 30801 29957
rect 30493 29946 30499 29948
rect 30555 29946 30579 29948
rect 30635 29946 30659 29948
rect 30715 29946 30739 29948
rect 30795 29946 30801 29948
rect 30555 29894 30557 29946
rect 30737 29894 30739 29946
rect 30493 29892 30499 29894
rect 30555 29892 30579 29894
rect 30635 29892 30659 29894
rect 30715 29892 30739 29894
rect 30795 29892 30801 29894
rect 30493 29883 30801 29892
rect 29828 29640 29880 29646
rect 29828 29582 29880 29588
rect 28908 29572 28960 29578
rect 28908 29514 28960 29520
rect 28920 29306 28948 29514
rect 30852 29510 30880 31198
rect 30932 31136 30984 31142
rect 30932 31078 30984 31084
rect 31024 31136 31076 31142
rect 31024 31078 31076 31084
rect 30944 30394 30972 31078
rect 31036 30938 31064 31078
rect 31024 30932 31076 30938
rect 31024 30874 31076 30880
rect 30932 30388 30984 30394
rect 30932 30330 30984 30336
rect 31220 30122 31248 31758
rect 31312 31142 31340 32388
rect 31392 32224 31444 32230
rect 31392 32166 31444 32172
rect 32036 32224 32088 32230
rect 32036 32166 32088 32172
rect 31404 32026 31432 32166
rect 31392 32020 31444 32026
rect 31392 31962 31444 31968
rect 31404 31346 31432 31962
rect 31668 31884 31720 31890
rect 31668 31826 31720 31832
rect 31680 31414 31708 31826
rect 32048 31822 32076 32166
rect 32232 31890 32260 33458
rect 32220 31884 32272 31890
rect 32220 31826 32272 31832
rect 31852 31816 31904 31822
rect 31852 31758 31904 31764
rect 32036 31816 32088 31822
rect 32036 31758 32088 31764
rect 31668 31408 31720 31414
rect 31668 31350 31720 31356
rect 31392 31340 31444 31346
rect 31392 31282 31444 31288
rect 31300 31136 31352 31142
rect 31300 31078 31352 31084
rect 31680 30938 31708 31350
rect 31668 30932 31720 30938
rect 31668 30874 31720 30880
rect 31392 30660 31444 30666
rect 31392 30602 31444 30608
rect 31404 30394 31432 30602
rect 31392 30388 31444 30394
rect 31392 30330 31444 30336
rect 31864 30258 31892 31758
rect 32128 31680 32180 31686
rect 32128 31622 32180 31628
rect 31944 31340 31996 31346
rect 31944 31282 31996 31288
rect 31852 30252 31904 30258
rect 31852 30194 31904 30200
rect 31208 30116 31260 30122
rect 31208 30058 31260 30064
rect 30840 29504 30892 29510
rect 30840 29446 30892 29452
rect 28908 29300 28960 29306
rect 28908 29242 28960 29248
rect 30493 28860 30801 28869
rect 30493 28858 30499 28860
rect 30555 28858 30579 28860
rect 30635 28858 30659 28860
rect 30715 28858 30739 28860
rect 30795 28858 30801 28860
rect 30555 28806 30557 28858
rect 30737 28806 30739 28858
rect 30493 28804 30499 28806
rect 30555 28804 30579 28806
rect 30635 28804 30659 28806
rect 30715 28804 30739 28806
rect 30795 28804 30801 28806
rect 30493 28795 30801 28804
rect 29000 28620 29052 28626
rect 29000 28562 29052 28568
rect 29012 28218 29040 28562
rect 30380 28484 30432 28490
rect 30380 28426 30432 28432
rect 30392 28218 30420 28426
rect 28816 28212 28868 28218
rect 28816 28154 28868 28160
rect 29000 28212 29052 28218
rect 29000 28154 29052 28160
rect 30380 28212 30432 28218
rect 30380 28154 30432 28160
rect 29000 28076 29052 28082
rect 29000 28018 29052 28024
rect 29184 28076 29236 28082
rect 29184 28018 29236 28024
rect 29012 27606 29040 28018
rect 29000 27600 29052 27606
rect 29000 27542 29052 27548
rect 27948 27424 28028 27452
rect 28264 27464 28316 27470
rect 27896 27406 27948 27412
rect 28264 27406 28316 27412
rect 28724 27464 28776 27470
rect 28724 27406 28776 27412
rect 28908 27464 28960 27470
rect 28908 27406 28960 27412
rect 28736 26518 28764 27406
rect 28816 27396 28868 27402
rect 28816 27338 28868 27344
rect 28828 26994 28856 27338
rect 28920 27130 28948 27406
rect 28908 27124 28960 27130
rect 28908 27066 28960 27072
rect 29012 26994 29040 27542
rect 29092 27328 29144 27334
rect 29092 27270 29144 27276
rect 28816 26988 28868 26994
rect 28816 26930 28868 26936
rect 29000 26988 29052 26994
rect 29000 26930 29052 26936
rect 28828 26874 28856 26930
rect 29104 26926 29132 27270
rect 29196 27130 29224 28018
rect 29368 27940 29420 27946
rect 29368 27882 29420 27888
rect 29380 27130 29408 27882
rect 30493 27772 30801 27781
rect 30493 27770 30499 27772
rect 30555 27770 30579 27772
rect 30635 27770 30659 27772
rect 30715 27770 30739 27772
rect 30795 27770 30801 27772
rect 30555 27718 30557 27770
rect 30737 27718 30739 27770
rect 30493 27716 30499 27718
rect 30555 27716 30579 27718
rect 30635 27716 30659 27718
rect 30715 27716 30739 27718
rect 30795 27716 30801 27718
rect 30493 27707 30801 27716
rect 29184 27124 29236 27130
rect 29184 27066 29236 27072
rect 29368 27124 29420 27130
rect 29368 27066 29420 27072
rect 29092 26920 29144 26926
rect 28828 26846 28948 26874
rect 29092 26862 29144 26868
rect 28724 26512 28776 26518
rect 28724 26454 28776 26460
rect 27804 26444 27856 26450
rect 27804 26386 27856 26392
rect 28632 26376 28684 26382
rect 28632 26318 28684 26324
rect 27712 26240 27764 26246
rect 27712 26182 27764 26188
rect 27804 26240 27856 26246
rect 27804 26182 27856 26188
rect 27620 26036 27672 26042
rect 27620 25978 27672 25984
rect 27724 25838 27752 26182
rect 27436 25832 27488 25838
rect 27436 25774 27488 25780
rect 27712 25832 27764 25838
rect 27712 25774 27764 25780
rect 27252 25696 27304 25702
rect 27252 25638 27304 25644
rect 26700 25492 26752 25498
rect 26700 25434 26752 25440
rect 26272 25052 26580 25061
rect 26272 25050 26278 25052
rect 26334 25050 26358 25052
rect 26414 25050 26438 25052
rect 26494 25050 26518 25052
rect 26574 25050 26580 25052
rect 26334 24998 26336 25050
rect 26516 24998 26518 25050
rect 26272 24996 26278 24998
rect 26334 24996 26358 24998
rect 26414 24996 26438 24998
rect 26494 24996 26518 24998
rect 26574 24996 26580 24998
rect 26272 24987 26580 24996
rect 26712 24818 26740 25434
rect 27448 24818 27476 25774
rect 27816 25294 27844 26182
rect 28644 25906 28672 26318
rect 27896 25900 27948 25906
rect 27896 25842 27948 25848
rect 28632 25900 28684 25906
rect 28632 25842 28684 25848
rect 27908 25498 27936 25842
rect 28644 25498 28672 25842
rect 27896 25492 27948 25498
rect 27896 25434 27948 25440
rect 28632 25492 28684 25498
rect 28632 25434 28684 25440
rect 27804 25288 27856 25294
rect 27804 25230 27856 25236
rect 26056 24812 26108 24818
rect 26056 24754 26108 24760
rect 26700 24812 26752 24818
rect 26700 24754 26752 24760
rect 27436 24812 27488 24818
rect 27436 24754 27488 24760
rect 26148 24676 26200 24682
rect 26148 24618 26200 24624
rect 26056 24064 26108 24070
rect 26056 24006 26108 24012
rect 25596 23860 25648 23866
rect 25596 23802 25648 23808
rect 25872 23656 25924 23662
rect 25872 23598 25924 23604
rect 25504 23316 25556 23322
rect 25504 23258 25556 23264
rect 25412 23112 25464 23118
rect 25412 23054 25464 23060
rect 25424 22778 25452 23054
rect 24952 22772 25004 22778
rect 24952 22714 25004 22720
rect 25412 22772 25464 22778
rect 25412 22714 25464 22720
rect 25424 22642 25452 22714
rect 25412 22636 25464 22642
rect 25412 22578 25464 22584
rect 25044 22500 25096 22506
rect 25044 22442 25096 22448
rect 25056 21622 25084 22442
rect 25136 22432 25188 22438
rect 25136 22374 25188 22380
rect 25044 21616 25096 21622
rect 25044 21558 25096 21564
rect 25056 21434 25084 21558
rect 25148 21554 25176 22374
rect 25516 22094 25544 23258
rect 25884 23118 25912 23598
rect 26068 23322 26096 24006
rect 26160 23798 26188 24618
rect 28540 24608 28592 24614
rect 28540 24550 28592 24556
rect 28552 24410 28580 24550
rect 28540 24404 28592 24410
rect 28540 24346 28592 24352
rect 26272 23964 26580 23973
rect 26272 23962 26278 23964
rect 26334 23962 26358 23964
rect 26414 23962 26438 23964
rect 26494 23962 26518 23964
rect 26574 23962 26580 23964
rect 26334 23910 26336 23962
rect 26516 23910 26518 23962
rect 26272 23908 26278 23910
rect 26334 23908 26358 23910
rect 26414 23908 26438 23910
rect 26494 23908 26518 23910
rect 26574 23908 26580 23910
rect 26272 23899 26580 23908
rect 26148 23792 26200 23798
rect 26148 23734 26200 23740
rect 26516 23724 26568 23730
rect 26792 23724 26844 23730
rect 26568 23684 26648 23712
rect 26516 23666 26568 23672
rect 26332 23520 26384 23526
rect 26332 23462 26384 23468
rect 26056 23316 26108 23322
rect 26056 23258 26108 23264
rect 25872 23112 25924 23118
rect 25872 23054 25924 23060
rect 25884 22234 25912 23054
rect 26068 22642 26096 23258
rect 26344 23050 26372 23462
rect 26332 23044 26384 23050
rect 26332 22986 26384 22992
rect 26272 22876 26580 22885
rect 26272 22874 26278 22876
rect 26334 22874 26358 22876
rect 26414 22874 26438 22876
rect 26494 22874 26518 22876
rect 26574 22874 26580 22876
rect 26334 22822 26336 22874
rect 26516 22822 26518 22874
rect 26272 22820 26278 22822
rect 26334 22820 26358 22822
rect 26414 22820 26438 22822
rect 26494 22820 26518 22822
rect 26574 22820 26580 22822
rect 26272 22811 26580 22820
rect 26620 22778 26648 23684
rect 26792 23666 26844 23672
rect 26148 22772 26200 22778
rect 26148 22714 26200 22720
rect 26608 22772 26660 22778
rect 26608 22714 26660 22720
rect 26056 22636 26108 22642
rect 26056 22578 26108 22584
rect 25872 22228 25924 22234
rect 25872 22170 25924 22176
rect 25424 22066 25544 22094
rect 25320 21888 25372 21894
rect 25320 21830 25372 21836
rect 25332 21622 25360 21830
rect 25320 21616 25372 21622
rect 25320 21558 25372 21564
rect 25136 21548 25188 21554
rect 25136 21490 25188 21496
rect 25056 21418 25268 21434
rect 25056 21412 25280 21418
rect 25056 21406 25228 21412
rect 25228 21354 25280 21360
rect 25136 21344 25188 21350
rect 25136 21286 25188 21292
rect 25148 21010 25176 21286
rect 25136 21004 25188 21010
rect 25136 20946 25188 20952
rect 25332 20942 25360 21558
rect 25320 20936 25372 20942
rect 25320 20878 25372 20884
rect 24860 19508 24912 19514
rect 24860 19450 24912 19456
rect 24860 19372 24912 19378
rect 24860 19314 24912 19320
rect 25044 19372 25096 19378
rect 25044 19314 25096 19320
rect 24676 18080 24728 18086
rect 24676 18022 24728 18028
rect 24688 17678 24716 18022
rect 24676 17672 24728 17678
rect 24676 17614 24728 17620
rect 24400 17332 24452 17338
rect 24400 17274 24452 17280
rect 24872 17202 24900 19314
rect 24952 18284 25004 18290
rect 24952 18226 25004 18232
rect 24964 17338 24992 18226
rect 25056 17610 25084 19314
rect 25044 17604 25096 17610
rect 25044 17546 25096 17552
rect 24952 17332 25004 17338
rect 24952 17274 25004 17280
rect 24860 17196 24912 17202
rect 24860 17138 24912 17144
rect 25228 17196 25280 17202
rect 25228 17138 25280 17144
rect 24492 15904 24544 15910
rect 24492 15846 24544 15852
rect 24584 15904 24636 15910
rect 24584 15846 24636 15852
rect 24400 15496 24452 15502
rect 24400 15438 24452 15444
rect 24308 15428 24360 15434
rect 24308 15370 24360 15376
rect 24216 15360 24268 15366
rect 24216 15302 24268 15308
rect 24228 15094 24256 15302
rect 22652 15088 22704 15094
rect 19996 15026 20116 15042
rect 22652 15030 22704 15036
rect 24216 15088 24268 15094
rect 24216 15030 24268 15036
rect 19996 15020 20128 15026
rect 19996 15014 20076 15020
rect 20076 14962 20128 14968
rect 23296 15020 23348 15026
rect 23296 14962 23348 14968
rect 22052 14716 22360 14725
rect 22052 14714 22058 14716
rect 22114 14714 22138 14716
rect 22194 14714 22218 14716
rect 22274 14714 22298 14716
rect 22354 14714 22360 14716
rect 22114 14662 22116 14714
rect 22296 14662 22298 14714
rect 22052 14660 22058 14662
rect 22114 14660 22138 14662
rect 22194 14660 22218 14662
rect 22274 14660 22298 14662
rect 22354 14660 22360 14662
rect 22052 14651 22360 14660
rect 23308 14618 23336 14962
rect 24320 14958 24348 15370
rect 24412 15026 24440 15438
rect 24400 15020 24452 15026
rect 24400 14962 24452 14968
rect 24308 14952 24360 14958
rect 24308 14894 24360 14900
rect 23296 14612 23348 14618
rect 23296 14554 23348 14560
rect 24504 14414 24532 15846
rect 24596 15706 24624 15846
rect 24584 15700 24636 15706
rect 24584 15642 24636 15648
rect 24872 15434 24900 17138
rect 25240 16250 25268 17138
rect 25228 16244 25280 16250
rect 25228 16186 25280 16192
rect 24676 15428 24728 15434
rect 24676 15370 24728 15376
rect 24860 15428 24912 15434
rect 24860 15370 24912 15376
rect 24688 14618 24716 15370
rect 24676 14612 24728 14618
rect 24676 14554 24728 14560
rect 25424 14482 25452 22066
rect 25780 21956 25832 21962
rect 25780 21898 25832 21904
rect 25792 21690 25820 21898
rect 25596 21684 25648 21690
rect 25596 21626 25648 21632
rect 25780 21684 25832 21690
rect 25780 21626 25832 21632
rect 25608 21486 25636 21626
rect 25596 21480 25648 21486
rect 25596 21422 25648 21428
rect 25608 20942 25636 21422
rect 25596 20936 25648 20942
rect 25596 20878 25648 20884
rect 25884 19786 25912 22170
rect 26160 22030 26188 22714
rect 26700 22636 26752 22642
rect 26700 22578 26752 22584
rect 26240 22568 26292 22574
rect 26240 22510 26292 22516
rect 26148 22024 26200 22030
rect 26148 21966 26200 21972
rect 26252 21876 26280 22510
rect 26712 22234 26740 22578
rect 26700 22228 26752 22234
rect 26700 22170 26752 22176
rect 26804 22098 26832 23666
rect 27896 23520 27948 23526
rect 27896 23462 27948 23468
rect 27908 23118 27936 23462
rect 27896 23112 27948 23118
rect 27896 23054 27948 23060
rect 27252 22976 27304 22982
rect 27252 22918 27304 22924
rect 27344 22976 27396 22982
rect 27344 22918 27396 22924
rect 27264 22506 27292 22918
rect 27252 22500 27304 22506
rect 27252 22442 27304 22448
rect 27264 22098 27292 22442
rect 26332 22092 26384 22098
rect 26332 22034 26384 22040
rect 26792 22092 26844 22098
rect 26792 22034 26844 22040
rect 27252 22092 27304 22098
rect 27252 22034 27304 22040
rect 26344 21962 26372 22034
rect 26332 21956 26384 21962
rect 26332 21898 26384 21904
rect 26160 21848 26280 21876
rect 26884 21888 26936 21894
rect 26056 21480 26108 21486
rect 26056 21422 26108 21428
rect 26068 21078 26096 21422
rect 26056 21072 26108 21078
rect 26056 21014 26108 21020
rect 26160 20466 26188 21848
rect 26884 21830 26936 21836
rect 26272 21788 26580 21797
rect 26272 21786 26278 21788
rect 26334 21786 26358 21788
rect 26414 21786 26438 21788
rect 26494 21786 26518 21788
rect 26574 21786 26580 21788
rect 26334 21734 26336 21786
rect 26516 21734 26518 21786
rect 26272 21732 26278 21734
rect 26334 21732 26358 21734
rect 26414 21732 26438 21734
rect 26494 21732 26518 21734
rect 26574 21732 26580 21734
rect 26272 21723 26580 21732
rect 26608 20936 26660 20942
rect 26608 20878 26660 20884
rect 26792 20936 26844 20942
rect 26792 20878 26844 20884
rect 26272 20700 26580 20709
rect 26272 20698 26278 20700
rect 26334 20698 26358 20700
rect 26414 20698 26438 20700
rect 26494 20698 26518 20700
rect 26574 20698 26580 20700
rect 26334 20646 26336 20698
rect 26516 20646 26518 20698
rect 26272 20644 26278 20646
rect 26334 20644 26358 20646
rect 26414 20644 26438 20646
rect 26494 20644 26518 20646
rect 26574 20644 26580 20646
rect 26272 20635 26580 20644
rect 26620 20602 26648 20878
rect 26700 20800 26752 20806
rect 26700 20742 26752 20748
rect 26608 20596 26660 20602
rect 26608 20538 26660 20544
rect 26148 20460 26200 20466
rect 26148 20402 26200 20408
rect 25872 19780 25924 19786
rect 25872 19722 25924 19728
rect 25688 19508 25740 19514
rect 25688 19450 25740 19456
rect 25504 19372 25556 19378
rect 25504 19314 25556 19320
rect 25516 18426 25544 19314
rect 25596 19168 25648 19174
rect 25596 19110 25648 19116
rect 25504 18420 25556 18426
rect 25504 18362 25556 18368
rect 25608 17338 25636 19110
rect 25596 17332 25648 17338
rect 25596 17274 25648 17280
rect 25700 17066 25728 19450
rect 26160 19174 26188 20402
rect 26424 20256 26476 20262
rect 26424 20198 26476 20204
rect 26436 20058 26464 20198
rect 26424 20052 26476 20058
rect 26424 19994 26476 20000
rect 26272 19612 26580 19621
rect 26272 19610 26278 19612
rect 26334 19610 26358 19612
rect 26414 19610 26438 19612
rect 26494 19610 26518 19612
rect 26574 19610 26580 19612
rect 26334 19558 26336 19610
rect 26516 19558 26518 19610
rect 26272 19556 26278 19558
rect 26334 19556 26358 19558
rect 26414 19556 26438 19558
rect 26494 19556 26518 19558
rect 26574 19556 26580 19558
rect 26272 19547 26580 19556
rect 26148 19168 26200 19174
rect 26148 19110 26200 19116
rect 26608 18828 26660 18834
rect 26608 18770 26660 18776
rect 26272 18524 26580 18533
rect 26272 18522 26278 18524
rect 26334 18522 26358 18524
rect 26414 18522 26438 18524
rect 26494 18522 26518 18524
rect 26574 18522 26580 18524
rect 26334 18470 26336 18522
rect 26516 18470 26518 18522
rect 26272 18468 26278 18470
rect 26334 18468 26358 18470
rect 26414 18468 26438 18470
rect 26494 18468 26518 18470
rect 26574 18468 26580 18470
rect 26272 18459 26580 18468
rect 25872 18284 25924 18290
rect 25872 18226 25924 18232
rect 26056 18284 26108 18290
rect 26056 18226 26108 18232
rect 26516 18284 26568 18290
rect 26620 18272 26648 18770
rect 26712 18290 26740 20742
rect 26804 20058 26832 20878
rect 26896 20534 26924 21830
rect 27068 21548 27120 21554
rect 27068 21490 27120 21496
rect 26976 21344 27028 21350
rect 26976 21286 27028 21292
rect 26988 20942 27016 21286
rect 27080 21146 27108 21490
rect 27356 21146 27384 22918
rect 27908 22642 27936 23054
rect 27988 22976 28040 22982
rect 27988 22918 28040 22924
rect 28000 22778 28028 22918
rect 27988 22772 28040 22778
rect 27988 22714 28040 22720
rect 27896 22636 27948 22642
rect 27896 22578 27948 22584
rect 28736 22438 28764 26454
rect 28816 26376 28868 26382
rect 28816 26318 28868 26324
rect 28828 26042 28856 26318
rect 28920 26314 28948 26846
rect 29104 26586 29132 26862
rect 30493 26684 30801 26693
rect 30493 26682 30499 26684
rect 30555 26682 30579 26684
rect 30635 26682 30659 26684
rect 30715 26682 30739 26684
rect 30795 26682 30801 26684
rect 30555 26630 30557 26682
rect 30737 26630 30739 26682
rect 30493 26628 30499 26630
rect 30555 26628 30579 26630
rect 30635 26628 30659 26630
rect 30715 26628 30739 26630
rect 30795 26628 30801 26630
rect 30493 26619 30801 26628
rect 29092 26580 29144 26586
rect 29092 26522 29144 26528
rect 29552 26512 29604 26518
rect 29552 26454 29604 26460
rect 28908 26308 28960 26314
rect 28908 26250 28960 26256
rect 28816 26036 28868 26042
rect 28816 25978 28868 25984
rect 28920 25838 28948 26250
rect 29564 26042 29592 26454
rect 30852 26450 30880 29446
rect 31220 29102 31248 30058
rect 31576 30048 31628 30054
rect 31576 29990 31628 29996
rect 31588 29646 31616 29990
rect 31956 29850 31984 31282
rect 32140 30870 32168 31622
rect 32680 31340 32732 31346
rect 32680 31282 32732 31288
rect 32692 30938 32720 31282
rect 32680 30932 32732 30938
rect 32680 30874 32732 30880
rect 32128 30864 32180 30870
rect 32128 30806 32180 30812
rect 34164 30598 34192 39306
rect 34713 39196 35021 39205
rect 34713 39194 34719 39196
rect 34775 39194 34799 39196
rect 34855 39194 34879 39196
rect 34935 39194 34959 39196
rect 35015 39194 35021 39196
rect 34775 39142 34777 39194
rect 34957 39142 34959 39194
rect 34713 39140 34719 39142
rect 34775 39140 34799 39142
rect 34855 39140 34879 39142
rect 34935 39140 34959 39142
rect 35015 39140 35021 39142
rect 34713 39131 35021 39140
rect 34713 38108 35021 38117
rect 34713 38106 34719 38108
rect 34775 38106 34799 38108
rect 34855 38106 34879 38108
rect 34935 38106 34959 38108
rect 35015 38106 35021 38108
rect 34775 38054 34777 38106
rect 34957 38054 34959 38106
rect 34713 38052 34719 38054
rect 34775 38052 34799 38054
rect 34855 38052 34879 38054
rect 34935 38052 34959 38054
rect 35015 38052 35021 38054
rect 34713 38043 35021 38052
rect 34713 37020 35021 37029
rect 34713 37018 34719 37020
rect 34775 37018 34799 37020
rect 34855 37018 34879 37020
rect 34935 37018 34959 37020
rect 35015 37018 35021 37020
rect 34775 36966 34777 37018
rect 34957 36966 34959 37018
rect 34713 36964 34719 36966
rect 34775 36964 34799 36966
rect 34855 36964 34879 36966
rect 34935 36964 34959 36966
rect 35015 36964 35021 36966
rect 34713 36955 35021 36964
rect 34713 35932 35021 35941
rect 34713 35930 34719 35932
rect 34775 35930 34799 35932
rect 34855 35930 34879 35932
rect 34935 35930 34959 35932
rect 35015 35930 35021 35932
rect 34775 35878 34777 35930
rect 34957 35878 34959 35930
rect 34713 35876 34719 35878
rect 34775 35876 34799 35878
rect 34855 35876 34879 35878
rect 34935 35876 34959 35878
rect 35015 35876 35021 35878
rect 34713 35867 35021 35876
rect 34713 34844 35021 34853
rect 34713 34842 34719 34844
rect 34775 34842 34799 34844
rect 34855 34842 34879 34844
rect 34935 34842 34959 34844
rect 35015 34842 35021 34844
rect 34775 34790 34777 34842
rect 34957 34790 34959 34842
rect 34713 34788 34719 34790
rect 34775 34788 34799 34790
rect 34855 34788 34879 34790
rect 34935 34788 34959 34790
rect 35015 34788 35021 34790
rect 34713 34779 35021 34788
rect 34713 33756 35021 33765
rect 34713 33754 34719 33756
rect 34775 33754 34799 33756
rect 34855 33754 34879 33756
rect 34935 33754 34959 33756
rect 35015 33754 35021 33756
rect 34775 33702 34777 33754
rect 34957 33702 34959 33754
rect 34713 33700 34719 33702
rect 34775 33700 34799 33702
rect 34855 33700 34879 33702
rect 34935 33700 34959 33702
rect 35015 33700 35021 33702
rect 34713 33691 35021 33700
rect 34713 32668 35021 32677
rect 34713 32666 34719 32668
rect 34775 32666 34799 32668
rect 34855 32666 34879 32668
rect 34935 32666 34959 32668
rect 35015 32666 35021 32668
rect 34775 32614 34777 32666
rect 34957 32614 34959 32666
rect 34713 32612 34719 32614
rect 34775 32612 34799 32614
rect 34855 32612 34879 32614
rect 34935 32612 34959 32614
rect 35015 32612 35021 32614
rect 34713 32603 35021 32612
rect 34888 32428 34940 32434
rect 34888 32370 34940 32376
rect 34900 32065 34928 32370
rect 34886 32056 34942 32065
rect 34886 31991 34942 32000
rect 34713 31580 35021 31589
rect 34713 31578 34719 31580
rect 34775 31578 34799 31580
rect 34855 31578 34879 31580
rect 34935 31578 34959 31580
rect 35015 31578 35021 31580
rect 34775 31526 34777 31578
rect 34957 31526 34959 31578
rect 34713 31524 34719 31526
rect 34775 31524 34799 31526
rect 34855 31524 34879 31526
rect 34935 31524 34959 31526
rect 35015 31524 35021 31526
rect 34713 31515 35021 31524
rect 34152 30592 34204 30598
rect 34152 30534 34204 30540
rect 34713 30492 35021 30501
rect 34713 30490 34719 30492
rect 34775 30490 34799 30492
rect 34855 30490 34879 30492
rect 34935 30490 34959 30492
rect 35015 30490 35021 30492
rect 34775 30438 34777 30490
rect 34957 30438 34959 30490
rect 34713 30436 34719 30438
rect 34775 30436 34799 30438
rect 34855 30436 34879 30438
rect 34935 30436 34959 30438
rect 35015 30436 35021 30438
rect 34713 30427 35021 30436
rect 31944 29844 31996 29850
rect 31944 29786 31996 29792
rect 31576 29640 31628 29646
rect 31576 29582 31628 29588
rect 31576 29504 31628 29510
rect 31576 29446 31628 29452
rect 32404 29504 32456 29510
rect 32404 29446 32456 29452
rect 31208 29096 31260 29102
rect 31208 29038 31260 29044
rect 31024 28552 31076 28558
rect 31024 28494 31076 28500
rect 30932 28076 30984 28082
rect 30932 28018 30984 28024
rect 30944 26994 30972 28018
rect 31036 27470 31064 28494
rect 31220 28218 31248 29038
rect 31392 28416 31444 28422
rect 31392 28358 31444 28364
rect 31208 28212 31260 28218
rect 31208 28154 31260 28160
rect 31116 28076 31168 28082
rect 31116 28018 31168 28024
rect 31024 27464 31076 27470
rect 31024 27406 31076 27412
rect 30932 26988 30984 26994
rect 30932 26930 30984 26936
rect 30840 26444 30892 26450
rect 30840 26386 30892 26392
rect 31036 26382 31064 27406
rect 31128 27130 31156 28018
rect 31116 27124 31168 27130
rect 31116 27066 31168 27072
rect 31220 26994 31248 28154
rect 31404 28150 31432 28358
rect 31392 28144 31444 28150
rect 31392 28086 31444 28092
rect 31300 27872 31352 27878
rect 31300 27814 31352 27820
rect 31312 27470 31340 27814
rect 31588 27614 31616 29446
rect 32416 29102 32444 29446
rect 34713 29404 35021 29413
rect 34713 29402 34719 29404
rect 34775 29402 34799 29404
rect 34855 29402 34879 29404
rect 34935 29402 34959 29404
rect 35015 29402 35021 29404
rect 34775 29350 34777 29402
rect 34957 29350 34959 29402
rect 34713 29348 34719 29350
rect 34775 29348 34799 29350
rect 34855 29348 34879 29350
rect 34935 29348 34959 29350
rect 35015 29348 35021 29350
rect 34713 29339 35021 29348
rect 32404 29096 32456 29102
rect 32404 29038 32456 29044
rect 31852 28960 31904 28966
rect 31852 28902 31904 28908
rect 31864 28558 31892 28902
rect 31852 28552 31904 28558
rect 31852 28494 31904 28500
rect 32128 28416 32180 28422
rect 32128 28358 32180 28364
rect 31760 28212 31812 28218
rect 31760 28154 31812 28160
rect 31772 27962 31800 28154
rect 32140 28082 32168 28358
rect 32416 28218 32444 29038
rect 34713 28316 35021 28325
rect 34713 28314 34719 28316
rect 34775 28314 34799 28316
rect 34855 28314 34879 28316
rect 34935 28314 34959 28316
rect 35015 28314 35021 28316
rect 34775 28262 34777 28314
rect 34957 28262 34959 28314
rect 34713 28260 34719 28262
rect 34775 28260 34799 28262
rect 34855 28260 34879 28262
rect 34935 28260 34959 28262
rect 35015 28260 35021 28262
rect 34713 28251 35021 28260
rect 32404 28212 32456 28218
rect 32404 28154 32456 28160
rect 32128 28076 32180 28082
rect 32128 28018 32180 28024
rect 32404 28076 32456 28082
rect 32404 28018 32456 28024
rect 31680 27934 31800 27962
rect 31680 27878 31708 27934
rect 31668 27872 31720 27878
rect 31668 27814 31720 27820
rect 32416 27674 32444 28018
rect 32496 27872 32548 27878
rect 32496 27814 32548 27820
rect 32772 27872 32824 27878
rect 32772 27814 32824 27820
rect 31496 27586 31616 27614
rect 32404 27668 32456 27674
rect 32404 27610 32456 27616
rect 31300 27464 31352 27470
rect 31300 27406 31352 27412
rect 31496 27334 31524 27586
rect 31484 27328 31536 27334
rect 31484 27270 31536 27276
rect 31208 26988 31260 26994
rect 31208 26930 31260 26936
rect 29828 26376 29880 26382
rect 29828 26318 29880 26324
rect 31024 26376 31076 26382
rect 31024 26318 31076 26324
rect 29552 26036 29604 26042
rect 29552 25978 29604 25984
rect 28908 25832 28960 25838
rect 28908 25774 28960 25780
rect 28920 25362 28948 25774
rect 29368 25696 29420 25702
rect 29368 25638 29420 25644
rect 29380 25498 29408 25638
rect 29368 25492 29420 25498
rect 29368 25434 29420 25440
rect 28908 25356 28960 25362
rect 28908 25298 28960 25304
rect 29184 25288 29236 25294
rect 29090 25256 29146 25265
rect 29184 25230 29236 25236
rect 29368 25288 29420 25294
rect 29368 25230 29420 25236
rect 29090 25191 29092 25200
rect 29144 25191 29146 25200
rect 29092 25162 29144 25168
rect 29196 24954 29224 25230
rect 29184 24948 29236 24954
rect 29184 24890 29236 24896
rect 28908 24812 28960 24818
rect 28908 24754 28960 24760
rect 28920 24410 28948 24754
rect 29380 24732 29408 25230
rect 29564 25226 29592 25978
rect 29736 25832 29788 25838
rect 29736 25774 29788 25780
rect 29748 25498 29776 25774
rect 29736 25492 29788 25498
rect 29736 25434 29788 25440
rect 29840 25430 29868 26318
rect 30012 26240 30064 26246
rect 30012 26182 30064 26188
rect 30024 25906 30052 26182
rect 31220 26042 31248 26930
rect 31208 26036 31260 26042
rect 31208 25978 31260 25984
rect 30012 25900 30064 25906
rect 30012 25842 30064 25848
rect 30104 25900 30156 25906
rect 30104 25842 30156 25848
rect 30116 25786 30144 25842
rect 30024 25758 30144 25786
rect 30380 25764 30432 25770
rect 29920 25696 29972 25702
rect 30024 25684 30052 25758
rect 30380 25706 30432 25712
rect 29972 25656 30052 25684
rect 30104 25696 30156 25702
rect 29920 25638 29972 25644
rect 30104 25638 30156 25644
rect 30116 25498 30144 25638
rect 30104 25492 30156 25498
rect 30104 25434 30156 25440
rect 29828 25424 29880 25430
rect 29828 25366 29880 25372
rect 29552 25220 29604 25226
rect 29552 25162 29604 25168
rect 29564 24886 29592 25162
rect 29552 24880 29604 24886
rect 29552 24822 29604 24828
rect 29736 24744 29788 24750
rect 29380 24704 29736 24732
rect 29736 24686 29788 24692
rect 29552 24608 29604 24614
rect 29552 24550 29604 24556
rect 28908 24404 28960 24410
rect 28908 24346 28960 24352
rect 29564 24138 29592 24550
rect 29552 24132 29604 24138
rect 29552 24074 29604 24080
rect 29276 23724 29328 23730
rect 29276 23666 29328 23672
rect 29288 23186 29316 23666
rect 29276 23180 29328 23186
rect 29276 23122 29328 23128
rect 29000 23044 29052 23050
rect 29000 22986 29052 22992
rect 29184 23044 29236 23050
rect 29184 22986 29236 22992
rect 29012 22778 29040 22986
rect 29000 22772 29052 22778
rect 29000 22714 29052 22720
rect 27804 22432 27856 22438
rect 27804 22374 27856 22380
rect 28356 22432 28408 22438
rect 28356 22374 28408 22380
rect 28724 22432 28776 22438
rect 28724 22374 28776 22380
rect 27816 22094 27844 22374
rect 28368 22094 28396 22374
rect 27816 22066 27936 22094
rect 27528 21956 27580 21962
rect 27528 21898 27580 21904
rect 27068 21140 27120 21146
rect 27068 21082 27120 21088
rect 27344 21140 27396 21146
rect 27344 21082 27396 21088
rect 26976 20936 27028 20942
rect 26976 20878 27028 20884
rect 27436 20936 27488 20942
rect 27436 20878 27488 20884
rect 26884 20528 26936 20534
rect 26884 20470 26936 20476
rect 26792 20052 26844 20058
rect 26792 19994 26844 20000
rect 26804 19378 26832 19994
rect 26792 19372 26844 19378
rect 26792 19314 26844 19320
rect 26896 18766 26924 20470
rect 27448 20466 27476 20878
rect 27160 20460 27212 20466
rect 27160 20402 27212 20408
rect 27436 20460 27488 20466
rect 27436 20402 27488 20408
rect 26976 20256 27028 20262
rect 26976 20198 27028 20204
rect 26988 19854 27016 20198
rect 26976 19848 27028 19854
rect 26976 19790 27028 19796
rect 27172 19514 27200 20402
rect 27160 19508 27212 19514
rect 27160 19450 27212 19456
rect 26884 18760 26936 18766
rect 26884 18702 26936 18708
rect 27436 18760 27488 18766
rect 27540 18748 27568 21898
rect 27712 21072 27764 21078
rect 27712 21014 27764 21020
rect 27724 20602 27752 21014
rect 27804 20936 27856 20942
rect 27804 20878 27856 20884
rect 27816 20602 27844 20878
rect 27712 20596 27764 20602
rect 27712 20538 27764 20544
rect 27804 20596 27856 20602
rect 27804 20538 27856 20544
rect 27816 20058 27844 20538
rect 27908 20466 27936 22066
rect 28184 22066 28396 22094
rect 28184 22030 28212 22066
rect 28172 22024 28224 22030
rect 28172 21966 28224 21972
rect 28356 21888 28408 21894
rect 28356 21830 28408 21836
rect 28368 21622 28396 21830
rect 28356 21616 28408 21622
rect 28356 21558 28408 21564
rect 27988 21344 28040 21350
rect 27988 21286 28040 21292
rect 28000 20942 28028 21286
rect 27988 20936 28040 20942
rect 27988 20878 28040 20884
rect 27896 20460 27948 20466
rect 27896 20402 27948 20408
rect 28000 20330 28028 20878
rect 28736 20806 28764 22374
rect 29000 20868 29052 20874
rect 29000 20810 29052 20816
rect 28724 20800 28776 20806
rect 28724 20742 28776 20748
rect 28172 20460 28224 20466
rect 28172 20402 28224 20408
rect 27988 20324 28040 20330
rect 27988 20266 28040 20272
rect 27804 20052 27856 20058
rect 27804 19994 27856 20000
rect 28184 19446 28212 20402
rect 28172 19440 28224 19446
rect 28172 19382 28224 19388
rect 28736 19378 28764 20742
rect 29012 20602 29040 20810
rect 29000 20596 29052 20602
rect 29000 20538 29052 20544
rect 29196 20058 29224 22986
rect 29288 21554 29316 23122
rect 29564 22710 29592 24074
rect 29840 23866 29868 25366
rect 30104 25288 30156 25294
rect 30102 25256 30104 25265
rect 30156 25256 30158 25265
rect 30102 25191 30158 25200
rect 30392 24954 30420 25706
rect 30840 25696 30892 25702
rect 30840 25638 30892 25644
rect 30493 25596 30801 25605
rect 30493 25594 30499 25596
rect 30555 25594 30579 25596
rect 30635 25594 30659 25596
rect 30715 25594 30739 25596
rect 30795 25594 30801 25596
rect 30555 25542 30557 25594
rect 30737 25542 30739 25594
rect 30493 25540 30499 25542
rect 30555 25540 30579 25542
rect 30635 25540 30659 25542
rect 30715 25540 30739 25542
rect 30795 25540 30801 25542
rect 30493 25531 30801 25540
rect 30852 25294 30880 25638
rect 30840 25288 30892 25294
rect 30840 25230 30892 25236
rect 30380 24948 30432 24954
rect 30380 24890 30432 24896
rect 31220 24818 31248 25978
rect 31496 25906 31524 27270
rect 32416 27130 32444 27610
rect 32404 27124 32456 27130
rect 32404 27066 32456 27072
rect 32220 26784 32272 26790
rect 32220 26726 32272 26732
rect 32232 26382 32260 26726
rect 31760 26376 31812 26382
rect 31760 26318 31812 26324
rect 32220 26376 32272 26382
rect 32220 26318 32272 26324
rect 31484 25900 31536 25906
rect 31484 25842 31536 25848
rect 30840 24812 30892 24818
rect 30840 24754 30892 24760
rect 31116 24812 31168 24818
rect 31116 24754 31168 24760
rect 31208 24812 31260 24818
rect 31208 24754 31260 24760
rect 30493 24508 30801 24517
rect 30493 24506 30499 24508
rect 30555 24506 30579 24508
rect 30635 24506 30659 24508
rect 30715 24506 30739 24508
rect 30795 24506 30801 24508
rect 30555 24454 30557 24506
rect 30737 24454 30739 24506
rect 30493 24452 30499 24454
rect 30555 24452 30579 24454
rect 30635 24452 30659 24454
rect 30715 24452 30739 24454
rect 30795 24452 30801 24454
rect 30493 24443 30801 24452
rect 30852 24410 30880 24754
rect 30932 24744 30984 24750
rect 30932 24686 30984 24692
rect 30840 24404 30892 24410
rect 30840 24346 30892 24352
rect 29828 23860 29880 23866
rect 29828 23802 29880 23808
rect 29644 23724 29696 23730
rect 29644 23666 29696 23672
rect 30196 23724 30248 23730
rect 30196 23666 30248 23672
rect 29552 22704 29604 22710
rect 29552 22646 29604 22652
rect 29656 21962 29684 23666
rect 29920 23520 29972 23526
rect 29920 23462 29972 23468
rect 29932 23050 29960 23462
rect 30208 23322 30236 23666
rect 30493 23420 30801 23429
rect 30493 23418 30499 23420
rect 30555 23418 30579 23420
rect 30635 23418 30659 23420
rect 30715 23418 30739 23420
rect 30795 23418 30801 23420
rect 30555 23366 30557 23418
rect 30737 23366 30739 23418
rect 30493 23364 30499 23366
rect 30555 23364 30579 23366
rect 30635 23364 30659 23366
rect 30715 23364 30739 23366
rect 30795 23364 30801 23366
rect 30493 23355 30801 23364
rect 30944 23322 30972 24686
rect 31024 24608 31076 24614
rect 31024 24550 31076 24556
rect 31036 24410 31064 24550
rect 31024 24404 31076 24410
rect 31024 24346 31076 24352
rect 31024 24064 31076 24070
rect 31024 24006 31076 24012
rect 31036 23866 31064 24006
rect 31024 23860 31076 23866
rect 31024 23802 31076 23808
rect 30196 23316 30248 23322
rect 30196 23258 30248 23264
rect 30932 23316 30984 23322
rect 30932 23258 30984 23264
rect 30380 23112 30432 23118
rect 30380 23054 30432 23060
rect 29920 23044 29972 23050
rect 29920 22986 29972 22992
rect 30392 22574 30420 23054
rect 31024 22976 31076 22982
rect 31024 22918 31076 22924
rect 31036 22778 31064 22918
rect 31024 22772 31076 22778
rect 31024 22714 31076 22720
rect 30380 22568 30432 22574
rect 30380 22510 30432 22516
rect 30392 22234 30420 22510
rect 31128 22438 31156 24754
rect 31208 24676 31260 24682
rect 31208 24618 31260 24624
rect 31220 24410 31248 24618
rect 31496 24614 31524 25842
rect 31772 25702 31800 26318
rect 32312 25832 32364 25838
rect 32312 25774 32364 25780
rect 31576 25696 31628 25702
rect 31576 25638 31628 25644
rect 31760 25696 31812 25702
rect 31760 25638 31812 25644
rect 32128 25696 32180 25702
rect 32128 25638 32180 25644
rect 31588 25294 31616 25638
rect 31576 25288 31628 25294
rect 31576 25230 31628 25236
rect 31760 25220 31812 25226
rect 31760 25162 31812 25168
rect 31576 25152 31628 25158
rect 31576 25094 31628 25100
rect 31588 24818 31616 25094
rect 31772 24954 31800 25162
rect 31760 24948 31812 24954
rect 31760 24890 31812 24896
rect 31576 24812 31628 24818
rect 31576 24754 31628 24760
rect 32140 24682 32168 25638
rect 32324 25498 32352 25774
rect 32312 25492 32364 25498
rect 32312 25434 32364 25440
rect 32324 24818 32352 25434
rect 32508 24818 32536 27814
rect 32588 26036 32640 26042
rect 32588 25978 32640 25984
rect 32312 24812 32364 24818
rect 32312 24754 32364 24760
rect 32496 24812 32548 24818
rect 32496 24754 32548 24760
rect 32220 24744 32272 24750
rect 32220 24686 32272 24692
rect 32128 24676 32180 24682
rect 32128 24618 32180 24624
rect 31484 24608 31536 24614
rect 31484 24550 31536 24556
rect 31208 24404 31260 24410
rect 31208 24346 31260 24352
rect 32036 24132 32088 24138
rect 32036 24074 32088 24080
rect 31300 24064 31352 24070
rect 31300 24006 31352 24012
rect 31312 23866 31340 24006
rect 31300 23860 31352 23866
rect 31300 23802 31352 23808
rect 31944 23724 31996 23730
rect 31944 23666 31996 23672
rect 31208 23112 31260 23118
rect 31208 23054 31260 23060
rect 31116 22432 31168 22438
rect 31116 22374 31168 22380
rect 30493 22332 30801 22341
rect 30493 22330 30499 22332
rect 30555 22330 30579 22332
rect 30635 22330 30659 22332
rect 30715 22330 30739 22332
rect 30795 22330 30801 22332
rect 30555 22278 30557 22330
rect 30737 22278 30739 22330
rect 30493 22276 30499 22278
rect 30555 22276 30579 22278
rect 30635 22276 30659 22278
rect 30715 22276 30739 22278
rect 30795 22276 30801 22278
rect 30493 22267 30801 22276
rect 31220 22234 31248 23054
rect 31392 22432 31444 22438
rect 31392 22374 31444 22380
rect 31760 22432 31812 22438
rect 31760 22374 31812 22380
rect 30380 22228 30432 22234
rect 30380 22170 30432 22176
rect 31208 22228 31260 22234
rect 31208 22170 31260 22176
rect 30392 22094 30420 22170
rect 30024 22066 30420 22094
rect 29920 22024 29972 22030
rect 29920 21966 29972 21972
rect 29644 21956 29696 21962
rect 29644 21898 29696 21904
rect 29276 21548 29328 21554
rect 29276 21490 29328 21496
rect 29288 20942 29316 21490
rect 29932 21146 29960 21966
rect 30024 21554 30052 22066
rect 31404 22030 31432 22374
rect 31772 22098 31800 22374
rect 31760 22092 31812 22098
rect 31760 22034 31812 22040
rect 30472 22024 30524 22030
rect 30392 21984 30472 22012
rect 30196 21888 30248 21894
rect 30196 21830 30248 21836
rect 30208 21622 30236 21830
rect 30196 21616 30248 21622
rect 30196 21558 30248 21564
rect 30012 21548 30064 21554
rect 30012 21490 30064 21496
rect 29920 21140 29972 21146
rect 29920 21082 29972 21088
rect 30024 21010 30052 21490
rect 30012 21004 30064 21010
rect 30012 20946 30064 20952
rect 29276 20936 29328 20942
rect 29276 20878 29328 20884
rect 30392 20874 30420 21984
rect 30472 21966 30524 21972
rect 31116 22024 31168 22030
rect 31116 21966 31168 21972
rect 31208 22024 31260 22030
rect 31208 21966 31260 21972
rect 31392 22024 31444 22030
rect 31392 21966 31444 21972
rect 30840 21888 30892 21894
rect 30840 21830 30892 21836
rect 30493 21244 30801 21253
rect 30493 21242 30499 21244
rect 30555 21242 30579 21244
rect 30635 21242 30659 21244
rect 30715 21242 30739 21244
rect 30795 21242 30801 21244
rect 30555 21190 30557 21242
rect 30737 21190 30739 21242
rect 30493 21188 30499 21190
rect 30555 21188 30579 21190
rect 30635 21188 30659 21190
rect 30715 21188 30739 21190
rect 30795 21188 30801 21190
rect 30493 21179 30801 21188
rect 30852 20942 30880 21830
rect 31128 21690 31156 21966
rect 31116 21684 31168 21690
rect 31116 21626 31168 21632
rect 31220 21622 31248 21966
rect 31300 21888 31352 21894
rect 31300 21830 31352 21836
rect 31208 21616 31260 21622
rect 31208 21558 31260 21564
rect 31312 21418 31340 21830
rect 31772 21418 31800 22034
rect 31956 22030 31984 23666
rect 32048 22778 32076 24074
rect 32232 23662 32260 24686
rect 32600 24596 32628 25978
rect 32784 25838 32812 27814
rect 34713 27228 35021 27237
rect 34713 27226 34719 27228
rect 34775 27226 34799 27228
rect 34855 27226 34879 27228
rect 34935 27226 34959 27228
rect 35015 27226 35021 27228
rect 34775 27174 34777 27226
rect 34957 27174 34959 27226
rect 34713 27172 34719 27174
rect 34775 27172 34799 27174
rect 34855 27172 34879 27174
rect 34935 27172 34959 27174
rect 35015 27172 35021 27174
rect 34713 27163 35021 27172
rect 33048 26852 33100 26858
rect 33048 26794 33100 26800
rect 32956 26512 33008 26518
rect 32956 26454 33008 26460
rect 32968 25906 32996 26454
rect 32956 25900 33008 25906
rect 32956 25842 33008 25848
rect 32680 25832 32732 25838
rect 32680 25774 32732 25780
rect 32772 25832 32824 25838
rect 32772 25774 32824 25780
rect 32692 24818 32720 25774
rect 32680 24812 32732 24818
rect 32680 24754 32732 24760
rect 32864 24812 32916 24818
rect 32968 24800 32996 25842
rect 33060 24818 33088 26794
rect 34713 26140 35021 26149
rect 34713 26138 34719 26140
rect 34775 26138 34799 26140
rect 34855 26138 34879 26140
rect 34935 26138 34959 26140
rect 35015 26138 35021 26140
rect 34775 26086 34777 26138
rect 34957 26086 34959 26138
rect 34713 26084 34719 26086
rect 34775 26084 34799 26086
rect 34855 26084 34879 26086
rect 34935 26084 34959 26086
rect 35015 26084 35021 26086
rect 34713 26075 35021 26084
rect 34713 25052 35021 25061
rect 34713 25050 34719 25052
rect 34775 25050 34799 25052
rect 34855 25050 34879 25052
rect 34935 25050 34959 25052
rect 35015 25050 35021 25052
rect 34775 24998 34777 25050
rect 34957 24998 34959 25050
rect 34713 24996 34719 24998
rect 34775 24996 34799 24998
rect 34855 24996 34879 24998
rect 34935 24996 34959 24998
rect 35015 24996 35021 24998
rect 34713 24987 35021 24996
rect 32916 24772 32996 24800
rect 33048 24812 33100 24818
rect 32864 24754 32916 24760
rect 33048 24754 33100 24760
rect 32680 24608 32732 24614
rect 32600 24568 32680 24596
rect 32680 24550 32732 24556
rect 32588 24132 32640 24138
rect 32588 24074 32640 24080
rect 32600 23866 32628 24074
rect 32588 23860 32640 23866
rect 32588 23802 32640 23808
rect 32220 23656 32272 23662
rect 32220 23598 32272 23604
rect 33060 23474 33088 24754
rect 33324 24608 33376 24614
rect 33324 24550 33376 24556
rect 33336 24410 33364 24550
rect 33324 24404 33376 24410
rect 33324 24346 33376 24352
rect 34713 23964 35021 23973
rect 34713 23962 34719 23964
rect 34775 23962 34799 23964
rect 34855 23962 34879 23964
rect 34935 23962 34959 23964
rect 35015 23962 35021 23964
rect 34775 23910 34777 23962
rect 34957 23910 34959 23962
rect 34713 23908 34719 23910
rect 34775 23908 34799 23910
rect 34855 23908 34879 23910
rect 34935 23908 34959 23910
rect 35015 23908 35021 23910
rect 34713 23899 35021 23908
rect 32784 23446 33088 23474
rect 32036 22772 32088 22778
rect 32036 22714 32088 22720
rect 32784 22642 32812 23446
rect 34713 22876 35021 22885
rect 34713 22874 34719 22876
rect 34775 22874 34799 22876
rect 34855 22874 34879 22876
rect 34935 22874 34959 22876
rect 35015 22874 35021 22876
rect 34775 22822 34777 22874
rect 34957 22822 34959 22874
rect 34713 22820 34719 22822
rect 34775 22820 34799 22822
rect 34855 22820 34879 22822
rect 34935 22820 34959 22822
rect 35015 22820 35021 22822
rect 34713 22811 35021 22820
rect 32864 22704 32916 22710
rect 32864 22646 32916 22652
rect 32772 22636 32824 22642
rect 32772 22578 32824 22584
rect 32220 22500 32272 22506
rect 32220 22442 32272 22448
rect 32232 22030 32260 22442
rect 32784 22234 32812 22578
rect 32772 22228 32824 22234
rect 32772 22170 32824 22176
rect 31944 22024 31996 22030
rect 31944 21966 31996 21972
rect 32220 22024 32272 22030
rect 32220 21966 32272 21972
rect 32404 21548 32456 21554
rect 32404 21490 32456 21496
rect 32772 21548 32824 21554
rect 32772 21490 32824 21496
rect 31300 21412 31352 21418
rect 31300 21354 31352 21360
rect 31760 21412 31812 21418
rect 31760 21354 31812 21360
rect 32416 21146 32444 21490
rect 32496 21344 32548 21350
rect 32496 21286 32548 21292
rect 31944 21140 31996 21146
rect 31944 21082 31996 21088
rect 32404 21140 32456 21146
rect 32404 21082 32456 21088
rect 30840 20936 30892 20942
rect 30840 20878 30892 20884
rect 30380 20868 30432 20874
rect 30380 20810 30432 20816
rect 30932 20868 30984 20874
rect 30932 20810 30984 20816
rect 30392 20618 30420 20810
rect 30392 20590 30604 20618
rect 30576 20534 30604 20590
rect 30564 20528 30616 20534
rect 30564 20470 30616 20476
rect 30493 20156 30801 20165
rect 30493 20154 30499 20156
rect 30555 20154 30579 20156
rect 30635 20154 30659 20156
rect 30715 20154 30739 20156
rect 30795 20154 30801 20156
rect 30555 20102 30557 20154
rect 30737 20102 30739 20154
rect 30493 20100 30499 20102
rect 30555 20100 30579 20102
rect 30635 20100 30659 20102
rect 30715 20100 30739 20102
rect 30795 20100 30801 20102
rect 30493 20091 30801 20100
rect 29184 20052 29236 20058
rect 29184 19994 29236 20000
rect 29552 20052 29604 20058
rect 29552 19994 29604 20000
rect 29368 19780 29420 19786
rect 29368 19722 29420 19728
rect 29380 19514 29408 19722
rect 29368 19508 29420 19514
rect 29368 19450 29420 19456
rect 29276 19440 29328 19446
rect 29276 19382 29328 19388
rect 28264 19372 28316 19378
rect 28264 19314 28316 19320
rect 28724 19372 28776 19378
rect 28724 19314 28776 19320
rect 29000 19372 29052 19378
rect 29000 19314 29052 19320
rect 29092 19372 29144 19378
rect 29092 19314 29144 19320
rect 28276 18970 28304 19314
rect 28448 19168 28500 19174
rect 28448 19110 28500 19116
rect 28264 18964 28316 18970
rect 28264 18906 28316 18912
rect 27488 18720 27568 18748
rect 27436 18702 27488 18708
rect 27540 18290 27568 18720
rect 27620 18692 27672 18698
rect 27620 18634 27672 18640
rect 27632 18426 27660 18634
rect 27620 18420 27672 18426
rect 27620 18362 27672 18368
rect 28460 18358 28488 19110
rect 29012 18970 29040 19314
rect 29000 18964 29052 18970
rect 29000 18906 29052 18912
rect 29104 18834 29132 19314
rect 29092 18828 29144 18834
rect 29092 18770 29144 18776
rect 29184 18692 29236 18698
rect 29184 18634 29236 18640
rect 28540 18624 28592 18630
rect 28540 18566 28592 18572
rect 28448 18352 28500 18358
rect 28448 18294 28500 18300
rect 26568 18244 26648 18272
rect 26516 18226 26568 18232
rect 25780 18148 25832 18154
rect 25780 18090 25832 18096
rect 25792 17882 25820 18090
rect 25780 17876 25832 17882
rect 25780 17818 25832 17824
rect 25884 17338 25912 18226
rect 25964 17604 26016 17610
rect 25964 17546 26016 17552
rect 25976 17338 26004 17546
rect 25872 17332 25924 17338
rect 25872 17274 25924 17280
rect 25964 17332 26016 17338
rect 25964 17274 26016 17280
rect 25688 17060 25740 17066
rect 25688 17002 25740 17008
rect 26068 16794 26096 18226
rect 26240 18080 26292 18086
rect 26240 18022 26292 18028
rect 26252 17524 26280 18022
rect 26160 17496 26280 17524
rect 26160 17338 26188 17496
rect 26272 17436 26580 17445
rect 26272 17434 26278 17436
rect 26334 17434 26358 17436
rect 26414 17434 26438 17436
rect 26494 17434 26518 17436
rect 26574 17434 26580 17436
rect 26334 17382 26336 17434
rect 26516 17382 26518 17434
rect 26272 17380 26278 17382
rect 26334 17380 26358 17382
rect 26414 17380 26438 17382
rect 26494 17380 26518 17382
rect 26574 17380 26580 17382
rect 26272 17371 26580 17380
rect 26620 17338 26648 18244
rect 26700 18284 26752 18290
rect 26700 18226 26752 18232
rect 26976 18284 27028 18290
rect 26976 18226 27028 18232
rect 27528 18284 27580 18290
rect 27528 18226 27580 18232
rect 26988 17338 27016 18226
rect 27896 18080 27948 18086
rect 27896 18022 27948 18028
rect 27908 17678 27936 18022
rect 27896 17672 27948 17678
rect 27896 17614 27948 17620
rect 28552 17542 28580 18566
rect 27252 17536 27304 17542
rect 27252 17478 27304 17484
rect 27344 17536 27396 17542
rect 27344 17478 27396 17484
rect 28540 17536 28592 17542
rect 28540 17478 28592 17484
rect 27264 17338 27292 17478
rect 26148 17332 26200 17338
rect 26148 17274 26200 17280
rect 26608 17332 26660 17338
rect 26608 17274 26660 17280
rect 26976 17332 27028 17338
rect 26976 17274 27028 17280
rect 27252 17332 27304 17338
rect 27252 17274 27304 17280
rect 26148 17196 26200 17202
rect 26148 17138 26200 17144
rect 26240 17196 26292 17202
rect 26240 17138 26292 17144
rect 26976 17196 27028 17202
rect 26976 17138 27028 17144
rect 26160 17066 26188 17138
rect 26148 17060 26200 17066
rect 26148 17002 26200 17008
rect 26160 16794 26188 17002
rect 26056 16788 26108 16794
rect 26056 16730 26108 16736
rect 26148 16788 26200 16794
rect 26148 16730 26200 16736
rect 26252 16726 26280 17138
rect 26424 17128 26476 17134
rect 26424 17070 26476 17076
rect 26332 16992 26384 16998
rect 26332 16934 26384 16940
rect 26240 16720 26292 16726
rect 26240 16662 26292 16668
rect 26240 16584 26292 16590
rect 26160 16532 26240 16538
rect 26160 16526 26292 16532
rect 26160 16510 26280 16526
rect 26344 16522 26372 16934
rect 26436 16794 26464 17070
rect 26700 17060 26752 17066
rect 26700 17002 26752 17008
rect 26424 16788 26476 16794
rect 26424 16730 26476 16736
rect 26608 16584 26660 16590
rect 26608 16526 26660 16532
rect 26332 16516 26384 16522
rect 26160 16250 26188 16510
rect 26332 16458 26384 16464
rect 26272 16348 26580 16357
rect 26272 16346 26278 16348
rect 26334 16346 26358 16348
rect 26414 16346 26438 16348
rect 26494 16346 26518 16348
rect 26574 16346 26580 16348
rect 26334 16294 26336 16346
rect 26516 16294 26518 16346
rect 26272 16292 26278 16294
rect 26334 16292 26358 16294
rect 26414 16292 26438 16294
rect 26494 16292 26518 16294
rect 26574 16292 26580 16294
rect 26272 16283 26580 16292
rect 26620 16250 26648 16526
rect 26148 16244 26200 16250
rect 26148 16186 26200 16192
rect 26608 16244 26660 16250
rect 26608 16186 26660 16192
rect 25780 16108 25832 16114
rect 25780 16050 25832 16056
rect 25964 16108 26016 16114
rect 25964 16050 26016 16056
rect 25792 14822 25820 16050
rect 25872 15904 25924 15910
rect 25872 15846 25924 15852
rect 25780 14816 25832 14822
rect 25780 14758 25832 14764
rect 25412 14476 25464 14482
rect 25412 14418 25464 14424
rect 25884 14414 25912 15846
rect 25976 15094 26004 16050
rect 26056 16040 26108 16046
rect 26056 15982 26108 15988
rect 26068 15706 26096 15982
rect 26240 15972 26292 15978
rect 26240 15914 26292 15920
rect 26056 15700 26108 15706
rect 26056 15642 26108 15648
rect 25964 15088 26016 15094
rect 25964 15030 26016 15036
rect 25976 14618 26004 15030
rect 26068 15026 26096 15642
rect 26252 15434 26280 15914
rect 26712 15586 26740 17002
rect 26792 16448 26844 16454
rect 26792 16390 26844 16396
rect 26804 16250 26832 16390
rect 26988 16250 27016 17138
rect 27356 16998 27384 17478
rect 27344 16992 27396 16998
rect 27344 16934 27396 16940
rect 28264 16584 28316 16590
rect 28264 16526 28316 16532
rect 26792 16244 26844 16250
rect 26792 16186 26844 16192
rect 26976 16244 27028 16250
rect 26976 16186 27028 16192
rect 27620 16108 27672 16114
rect 27620 16050 27672 16056
rect 26620 15558 26740 15586
rect 26240 15428 26292 15434
rect 26240 15370 26292 15376
rect 26148 15360 26200 15366
rect 26148 15302 26200 15308
rect 26160 15042 26188 15302
rect 26272 15260 26580 15269
rect 26272 15258 26278 15260
rect 26334 15258 26358 15260
rect 26414 15258 26438 15260
rect 26494 15258 26518 15260
rect 26574 15258 26580 15260
rect 26334 15206 26336 15258
rect 26516 15206 26518 15258
rect 26272 15204 26278 15206
rect 26334 15204 26358 15206
rect 26414 15204 26438 15206
rect 26494 15204 26518 15206
rect 26574 15204 26580 15206
rect 26272 15195 26580 15204
rect 26620 15162 26648 15558
rect 27632 15502 27660 16050
rect 28276 15706 28304 16526
rect 28448 16448 28500 16454
rect 28448 16390 28500 16396
rect 28460 16250 28488 16390
rect 28448 16244 28500 16250
rect 28448 16186 28500 16192
rect 28552 16114 28580 17478
rect 29092 16584 29144 16590
rect 29092 16526 29144 16532
rect 29104 16250 29132 16526
rect 29196 16454 29224 18634
rect 29288 17338 29316 19382
rect 29564 18766 29592 19994
rect 30944 19922 30972 20810
rect 31956 20806 31984 21082
rect 31944 20800 31996 20806
rect 31944 20742 31996 20748
rect 32508 20602 32536 21286
rect 32784 21146 32812 21490
rect 32772 21140 32824 21146
rect 32772 21082 32824 21088
rect 32496 20596 32548 20602
rect 32496 20538 32548 20544
rect 32876 20534 32904 22646
rect 34888 22024 34940 22030
rect 34886 21992 34888 22001
rect 34940 21992 34942 22001
rect 34886 21927 34942 21936
rect 33508 21888 33560 21894
rect 33508 21830 33560 21836
rect 33520 21690 33548 21830
rect 34713 21788 35021 21797
rect 34713 21786 34719 21788
rect 34775 21786 34799 21788
rect 34855 21786 34879 21788
rect 34935 21786 34959 21788
rect 35015 21786 35021 21788
rect 34775 21734 34777 21786
rect 34957 21734 34959 21786
rect 34713 21732 34719 21734
rect 34775 21732 34799 21734
rect 34855 21732 34879 21734
rect 34935 21732 34959 21734
rect 35015 21732 35021 21734
rect 34713 21723 35021 21732
rect 33508 21684 33560 21690
rect 33508 21626 33560 21632
rect 33520 21350 33548 21626
rect 33600 21480 33652 21486
rect 33600 21422 33652 21428
rect 33508 21344 33560 21350
rect 33508 21286 33560 21292
rect 33324 20868 33376 20874
rect 33324 20810 33376 20816
rect 33336 20602 33364 20810
rect 33324 20596 33376 20602
rect 33324 20538 33376 20544
rect 32864 20528 32916 20534
rect 32864 20470 32916 20476
rect 31208 20460 31260 20466
rect 31208 20402 31260 20408
rect 31944 20460 31996 20466
rect 31944 20402 31996 20408
rect 32404 20460 32456 20466
rect 32404 20402 32456 20408
rect 33232 20460 33284 20466
rect 33232 20402 33284 20408
rect 33508 20460 33560 20466
rect 33508 20402 33560 20408
rect 31220 20058 31248 20402
rect 31392 20256 31444 20262
rect 31392 20198 31444 20204
rect 31208 20052 31260 20058
rect 31208 19994 31260 20000
rect 30932 19916 30984 19922
rect 30932 19858 30984 19864
rect 31220 19496 31248 19994
rect 31404 19786 31432 20198
rect 31392 19780 31444 19786
rect 31392 19722 31444 19728
rect 31956 19514 31984 20402
rect 32220 20392 32272 20398
rect 32220 20334 32272 20340
rect 32128 19916 32180 19922
rect 32128 19858 32180 19864
rect 31944 19508 31996 19514
rect 31220 19468 31340 19496
rect 31208 19372 31260 19378
rect 31208 19314 31260 19320
rect 30840 19168 30892 19174
rect 30840 19110 30892 19116
rect 30493 19068 30801 19077
rect 30493 19066 30499 19068
rect 30555 19066 30579 19068
rect 30635 19066 30659 19068
rect 30715 19066 30739 19068
rect 30795 19066 30801 19068
rect 30555 19014 30557 19066
rect 30737 19014 30739 19066
rect 30493 19012 30499 19014
rect 30555 19012 30579 19014
rect 30635 19012 30659 19014
rect 30715 19012 30739 19014
rect 30795 19012 30801 19014
rect 30493 19003 30801 19012
rect 29644 18964 29696 18970
rect 29644 18906 29696 18912
rect 29552 18760 29604 18766
rect 29552 18702 29604 18708
rect 29460 18624 29512 18630
rect 29460 18566 29512 18572
rect 29472 18426 29500 18566
rect 29460 18420 29512 18426
rect 29460 18362 29512 18368
rect 29472 17882 29500 18362
rect 29460 17876 29512 17882
rect 29460 17818 29512 17824
rect 29276 17332 29328 17338
rect 29276 17274 29328 17280
rect 29472 17066 29500 17818
rect 29564 17338 29592 18702
rect 29656 18426 29684 18906
rect 30104 18760 30156 18766
rect 30104 18702 30156 18708
rect 30116 18426 30144 18702
rect 30380 18624 30432 18630
rect 30380 18566 30432 18572
rect 29644 18420 29696 18426
rect 29644 18362 29696 18368
rect 29736 18420 29788 18426
rect 29736 18362 29788 18368
rect 30104 18420 30156 18426
rect 30392 18408 30420 18566
rect 30104 18362 30156 18368
rect 30300 18380 30420 18408
rect 29656 17338 29684 18362
rect 29748 17338 29776 18362
rect 30300 17814 30328 18380
rect 30380 18284 30432 18290
rect 30380 18226 30432 18232
rect 30392 17882 30420 18226
rect 30852 18086 30880 19110
rect 31220 18970 31248 19314
rect 31208 18964 31260 18970
rect 31208 18906 31260 18912
rect 31312 18766 31340 19468
rect 31944 19450 31996 19456
rect 31956 18766 31984 19450
rect 32140 18834 32168 19858
rect 32232 19854 32260 20334
rect 32312 20324 32364 20330
rect 32312 20266 32364 20272
rect 32220 19848 32272 19854
rect 32220 19790 32272 19796
rect 32324 19310 32352 20266
rect 32416 19990 32444 20402
rect 32588 20256 32640 20262
rect 32588 20198 32640 20204
rect 33048 20256 33100 20262
rect 33048 20198 33100 20204
rect 32404 19984 32456 19990
rect 32404 19926 32456 19932
rect 32600 19718 32628 20198
rect 32588 19712 32640 19718
rect 32588 19654 32640 19660
rect 32864 19712 32916 19718
rect 32864 19654 32916 19660
rect 32312 19304 32364 19310
rect 32312 19246 32364 19252
rect 32128 18828 32180 18834
rect 32128 18770 32180 18776
rect 30932 18760 30984 18766
rect 30932 18702 30984 18708
rect 31300 18760 31352 18766
rect 31300 18702 31352 18708
rect 31944 18760 31996 18766
rect 31944 18702 31996 18708
rect 30840 18080 30892 18086
rect 30840 18022 30892 18028
rect 30493 17980 30801 17989
rect 30493 17978 30499 17980
rect 30555 17978 30579 17980
rect 30635 17978 30659 17980
rect 30715 17978 30739 17980
rect 30795 17978 30801 17980
rect 30555 17926 30557 17978
rect 30737 17926 30739 17978
rect 30493 17924 30499 17926
rect 30555 17924 30579 17926
rect 30635 17924 30659 17926
rect 30715 17924 30739 17926
rect 30795 17924 30801 17926
rect 30493 17915 30801 17924
rect 30380 17876 30432 17882
rect 30380 17818 30432 17824
rect 30288 17808 30340 17814
rect 30288 17750 30340 17756
rect 30840 17604 30892 17610
rect 30840 17546 30892 17552
rect 30852 17338 30880 17546
rect 29552 17332 29604 17338
rect 29552 17274 29604 17280
rect 29644 17332 29696 17338
rect 29644 17274 29696 17280
rect 29736 17332 29788 17338
rect 29736 17274 29788 17280
rect 30840 17332 30892 17338
rect 30840 17274 30892 17280
rect 30380 17196 30432 17202
rect 30380 17138 30432 17144
rect 29920 17128 29972 17134
rect 29920 17070 29972 17076
rect 29460 17060 29512 17066
rect 29460 17002 29512 17008
rect 29932 16794 29960 17070
rect 30392 16794 30420 17138
rect 30493 16892 30801 16901
rect 30493 16890 30499 16892
rect 30555 16890 30579 16892
rect 30635 16890 30659 16892
rect 30715 16890 30739 16892
rect 30795 16890 30801 16892
rect 30555 16838 30557 16890
rect 30737 16838 30739 16890
rect 30493 16836 30499 16838
rect 30555 16836 30579 16838
rect 30635 16836 30659 16838
rect 30715 16836 30739 16838
rect 30795 16836 30801 16838
rect 30493 16827 30801 16836
rect 30944 16794 30972 18702
rect 31392 18080 31444 18086
rect 31392 18022 31444 18028
rect 31404 17678 31432 18022
rect 32600 17954 32628 19654
rect 32876 19514 32904 19654
rect 32864 19508 32916 19514
rect 32864 19450 32916 19456
rect 33060 19446 33088 20198
rect 33140 19848 33192 19854
rect 33140 19790 33192 19796
rect 33152 19514 33180 19790
rect 33140 19508 33192 19514
rect 33140 19450 33192 19456
rect 33048 19440 33100 19446
rect 33048 19382 33100 19388
rect 33244 18970 33272 20402
rect 33520 20058 33548 20402
rect 33508 20052 33560 20058
rect 33508 19994 33560 20000
rect 33612 19854 33640 21422
rect 34713 20700 35021 20709
rect 34713 20698 34719 20700
rect 34775 20698 34799 20700
rect 34855 20698 34879 20700
rect 34935 20698 34959 20700
rect 35015 20698 35021 20700
rect 34775 20646 34777 20698
rect 34957 20646 34959 20698
rect 34713 20644 34719 20646
rect 34775 20644 34799 20646
rect 34855 20644 34879 20646
rect 34935 20644 34959 20646
rect 35015 20644 35021 20646
rect 34713 20635 35021 20644
rect 33600 19848 33652 19854
rect 33600 19790 33652 19796
rect 34713 19612 35021 19621
rect 34713 19610 34719 19612
rect 34775 19610 34799 19612
rect 34855 19610 34879 19612
rect 34935 19610 34959 19612
rect 35015 19610 35021 19612
rect 34775 19558 34777 19610
rect 34957 19558 34959 19610
rect 34713 19556 34719 19558
rect 34775 19556 34799 19558
rect 34855 19556 34879 19558
rect 34935 19556 34959 19558
rect 35015 19556 35021 19558
rect 34713 19547 35021 19556
rect 33232 18964 33284 18970
rect 33232 18906 33284 18912
rect 34713 18524 35021 18533
rect 34713 18522 34719 18524
rect 34775 18522 34799 18524
rect 34855 18522 34879 18524
rect 34935 18522 34959 18524
rect 35015 18522 35021 18524
rect 34775 18470 34777 18522
rect 34957 18470 34959 18522
rect 34713 18468 34719 18470
rect 34775 18468 34799 18470
rect 34855 18468 34879 18470
rect 34935 18468 34959 18470
rect 35015 18468 35021 18470
rect 34713 18459 35021 18468
rect 32232 17926 32628 17954
rect 31392 17672 31444 17678
rect 31392 17614 31444 17620
rect 29368 16788 29420 16794
rect 29368 16730 29420 16736
rect 29920 16788 29972 16794
rect 29920 16730 29972 16736
rect 30380 16788 30432 16794
rect 30380 16730 30432 16736
rect 30932 16788 30984 16794
rect 30932 16730 30984 16736
rect 29184 16448 29236 16454
rect 29184 16390 29236 16396
rect 29092 16244 29144 16250
rect 29092 16186 29144 16192
rect 28540 16108 28592 16114
rect 28540 16050 28592 16056
rect 28264 15700 28316 15706
rect 28264 15642 28316 15648
rect 28908 15632 28960 15638
rect 28908 15574 28960 15580
rect 28920 15502 28948 15574
rect 29104 15570 29132 16186
rect 29092 15564 29144 15570
rect 29092 15506 29144 15512
rect 27620 15496 27672 15502
rect 27620 15438 27672 15444
rect 28172 15496 28224 15502
rect 28172 15438 28224 15444
rect 28908 15496 28960 15502
rect 28908 15438 28960 15444
rect 26700 15428 26752 15434
rect 26700 15370 26752 15376
rect 26712 15162 26740 15370
rect 26608 15156 26660 15162
rect 26608 15098 26660 15104
rect 26700 15156 26752 15162
rect 26700 15098 26752 15104
rect 26160 15026 26280 15042
rect 27632 15026 27660 15438
rect 27988 15360 28040 15366
rect 27988 15302 28040 15308
rect 28000 15094 28028 15302
rect 27988 15088 28040 15094
rect 27988 15030 28040 15036
rect 26056 15020 26108 15026
rect 26160 15020 26292 15026
rect 26160 15014 26240 15020
rect 26056 14962 26108 14968
rect 26240 14962 26292 14968
rect 26516 15020 26568 15026
rect 26516 14962 26568 14968
rect 27620 15020 27672 15026
rect 27620 14962 27672 14968
rect 26528 14618 26556 14962
rect 27896 14816 27948 14822
rect 27896 14758 27948 14764
rect 25964 14612 26016 14618
rect 25964 14554 26016 14560
rect 26516 14612 26568 14618
rect 26516 14554 26568 14560
rect 27908 14414 27936 14758
rect 28184 14618 28212 15438
rect 29380 15434 29408 16730
rect 31404 16590 31432 17614
rect 30380 16584 30432 16590
rect 30380 16526 30432 16532
rect 30656 16584 30708 16590
rect 30656 16526 30708 16532
rect 31392 16584 31444 16590
rect 31392 16526 31444 16532
rect 29920 16448 29972 16454
rect 29920 16390 29972 16396
rect 30012 16448 30064 16454
rect 30012 16390 30064 16396
rect 29932 16250 29960 16390
rect 29920 16244 29972 16250
rect 29920 16186 29972 16192
rect 29736 16108 29788 16114
rect 29736 16050 29788 16056
rect 29748 15706 29776 16050
rect 30024 15706 30052 16390
rect 30392 16182 30420 16526
rect 30380 16176 30432 16182
rect 30380 16118 30432 16124
rect 30392 15706 30420 16118
rect 30668 15910 30696 16526
rect 31404 15994 31432 16526
rect 31484 16516 31536 16522
rect 31484 16458 31536 16464
rect 31312 15966 31432 15994
rect 30656 15904 30708 15910
rect 30656 15846 30708 15852
rect 30493 15804 30801 15813
rect 30493 15802 30499 15804
rect 30555 15802 30579 15804
rect 30635 15802 30659 15804
rect 30715 15802 30739 15804
rect 30795 15802 30801 15804
rect 30555 15750 30557 15802
rect 30737 15750 30739 15802
rect 30493 15748 30499 15750
rect 30555 15748 30579 15750
rect 30635 15748 30659 15750
rect 30715 15748 30739 15750
rect 30795 15748 30801 15750
rect 30493 15739 30801 15748
rect 29736 15700 29788 15706
rect 29736 15642 29788 15648
rect 30012 15700 30064 15706
rect 30012 15642 30064 15648
rect 30380 15700 30432 15706
rect 30380 15642 30432 15648
rect 31312 15502 31340 15966
rect 31392 15904 31444 15910
rect 31392 15846 31444 15852
rect 31300 15496 31352 15502
rect 31300 15438 31352 15444
rect 29368 15428 29420 15434
rect 29368 15370 29420 15376
rect 30564 15428 30616 15434
rect 30564 15370 30616 15376
rect 29380 15162 29408 15370
rect 30576 15162 30604 15370
rect 31404 15162 31432 15846
rect 31496 15706 31524 16458
rect 32232 16454 32260 17926
rect 34713 17436 35021 17445
rect 34713 17434 34719 17436
rect 34775 17434 34799 17436
rect 34855 17434 34879 17436
rect 34935 17434 34959 17436
rect 35015 17434 35021 17436
rect 34775 17382 34777 17434
rect 34957 17382 34959 17434
rect 34713 17380 34719 17382
rect 34775 17380 34799 17382
rect 34855 17380 34879 17382
rect 34935 17380 34959 17382
rect 35015 17380 35021 17382
rect 34713 17371 35021 17380
rect 32220 16448 32272 16454
rect 32220 16390 32272 16396
rect 34713 16348 35021 16357
rect 34713 16346 34719 16348
rect 34775 16346 34799 16348
rect 34855 16346 34879 16348
rect 34935 16346 34959 16348
rect 35015 16346 35021 16348
rect 34775 16294 34777 16346
rect 34957 16294 34959 16346
rect 34713 16292 34719 16294
rect 34775 16292 34799 16294
rect 34855 16292 34879 16294
rect 34935 16292 34959 16294
rect 35015 16292 35021 16294
rect 34713 16283 35021 16292
rect 31484 15700 31536 15706
rect 31484 15642 31536 15648
rect 31668 15496 31720 15502
rect 31668 15438 31720 15444
rect 31680 15162 31708 15438
rect 34713 15260 35021 15269
rect 34713 15258 34719 15260
rect 34775 15258 34799 15260
rect 34855 15258 34879 15260
rect 34935 15258 34959 15260
rect 35015 15258 35021 15260
rect 34775 15206 34777 15258
rect 34957 15206 34959 15258
rect 34713 15204 34719 15206
rect 34775 15204 34799 15206
rect 34855 15204 34879 15206
rect 34935 15204 34959 15206
rect 35015 15204 35021 15206
rect 34713 15195 35021 15204
rect 29368 15156 29420 15162
rect 29368 15098 29420 15104
rect 30564 15156 30616 15162
rect 30564 15098 30616 15104
rect 31392 15156 31444 15162
rect 31392 15098 31444 15104
rect 31668 15156 31720 15162
rect 31668 15098 31720 15104
rect 31484 15020 31536 15026
rect 31484 14962 31536 14968
rect 30493 14716 30801 14725
rect 30493 14714 30499 14716
rect 30555 14714 30579 14716
rect 30635 14714 30659 14716
rect 30715 14714 30739 14716
rect 30795 14714 30801 14716
rect 30555 14662 30557 14714
rect 30737 14662 30739 14714
rect 30493 14660 30499 14662
rect 30555 14660 30579 14662
rect 30635 14660 30659 14662
rect 30715 14660 30739 14662
rect 30795 14660 30801 14662
rect 30493 14651 30801 14660
rect 28172 14612 28224 14618
rect 28172 14554 28224 14560
rect 24492 14408 24544 14414
rect 24492 14350 24544 14356
rect 25872 14408 25924 14414
rect 25872 14350 25924 14356
rect 27896 14408 27948 14414
rect 27896 14350 27948 14356
rect 28448 14408 28500 14414
rect 28448 14350 28500 14356
rect 26272 14172 26580 14181
rect 26272 14170 26278 14172
rect 26334 14170 26358 14172
rect 26414 14170 26438 14172
rect 26494 14170 26518 14172
rect 26574 14170 26580 14172
rect 26334 14118 26336 14170
rect 26516 14118 26518 14170
rect 26272 14116 26278 14118
rect 26334 14116 26358 14118
rect 26414 14116 26438 14118
rect 26494 14116 26518 14118
rect 26574 14116 26580 14118
rect 26272 14107 26580 14116
rect 22052 13628 22360 13637
rect 22052 13626 22058 13628
rect 22114 13626 22138 13628
rect 22194 13626 22218 13628
rect 22274 13626 22298 13628
rect 22354 13626 22360 13628
rect 22114 13574 22116 13626
rect 22296 13574 22298 13626
rect 22052 13572 22058 13574
rect 22114 13572 22138 13574
rect 22194 13572 22218 13574
rect 22274 13572 22298 13574
rect 22354 13572 22360 13574
rect 22052 13563 22360 13572
rect 26272 13084 26580 13093
rect 26272 13082 26278 13084
rect 26334 13082 26358 13084
rect 26414 13082 26438 13084
rect 26494 13082 26518 13084
rect 26574 13082 26580 13084
rect 26334 13030 26336 13082
rect 26516 13030 26518 13082
rect 26272 13028 26278 13030
rect 26334 13028 26358 13030
rect 26414 13028 26438 13030
rect 26494 13028 26518 13030
rect 26574 13028 26580 13030
rect 26272 13019 26580 13028
rect 22052 12540 22360 12549
rect 22052 12538 22058 12540
rect 22114 12538 22138 12540
rect 22194 12538 22218 12540
rect 22274 12538 22298 12540
rect 22354 12538 22360 12540
rect 22114 12486 22116 12538
rect 22296 12486 22298 12538
rect 22052 12484 22058 12486
rect 22114 12484 22138 12486
rect 22194 12484 22218 12486
rect 22274 12484 22298 12486
rect 22354 12484 22360 12486
rect 22052 12475 22360 12484
rect 26272 11996 26580 12005
rect 26272 11994 26278 11996
rect 26334 11994 26358 11996
rect 26414 11994 26438 11996
rect 26494 11994 26518 11996
rect 26574 11994 26580 11996
rect 26334 11942 26336 11994
rect 26516 11942 26518 11994
rect 26272 11940 26278 11942
rect 26334 11940 26358 11942
rect 26414 11940 26438 11942
rect 26494 11940 26518 11942
rect 26574 11940 26580 11942
rect 26272 11931 26580 11940
rect 22052 11452 22360 11461
rect 22052 11450 22058 11452
rect 22114 11450 22138 11452
rect 22194 11450 22218 11452
rect 22274 11450 22298 11452
rect 22354 11450 22360 11452
rect 22114 11398 22116 11450
rect 22296 11398 22298 11450
rect 22052 11396 22058 11398
rect 22114 11396 22138 11398
rect 22194 11396 22218 11398
rect 22274 11396 22298 11398
rect 22354 11396 22360 11398
rect 22052 11387 22360 11396
rect 26272 10908 26580 10917
rect 26272 10906 26278 10908
rect 26334 10906 26358 10908
rect 26414 10906 26438 10908
rect 26494 10906 26518 10908
rect 26574 10906 26580 10908
rect 26334 10854 26336 10906
rect 26516 10854 26518 10906
rect 26272 10852 26278 10854
rect 26334 10852 26358 10854
rect 26414 10852 26438 10854
rect 26494 10852 26518 10854
rect 26574 10852 26580 10854
rect 26272 10843 26580 10852
rect 22052 10364 22360 10373
rect 22052 10362 22058 10364
rect 22114 10362 22138 10364
rect 22194 10362 22218 10364
rect 22274 10362 22298 10364
rect 22354 10362 22360 10364
rect 22114 10310 22116 10362
rect 22296 10310 22298 10362
rect 22052 10308 22058 10310
rect 22114 10308 22138 10310
rect 22194 10308 22218 10310
rect 22274 10308 22298 10310
rect 22354 10308 22360 10310
rect 22052 10299 22360 10308
rect 26272 9820 26580 9829
rect 26272 9818 26278 9820
rect 26334 9818 26358 9820
rect 26414 9818 26438 9820
rect 26494 9818 26518 9820
rect 26574 9818 26580 9820
rect 26334 9766 26336 9818
rect 26516 9766 26518 9818
rect 26272 9764 26278 9766
rect 26334 9764 26358 9766
rect 26414 9764 26438 9766
rect 26494 9764 26518 9766
rect 26574 9764 26580 9766
rect 26272 9755 26580 9764
rect 22052 9276 22360 9285
rect 22052 9274 22058 9276
rect 22114 9274 22138 9276
rect 22194 9274 22218 9276
rect 22274 9274 22298 9276
rect 22354 9274 22360 9276
rect 22114 9222 22116 9274
rect 22296 9222 22298 9274
rect 22052 9220 22058 9222
rect 22114 9220 22138 9222
rect 22194 9220 22218 9222
rect 22274 9220 22298 9222
rect 22354 9220 22360 9222
rect 22052 9211 22360 9220
rect 26272 8732 26580 8741
rect 26272 8730 26278 8732
rect 26334 8730 26358 8732
rect 26414 8730 26438 8732
rect 26494 8730 26518 8732
rect 26574 8730 26580 8732
rect 26334 8678 26336 8730
rect 26516 8678 26518 8730
rect 26272 8676 26278 8678
rect 26334 8676 26358 8678
rect 26414 8676 26438 8678
rect 26494 8676 26518 8678
rect 26574 8676 26580 8678
rect 26272 8667 26580 8676
rect 22052 8188 22360 8197
rect 22052 8186 22058 8188
rect 22114 8186 22138 8188
rect 22194 8186 22218 8188
rect 22274 8186 22298 8188
rect 22354 8186 22360 8188
rect 22114 8134 22116 8186
rect 22296 8134 22298 8186
rect 22052 8132 22058 8134
rect 22114 8132 22138 8134
rect 22194 8132 22218 8134
rect 22274 8132 22298 8134
rect 22354 8132 22360 8134
rect 22052 8123 22360 8132
rect 26272 7644 26580 7653
rect 26272 7642 26278 7644
rect 26334 7642 26358 7644
rect 26414 7642 26438 7644
rect 26494 7642 26518 7644
rect 26574 7642 26580 7644
rect 26334 7590 26336 7642
rect 26516 7590 26518 7642
rect 26272 7588 26278 7590
rect 26334 7588 26358 7590
rect 26414 7588 26438 7590
rect 26494 7588 26518 7590
rect 26574 7588 26580 7590
rect 26272 7579 26580 7588
rect 22052 7100 22360 7109
rect 22052 7098 22058 7100
rect 22114 7098 22138 7100
rect 22194 7098 22218 7100
rect 22274 7098 22298 7100
rect 22354 7098 22360 7100
rect 22114 7046 22116 7098
rect 22296 7046 22298 7098
rect 22052 7044 22058 7046
rect 22114 7044 22138 7046
rect 22194 7044 22218 7046
rect 22274 7044 22298 7046
rect 22354 7044 22360 7046
rect 22052 7035 22360 7044
rect 19628 6886 19748 6914
rect 9390 6556 9698 6565
rect 9390 6554 9396 6556
rect 9452 6554 9476 6556
rect 9532 6554 9556 6556
rect 9612 6554 9636 6556
rect 9692 6554 9698 6556
rect 9452 6502 9454 6554
rect 9634 6502 9636 6554
rect 9390 6500 9396 6502
rect 9452 6500 9476 6502
rect 9532 6500 9556 6502
rect 9612 6500 9636 6502
rect 9692 6500 9698 6502
rect 9390 6491 9698 6500
rect 17831 6556 18139 6565
rect 17831 6554 17837 6556
rect 17893 6554 17917 6556
rect 17973 6554 17997 6556
rect 18053 6554 18077 6556
rect 18133 6554 18139 6556
rect 17893 6502 17895 6554
rect 18075 6502 18077 6554
rect 17831 6500 17837 6502
rect 17893 6500 17917 6502
rect 17973 6500 17997 6502
rect 18053 6500 18077 6502
rect 18133 6500 18139 6502
rect 17831 6491 18139 6500
rect 5170 6012 5478 6021
rect 5170 6010 5176 6012
rect 5232 6010 5256 6012
rect 5312 6010 5336 6012
rect 5392 6010 5416 6012
rect 5472 6010 5478 6012
rect 5232 5958 5234 6010
rect 5414 5958 5416 6010
rect 5170 5956 5176 5958
rect 5232 5956 5256 5958
rect 5312 5956 5336 5958
rect 5392 5956 5416 5958
rect 5472 5956 5478 5958
rect 5170 5947 5478 5956
rect 13611 6012 13919 6021
rect 13611 6010 13617 6012
rect 13673 6010 13697 6012
rect 13753 6010 13777 6012
rect 13833 6010 13857 6012
rect 13913 6010 13919 6012
rect 13673 5958 13675 6010
rect 13855 5958 13857 6010
rect 13611 5956 13617 5958
rect 13673 5956 13697 5958
rect 13753 5956 13777 5958
rect 13833 5956 13857 5958
rect 13913 5956 13919 5958
rect 13611 5947 13919 5956
rect 9390 5468 9698 5477
rect 9390 5466 9396 5468
rect 9452 5466 9476 5468
rect 9532 5466 9556 5468
rect 9612 5466 9636 5468
rect 9692 5466 9698 5468
rect 9452 5414 9454 5466
rect 9634 5414 9636 5466
rect 9390 5412 9396 5414
rect 9452 5412 9476 5414
rect 9532 5412 9556 5414
rect 9612 5412 9636 5414
rect 9692 5412 9698 5414
rect 9390 5403 9698 5412
rect 17831 5468 18139 5477
rect 17831 5466 17837 5468
rect 17893 5466 17917 5468
rect 17973 5466 17997 5468
rect 18053 5466 18077 5468
rect 18133 5466 18139 5468
rect 17893 5414 17895 5466
rect 18075 5414 18077 5466
rect 17831 5412 17837 5414
rect 17893 5412 17917 5414
rect 17973 5412 17997 5414
rect 18053 5412 18077 5414
rect 18133 5412 18139 5414
rect 17831 5403 18139 5412
rect 5170 4924 5478 4933
rect 5170 4922 5176 4924
rect 5232 4922 5256 4924
rect 5312 4922 5336 4924
rect 5392 4922 5416 4924
rect 5472 4922 5478 4924
rect 5232 4870 5234 4922
rect 5414 4870 5416 4922
rect 5170 4868 5176 4870
rect 5232 4868 5256 4870
rect 5312 4868 5336 4870
rect 5392 4868 5416 4870
rect 5472 4868 5478 4870
rect 5170 4859 5478 4868
rect 13611 4924 13919 4933
rect 13611 4922 13617 4924
rect 13673 4922 13697 4924
rect 13753 4922 13777 4924
rect 13833 4922 13857 4924
rect 13913 4922 13919 4924
rect 13673 4870 13675 4922
rect 13855 4870 13857 4922
rect 13611 4868 13617 4870
rect 13673 4868 13697 4870
rect 13753 4868 13777 4870
rect 13833 4868 13857 4870
rect 13913 4868 13919 4870
rect 13611 4859 13919 4868
rect 9390 4380 9698 4389
rect 9390 4378 9396 4380
rect 9452 4378 9476 4380
rect 9532 4378 9556 4380
rect 9612 4378 9636 4380
rect 9692 4378 9698 4380
rect 9452 4326 9454 4378
rect 9634 4326 9636 4378
rect 9390 4324 9396 4326
rect 9452 4324 9476 4326
rect 9532 4324 9556 4326
rect 9612 4324 9636 4326
rect 9692 4324 9698 4326
rect 9390 4315 9698 4324
rect 17831 4380 18139 4389
rect 17831 4378 17837 4380
rect 17893 4378 17917 4380
rect 17973 4378 17997 4380
rect 18053 4378 18077 4380
rect 18133 4378 18139 4380
rect 17893 4326 17895 4378
rect 18075 4326 18077 4378
rect 17831 4324 17837 4326
rect 17893 4324 17917 4326
rect 17973 4324 17997 4326
rect 18053 4324 18077 4326
rect 18133 4324 18139 4326
rect 17831 4315 18139 4324
rect 5170 3836 5478 3845
rect 5170 3834 5176 3836
rect 5232 3834 5256 3836
rect 5312 3834 5336 3836
rect 5392 3834 5416 3836
rect 5472 3834 5478 3836
rect 5232 3782 5234 3834
rect 5414 3782 5416 3834
rect 5170 3780 5176 3782
rect 5232 3780 5256 3782
rect 5312 3780 5336 3782
rect 5392 3780 5416 3782
rect 5472 3780 5478 3782
rect 5170 3771 5478 3780
rect 13611 3836 13919 3845
rect 13611 3834 13617 3836
rect 13673 3834 13697 3836
rect 13753 3834 13777 3836
rect 13833 3834 13857 3836
rect 13913 3834 13919 3836
rect 13673 3782 13675 3834
rect 13855 3782 13857 3834
rect 13611 3780 13617 3782
rect 13673 3780 13697 3782
rect 13753 3780 13777 3782
rect 13833 3780 13857 3782
rect 13913 3780 13919 3782
rect 13611 3771 13919 3780
rect 9390 3292 9698 3301
rect 9390 3290 9396 3292
rect 9452 3290 9476 3292
rect 9532 3290 9556 3292
rect 9612 3290 9636 3292
rect 9692 3290 9698 3292
rect 9452 3238 9454 3290
rect 9634 3238 9636 3290
rect 9390 3236 9396 3238
rect 9452 3236 9476 3238
rect 9532 3236 9556 3238
rect 9612 3236 9636 3238
rect 9692 3236 9698 3238
rect 9390 3227 9698 3236
rect 17831 3292 18139 3301
rect 17831 3290 17837 3292
rect 17893 3290 17917 3292
rect 17973 3290 17997 3292
rect 18053 3290 18077 3292
rect 18133 3290 18139 3292
rect 17893 3238 17895 3290
rect 18075 3238 18077 3290
rect 17831 3236 17837 3238
rect 17893 3236 17917 3238
rect 17973 3236 17997 3238
rect 18053 3236 18077 3238
rect 18133 3236 18139 3238
rect 17831 3227 18139 3236
rect 5170 2748 5478 2757
rect 5170 2746 5176 2748
rect 5232 2746 5256 2748
rect 5312 2746 5336 2748
rect 5392 2746 5416 2748
rect 5472 2746 5478 2748
rect 5232 2694 5234 2746
rect 5414 2694 5416 2746
rect 5170 2692 5176 2694
rect 5232 2692 5256 2694
rect 5312 2692 5336 2694
rect 5392 2692 5416 2694
rect 5472 2692 5478 2694
rect 5170 2683 5478 2692
rect 13611 2748 13919 2757
rect 13611 2746 13617 2748
rect 13673 2746 13697 2748
rect 13753 2746 13777 2748
rect 13833 2746 13857 2748
rect 13913 2746 13919 2748
rect 13673 2694 13675 2746
rect 13855 2694 13857 2746
rect 13611 2692 13617 2694
rect 13673 2692 13697 2694
rect 13753 2692 13777 2694
rect 13833 2692 13857 2694
rect 13913 2692 13919 2694
rect 13611 2683 13919 2692
rect 1676 2508 1728 2514
rect 1676 2450 1728 2456
rect 19628 2446 19656 6886
rect 26272 6556 26580 6565
rect 26272 6554 26278 6556
rect 26334 6554 26358 6556
rect 26414 6554 26438 6556
rect 26494 6554 26518 6556
rect 26574 6554 26580 6556
rect 26334 6502 26336 6554
rect 26516 6502 26518 6554
rect 26272 6500 26278 6502
rect 26334 6500 26358 6502
rect 26414 6500 26438 6502
rect 26494 6500 26518 6502
rect 26574 6500 26580 6502
rect 26272 6491 26580 6500
rect 22052 6012 22360 6021
rect 22052 6010 22058 6012
rect 22114 6010 22138 6012
rect 22194 6010 22218 6012
rect 22274 6010 22298 6012
rect 22354 6010 22360 6012
rect 22114 5958 22116 6010
rect 22296 5958 22298 6010
rect 22052 5956 22058 5958
rect 22114 5956 22138 5958
rect 22194 5956 22218 5958
rect 22274 5956 22298 5958
rect 22354 5956 22360 5958
rect 22052 5947 22360 5956
rect 26272 5468 26580 5477
rect 26272 5466 26278 5468
rect 26334 5466 26358 5468
rect 26414 5466 26438 5468
rect 26494 5466 26518 5468
rect 26574 5466 26580 5468
rect 26334 5414 26336 5466
rect 26516 5414 26518 5466
rect 26272 5412 26278 5414
rect 26334 5412 26358 5414
rect 26414 5412 26438 5414
rect 26494 5412 26518 5414
rect 26574 5412 26580 5414
rect 26272 5403 26580 5412
rect 22052 4924 22360 4933
rect 22052 4922 22058 4924
rect 22114 4922 22138 4924
rect 22194 4922 22218 4924
rect 22274 4922 22298 4924
rect 22354 4922 22360 4924
rect 22114 4870 22116 4922
rect 22296 4870 22298 4922
rect 22052 4868 22058 4870
rect 22114 4868 22138 4870
rect 22194 4868 22218 4870
rect 22274 4868 22298 4870
rect 22354 4868 22360 4870
rect 22052 4859 22360 4868
rect 26272 4380 26580 4389
rect 26272 4378 26278 4380
rect 26334 4378 26358 4380
rect 26414 4378 26438 4380
rect 26494 4378 26518 4380
rect 26574 4378 26580 4380
rect 26334 4326 26336 4378
rect 26516 4326 26518 4378
rect 26272 4324 26278 4326
rect 26334 4324 26358 4326
rect 26414 4324 26438 4326
rect 26494 4324 26518 4326
rect 26574 4324 26580 4326
rect 26272 4315 26580 4324
rect 22052 3836 22360 3845
rect 22052 3834 22058 3836
rect 22114 3834 22138 3836
rect 22194 3834 22218 3836
rect 22274 3834 22298 3836
rect 22354 3834 22360 3836
rect 22114 3782 22116 3834
rect 22296 3782 22298 3834
rect 22052 3780 22058 3782
rect 22114 3780 22138 3782
rect 22194 3780 22218 3782
rect 22274 3780 22298 3782
rect 22354 3780 22360 3782
rect 22052 3771 22360 3780
rect 26272 3292 26580 3301
rect 26272 3290 26278 3292
rect 26334 3290 26358 3292
rect 26414 3290 26438 3292
rect 26494 3290 26518 3292
rect 26574 3290 26580 3292
rect 26334 3238 26336 3290
rect 26516 3238 26518 3290
rect 26272 3236 26278 3238
rect 26334 3236 26358 3238
rect 26414 3236 26438 3238
rect 26494 3236 26518 3238
rect 26574 3236 26580 3238
rect 26272 3227 26580 3236
rect 22052 2748 22360 2757
rect 22052 2746 22058 2748
rect 22114 2746 22138 2748
rect 22194 2746 22218 2748
rect 22274 2746 22298 2748
rect 22354 2746 22360 2748
rect 22114 2694 22116 2746
rect 22296 2694 22298 2746
rect 22052 2692 22058 2694
rect 22114 2692 22138 2694
rect 22194 2692 22218 2694
rect 22274 2692 22298 2694
rect 22354 2692 22360 2694
rect 22052 2683 22360 2692
rect 28460 2650 28488 14350
rect 30493 13628 30801 13637
rect 30493 13626 30499 13628
rect 30555 13626 30579 13628
rect 30635 13626 30659 13628
rect 30715 13626 30739 13628
rect 30795 13626 30801 13628
rect 30555 13574 30557 13626
rect 30737 13574 30739 13626
rect 30493 13572 30499 13574
rect 30555 13572 30579 13574
rect 30635 13572 30659 13574
rect 30715 13572 30739 13574
rect 30795 13572 30801 13574
rect 30493 13563 30801 13572
rect 30493 12540 30801 12549
rect 30493 12538 30499 12540
rect 30555 12538 30579 12540
rect 30635 12538 30659 12540
rect 30715 12538 30739 12540
rect 30795 12538 30801 12540
rect 30555 12486 30557 12538
rect 30737 12486 30739 12538
rect 30493 12484 30499 12486
rect 30555 12484 30579 12486
rect 30635 12484 30659 12486
rect 30715 12484 30739 12486
rect 30795 12484 30801 12486
rect 30493 12475 30801 12484
rect 30493 11452 30801 11461
rect 30493 11450 30499 11452
rect 30555 11450 30579 11452
rect 30635 11450 30659 11452
rect 30715 11450 30739 11452
rect 30795 11450 30801 11452
rect 30555 11398 30557 11450
rect 30737 11398 30739 11450
rect 30493 11396 30499 11398
rect 30555 11396 30579 11398
rect 30635 11396 30659 11398
rect 30715 11396 30739 11398
rect 30795 11396 30801 11398
rect 30493 11387 30801 11396
rect 30493 10364 30801 10373
rect 30493 10362 30499 10364
rect 30555 10362 30579 10364
rect 30635 10362 30659 10364
rect 30715 10362 30739 10364
rect 30795 10362 30801 10364
rect 30555 10310 30557 10362
rect 30737 10310 30739 10362
rect 30493 10308 30499 10310
rect 30555 10308 30579 10310
rect 30635 10308 30659 10310
rect 30715 10308 30739 10310
rect 30795 10308 30801 10310
rect 30493 10299 30801 10308
rect 30493 9276 30801 9285
rect 30493 9274 30499 9276
rect 30555 9274 30579 9276
rect 30635 9274 30659 9276
rect 30715 9274 30739 9276
rect 30795 9274 30801 9276
rect 30555 9222 30557 9274
rect 30737 9222 30739 9274
rect 30493 9220 30499 9222
rect 30555 9220 30579 9222
rect 30635 9220 30659 9222
rect 30715 9220 30739 9222
rect 30795 9220 30801 9222
rect 30493 9211 30801 9220
rect 30493 8188 30801 8197
rect 30493 8186 30499 8188
rect 30555 8186 30579 8188
rect 30635 8186 30659 8188
rect 30715 8186 30739 8188
rect 30795 8186 30801 8188
rect 30555 8134 30557 8186
rect 30737 8134 30739 8186
rect 30493 8132 30499 8134
rect 30555 8132 30579 8134
rect 30635 8132 30659 8134
rect 30715 8132 30739 8134
rect 30795 8132 30801 8134
rect 30493 8123 30801 8132
rect 30493 7100 30801 7109
rect 30493 7098 30499 7100
rect 30555 7098 30579 7100
rect 30635 7098 30659 7100
rect 30715 7098 30739 7100
rect 30795 7098 30801 7100
rect 30555 7046 30557 7098
rect 30737 7046 30739 7098
rect 30493 7044 30499 7046
rect 30555 7044 30579 7046
rect 30635 7044 30659 7046
rect 30715 7044 30739 7046
rect 30795 7044 30801 7046
rect 30493 7035 30801 7044
rect 30493 6012 30801 6021
rect 30493 6010 30499 6012
rect 30555 6010 30579 6012
rect 30635 6010 30659 6012
rect 30715 6010 30739 6012
rect 30795 6010 30801 6012
rect 30555 5958 30557 6010
rect 30737 5958 30739 6010
rect 30493 5956 30499 5958
rect 30555 5956 30579 5958
rect 30635 5956 30659 5958
rect 30715 5956 30739 5958
rect 30795 5956 30801 5958
rect 30493 5947 30801 5956
rect 30493 4924 30801 4933
rect 30493 4922 30499 4924
rect 30555 4922 30579 4924
rect 30635 4922 30659 4924
rect 30715 4922 30739 4924
rect 30795 4922 30801 4924
rect 30555 4870 30557 4922
rect 30737 4870 30739 4922
rect 30493 4868 30499 4870
rect 30555 4868 30579 4870
rect 30635 4868 30659 4870
rect 30715 4868 30739 4870
rect 30795 4868 30801 4870
rect 30493 4859 30801 4868
rect 30493 3836 30801 3845
rect 30493 3834 30499 3836
rect 30555 3834 30579 3836
rect 30635 3834 30659 3836
rect 30715 3834 30739 3836
rect 30795 3834 30801 3836
rect 30555 3782 30557 3834
rect 30737 3782 30739 3834
rect 30493 3780 30499 3782
rect 30555 3780 30579 3782
rect 30635 3780 30659 3782
rect 30715 3780 30739 3782
rect 30795 3780 30801 3782
rect 30493 3771 30801 3780
rect 30493 2748 30801 2757
rect 30493 2746 30499 2748
rect 30555 2746 30579 2748
rect 30635 2746 30659 2748
rect 30715 2746 30739 2748
rect 30795 2746 30801 2748
rect 30555 2694 30557 2746
rect 30737 2694 30739 2746
rect 30493 2692 30499 2694
rect 30555 2692 30579 2694
rect 30635 2692 30659 2694
rect 30715 2692 30739 2694
rect 30795 2692 30801 2694
rect 30493 2683 30801 2692
rect 31496 2650 31524 14962
rect 34713 14172 35021 14181
rect 34713 14170 34719 14172
rect 34775 14170 34799 14172
rect 34855 14170 34879 14172
rect 34935 14170 34959 14172
rect 35015 14170 35021 14172
rect 34775 14118 34777 14170
rect 34957 14118 34959 14170
rect 34713 14116 34719 14118
rect 34775 14116 34799 14118
rect 34855 14116 34879 14118
rect 34935 14116 34959 14118
rect 35015 14116 35021 14118
rect 34713 14107 35021 14116
rect 34713 13084 35021 13093
rect 34713 13082 34719 13084
rect 34775 13082 34799 13084
rect 34855 13082 34879 13084
rect 34935 13082 34959 13084
rect 35015 13082 35021 13084
rect 34775 13030 34777 13082
rect 34957 13030 34959 13082
rect 34713 13028 34719 13030
rect 34775 13028 34799 13030
rect 34855 13028 34879 13030
rect 34935 13028 34959 13030
rect 35015 13028 35021 13030
rect 34713 13019 35021 13028
rect 34152 12096 34204 12102
rect 34152 12038 34204 12044
rect 34164 11898 34192 12038
rect 34713 11996 35021 12005
rect 34713 11994 34719 11996
rect 34775 11994 34799 11996
rect 34855 11994 34879 11996
rect 34935 11994 34959 11996
rect 35015 11994 35021 11996
rect 34775 11942 34777 11994
rect 34957 11942 34959 11994
rect 34713 11940 34719 11942
rect 34775 11940 34799 11942
rect 34855 11940 34879 11942
rect 34935 11940 34959 11942
rect 35015 11940 35021 11942
rect 34713 11931 35021 11940
rect 34152 11892 34204 11898
rect 34152 11834 34204 11840
rect 34518 11656 34574 11665
rect 34518 11591 34520 11600
rect 34572 11591 34574 11600
rect 34520 11562 34572 11568
rect 34713 10908 35021 10917
rect 34713 10906 34719 10908
rect 34775 10906 34799 10908
rect 34855 10906 34879 10908
rect 34935 10906 34959 10908
rect 35015 10906 35021 10908
rect 34775 10854 34777 10906
rect 34957 10854 34959 10906
rect 34713 10852 34719 10854
rect 34775 10852 34799 10854
rect 34855 10852 34879 10854
rect 34935 10852 34959 10854
rect 35015 10852 35021 10854
rect 34713 10843 35021 10852
rect 34713 9820 35021 9829
rect 34713 9818 34719 9820
rect 34775 9818 34799 9820
rect 34855 9818 34879 9820
rect 34935 9818 34959 9820
rect 35015 9818 35021 9820
rect 34775 9766 34777 9818
rect 34957 9766 34959 9818
rect 34713 9764 34719 9766
rect 34775 9764 34799 9766
rect 34855 9764 34879 9766
rect 34935 9764 34959 9766
rect 35015 9764 35021 9766
rect 34713 9755 35021 9764
rect 34713 8732 35021 8741
rect 34713 8730 34719 8732
rect 34775 8730 34799 8732
rect 34855 8730 34879 8732
rect 34935 8730 34959 8732
rect 35015 8730 35021 8732
rect 34775 8678 34777 8730
rect 34957 8678 34959 8730
rect 34713 8676 34719 8678
rect 34775 8676 34799 8678
rect 34855 8676 34879 8678
rect 34935 8676 34959 8678
rect 35015 8676 35021 8678
rect 34713 8667 35021 8676
rect 34713 7644 35021 7653
rect 34713 7642 34719 7644
rect 34775 7642 34799 7644
rect 34855 7642 34879 7644
rect 34935 7642 34959 7644
rect 35015 7642 35021 7644
rect 34775 7590 34777 7642
rect 34957 7590 34959 7642
rect 34713 7588 34719 7590
rect 34775 7588 34799 7590
rect 34855 7588 34879 7590
rect 34935 7588 34959 7590
rect 35015 7588 35021 7590
rect 34713 7579 35021 7588
rect 34713 6556 35021 6565
rect 34713 6554 34719 6556
rect 34775 6554 34799 6556
rect 34855 6554 34879 6556
rect 34935 6554 34959 6556
rect 35015 6554 35021 6556
rect 34775 6502 34777 6554
rect 34957 6502 34959 6554
rect 34713 6500 34719 6502
rect 34775 6500 34799 6502
rect 34855 6500 34879 6502
rect 34935 6500 34959 6502
rect 35015 6500 35021 6502
rect 34713 6491 35021 6500
rect 34713 5468 35021 5477
rect 34713 5466 34719 5468
rect 34775 5466 34799 5468
rect 34855 5466 34879 5468
rect 34935 5466 34959 5468
rect 35015 5466 35021 5468
rect 34775 5414 34777 5466
rect 34957 5414 34959 5466
rect 34713 5412 34719 5414
rect 34775 5412 34799 5414
rect 34855 5412 34879 5414
rect 34935 5412 34959 5414
rect 35015 5412 35021 5414
rect 34713 5403 35021 5412
rect 34713 4380 35021 4389
rect 34713 4378 34719 4380
rect 34775 4378 34799 4380
rect 34855 4378 34879 4380
rect 34935 4378 34959 4380
rect 35015 4378 35021 4380
rect 34775 4326 34777 4378
rect 34957 4326 34959 4378
rect 34713 4324 34719 4326
rect 34775 4324 34799 4326
rect 34855 4324 34879 4326
rect 34935 4324 34959 4326
rect 35015 4324 35021 4326
rect 34713 4315 35021 4324
rect 34713 3292 35021 3301
rect 34713 3290 34719 3292
rect 34775 3290 34799 3292
rect 34855 3290 34879 3292
rect 34935 3290 34959 3292
rect 35015 3290 35021 3292
rect 34775 3238 34777 3290
rect 34957 3238 34959 3290
rect 34713 3236 34719 3238
rect 34775 3236 34799 3238
rect 34855 3236 34879 3238
rect 34935 3236 34959 3238
rect 35015 3236 35021 3238
rect 34713 3227 35021 3236
rect 28448 2644 28500 2650
rect 28448 2586 28500 2592
rect 31484 2644 31536 2650
rect 31484 2586 31536 2592
rect 20 2440 72 2446
rect 20 2382 72 2388
rect 9128 2440 9180 2446
rect 9128 2382 9180 2388
rect 19616 2440 19668 2446
rect 19616 2382 19668 2388
rect 28356 2440 28408 2446
rect 28356 2382 28408 2388
rect 32 800 60 2382
rect 9140 1306 9168 2382
rect 18788 2304 18840 2310
rect 18788 2246 18840 2252
rect 9390 2204 9698 2213
rect 9390 2202 9396 2204
rect 9452 2202 9476 2204
rect 9532 2202 9556 2204
rect 9612 2202 9636 2204
rect 9692 2202 9698 2204
rect 9452 2150 9454 2202
rect 9634 2150 9636 2202
rect 9390 2148 9396 2150
rect 9452 2148 9476 2150
rect 9532 2148 9556 2150
rect 9612 2148 9636 2150
rect 9692 2148 9698 2150
rect 9390 2139 9698 2148
rect 17831 2204 18139 2213
rect 17831 2202 17837 2204
rect 17893 2202 17917 2204
rect 17973 2202 17997 2204
rect 18053 2202 18077 2204
rect 18133 2202 18139 2204
rect 17893 2150 17895 2202
rect 18075 2150 18077 2202
rect 17831 2148 17837 2150
rect 17893 2148 17917 2150
rect 17973 2148 17997 2150
rect 18053 2148 18077 2150
rect 18133 2148 18139 2150
rect 17831 2139 18139 2148
rect 9048 1278 9168 1306
rect 9048 800 9076 1278
rect 18800 1170 18828 2246
rect 26272 2204 26580 2213
rect 26272 2202 26278 2204
rect 26334 2202 26358 2204
rect 26414 2202 26438 2204
rect 26494 2202 26518 2204
rect 26574 2202 26580 2204
rect 26334 2150 26336 2202
rect 26516 2150 26518 2202
rect 26272 2148 26278 2150
rect 26334 2148 26358 2150
rect 26414 2148 26438 2150
rect 26494 2148 26518 2150
rect 26574 2148 26580 2150
rect 26272 2139 26580 2148
rect 18708 1142 18828 1170
rect 18708 800 18736 1142
rect 28368 800 28396 2382
rect 35164 2304 35216 2310
rect 35164 2246 35216 2252
rect 34713 2204 35021 2213
rect 34713 2202 34719 2204
rect 34775 2202 34799 2204
rect 34855 2202 34879 2204
rect 34935 2202 34959 2204
rect 35015 2202 35021 2204
rect 34775 2150 34777 2202
rect 34957 2150 34959 2202
rect 34713 2148 34719 2150
rect 34775 2148 34799 2150
rect 34855 2148 34879 2150
rect 34935 2148 34959 2150
rect 35015 2148 35021 2150
rect 34713 2139 35021 2148
rect 35176 2145 35204 2246
rect 35162 2136 35218 2145
rect 35162 2071 35218 2080
rect -10 0 102 800
rect 9006 0 9118 800
rect 18666 0 18778 800
rect 28326 0 28438 800
<< via2 >>
rect 5176 39738 5232 39740
rect 5256 39738 5312 39740
rect 5336 39738 5392 39740
rect 5416 39738 5472 39740
rect 5176 39686 5222 39738
rect 5222 39686 5232 39738
rect 5256 39686 5286 39738
rect 5286 39686 5298 39738
rect 5298 39686 5312 39738
rect 5336 39686 5350 39738
rect 5350 39686 5362 39738
rect 5362 39686 5392 39738
rect 5416 39686 5426 39738
rect 5426 39686 5472 39738
rect 5176 39684 5232 39686
rect 5256 39684 5312 39686
rect 5336 39684 5392 39686
rect 5416 39684 5472 39686
rect 938 39480 994 39536
rect 13617 39738 13673 39740
rect 13697 39738 13753 39740
rect 13777 39738 13833 39740
rect 13857 39738 13913 39740
rect 13617 39686 13663 39738
rect 13663 39686 13673 39738
rect 13697 39686 13727 39738
rect 13727 39686 13739 39738
rect 13739 39686 13753 39738
rect 13777 39686 13791 39738
rect 13791 39686 13803 39738
rect 13803 39686 13833 39738
rect 13857 39686 13867 39738
rect 13867 39686 13913 39738
rect 13617 39684 13673 39686
rect 13697 39684 13753 39686
rect 13777 39684 13833 39686
rect 13857 39684 13913 39686
rect 22058 39738 22114 39740
rect 22138 39738 22194 39740
rect 22218 39738 22274 39740
rect 22298 39738 22354 39740
rect 22058 39686 22104 39738
rect 22104 39686 22114 39738
rect 22138 39686 22168 39738
rect 22168 39686 22180 39738
rect 22180 39686 22194 39738
rect 22218 39686 22232 39738
rect 22232 39686 22244 39738
rect 22244 39686 22274 39738
rect 22298 39686 22308 39738
rect 22308 39686 22354 39738
rect 22058 39684 22114 39686
rect 22138 39684 22194 39686
rect 22218 39684 22274 39686
rect 22298 39684 22354 39686
rect 30499 39738 30555 39740
rect 30579 39738 30635 39740
rect 30659 39738 30715 39740
rect 30739 39738 30795 39740
rect 30499 39686 30545 39738
rect 30545 39686 30555 39738
rect 30579 39686 30609 39738
rect 30609 39686 30621 39738
rect 30621 39686 30635 39738
rect 30659 39686 30673 39738
rect 30673 39686 30685 39738
rect 30685 39686 30715 39738
rect 30739 39686 30749 39738
rect 30749 39686 30795 39738
rect 30499 39684 30555 39686
rect 30579 39684 30635 39686
rect 30659 39684 30715 39686
rect 30739 39684 30795 39686
rect 9396 39194 9452 39196
rect 9476 39194 9532 39196
rect 9556 39194 9612 39196
rect 9636 39194 9692 39196
rect 9396 39142 9442 39194
rect 9442 39142 9452 39194
rect 9476 39142 9506 39194
rect 9506 39142 9518 39194
rect 9518 39142 9532 39194
rect 9556 39142 9570 39194
rect 9570 39142 9582 39194
rect 9582 39142 9612 39194
rect 9636 39142 9646 39194
rect 9646 39142 9692 39194
rect 9396 39140 9452 39142
rect 9476 39140 9532 39142
rect 9556 39140 9612 39142
rect 9636 39140 9692 39142
rect 5176 38650 5232 38652
rect 5256 38650 5312 38652
rect 5336 38650 5392 38652
rect 5416 38650 5472 38652
rect 5176 38598 5222 38650
rect 5222 38598 5232 38650
rect 5256 38598 5286 38650
rect 5286 38598 5298 38650
rect 5298 38598 5312 38650
rect 5336 38598 5350 38650
rect 5350 38598 5362 38650
rect 5362 38598 5392 38650
rect 5416 38598 5426 38650
rect 5426 38598 5472 38650
rect 5176 38596 5232 38598
rect 5256 38596 5312 38598
rect 5336 38596 5392 38598
rect 5416 38596 5472 38598
rect 13617 38650 13673 38652
rect 13697 38650 13753 38652
rect 13777 38650 13833 38652
rect 13857 38650 13913 38652
rect 13617 38598 13663 38650
rect 13663 38598 13673 38650
rect 13697 38598 13727 38650
rect 13727 38598 13739 38650
rect 13739 38598 13753 38650
rect 13777 38598 13791 38650
rect 13791 38598 13803 38650
rect 13803 38598 13833 38650
rect 13857 38598 13867 38650
rect 13867 38598 13913 38650
rect 13617 38596 13673 38598
rect 13697 38596 13753 38598
rect 13777 38596 13833 38598
rect 13857 38596 13913 38598
rect 9396 38106 9452 38108
rect 9476 38106 9532 38108
rect 9556 38106 9612 38108
rect 9636 38106 9692 38108
rect 9396 38054 9442 38106
rect 9442 38054 9452 38106
rect 9476 38054 9506 38106
rect 9506 38054 9518 38106
rect 9518 38054 9532 38106
rect 9556 38054 9570 38106
rect 9570 38054 9582 38106
rect 9582 38054 9612 38106
rect 9636 38054 9646 38106
rect 9646 38054 9692 38106
rect 9396 38052 9452 38054
rect 9476 38052 9532 38054
rect 9556 38052 9612 38054
rect 9636 38052 9692 38054
rect 5176 37562 5232 37564
rect 5256 37562 5312 37564
rect 5336 37562 5392 37564
rect 5416 37562 5472 37564
rect 5176 37510 5222 37562
rect 5222 37510 5232 37562
rect 5256 37510 5286 37562
rect 5286 37510 5298 37562
rect 5298 37510 5312 37562
rect 5336 37510 5350 37562
rect 5350 37510 5362 37562
rect 5362 37510 5392 37562
rect 5416 37510 5426 37562
rect 5426 37510 5472 37562
rect 5176 37508 5232 37510
rect 5256 37508 5312 37510
rect 5336 37508 5392 37510
rect 5416 37508 5472 37510
rect 13617 37562 13673 37564
rect 13697 37562 13753 37564
rect 13777 37562 13833 37564
rect 13857 37562 13913 37564
rect 13617 37510 13663 37562
rect 13663 37510 13673 37562
rect 13697 37510 13727 37562
rect 13727 37510 13739 37562
rect 13739 37510 13753 37562
rect 13777 37510 13791 37562
rect 13791 37510 13803 37562
rect 13803 37510 13833 37562
rect 13857 37510 13867 37562
rect 13867 37510 13913 37562
rect 13617 37508 13673 37510
rect 13697 37508 13753 37510
rect 13777 37508 13833 37510
rect 13857 37508 13913 37510
rect 9396 37018 9452 37020
rect 9476 37018 9532 37020
rect 9556 37018 9612 37020
rect 9636 37018 9692 37020
rect 9396 36966 9442 37018
rect 9442 36966 9452 37018
rect 9476 36966 9506 37018
rect 9506 36966 9518 37018
rect 9518 36966 9532 37018
rect 9556 36966 9570 37018
rect 9570 36966 9582 37018
rect 9582 36966 9612 37018
rect 9636 36966 9646 37018
rect 9646 36966 9692 37018
rect 9396 36964 9452 36966
rect 9476 36964 9532 36966
rect 9556 36964 9612 36966
rect 9636 36964 9692 36966
rect 5176 36474 5232 36476
rect 5256 36474 5312 36476
rect 5336 36474 5392 36476
rect 5416 36474 5472 36476
rect 5176 36422 5222 36474
rect 5222 36422 5232 36474
rect 5256 36422 5286 36474
rect 5286 36422 5298 36474
rect 5298 36422 5312 36474
rect 5336 36422 5350 36474
rect 5350 36422 5362 36474
rect 5362 36422 5392 36474
rect 5416 36422 5426 36474
rect 5426 36422 5472 36474
rect 5176 36420 5232 36422
rect 5256 36420 5312 36422
rect 5336 36420 5392 36422
rect 5416 36420 5472 36422
rect 13617 36474 13673 36476
rect 13697 36474 13753 36476
rect 13777 36474 13833 36476
rect 13857 36474 13913 36476
rect 13617 36422 13663 36474
rect 13663 36422 13673 36474
rect 13697 36422 13727 36474
rect 13727 36422 13739 36474
rect 13739 36422 13753 36474
rect 13777 36422 13791 36474
rect 13791 36422 13803 36474
rect 13803 36422 13833 36474
rect 13857 36422 13867 36474
rect 13867 36422 13913 36474
rect 13617 36420 13673 36422
rect 13697 36420 13753 36422
rect 13777 36420 13833 36422
rect 13857 36420 13913 36422
rect 9396 35930 9452 35932
rect 9476 35930 9532 35932
rect 9556 35930 9612 35932
rect 9636 35930 9692 35932
rect 9396 35878 9442 35930
rect 9442 35878 9452 35930
rect 9476 35878 9506 35930
rect 9506 35878 9518 35930
rect 9518 35878 9532 35930
rect 9556 35878 9570 35930
rect 9570 35878 9582 35930
rect 9582 35878 9612 35930
rect 9636 35878 9646 35930
rect 9646 35878 9692 35930
rect 9396 35876 9452 35878
rect 9476 35876 9532 35878
rect 9556 35876 9612 35878
rect 9636 35876 9692 35878
rect 5176 35386 5232 35388
rect 5256 35386 5312 35388
rect 5336 35386 5392 35388
rect 5416 35386 5472 35388
rect 5176 35334 5222 35386
rect 5222 35334 5232 35386
rect 5256 35334 5286 35386
rect 5286 35334 5298 35386
rect 5298 35334 5312 35386
rect 5336 35334 5350 35386
rect 5350 35334 5362 35386
rect 5362 35334 5392 35386
rect 5416 35334 5426 35386
rect 5426 35334 5472 35386
rect 5176 35332 5232 35334
rect 5256 35332 5312 35334
rect 5336 35332 5392 35334
rect 5416 35332 5472 35334
rect 13617 35386 13673 35388
rect 13697 35386 13753 35388
rect 13777 35386 13833 35388
rect 13857 35386 13913 35388
rect 13617 35334 13663 35386
rect 13663 35334 13673 35386
rect 13697 35334 13727 35386
rect 13727 35334 13739 35386
rect 13739 35334 13753 35386
rect 13777 35334 13791 35386
rect 13791 35334 13803 35386
rect 13803 35334 13833 35386
rect 13857 35334 13867 35386
rect 13867 35334 13913 35386
rect 13617 35332 13673 35334
rect 13697 35332 13753 35334
rect 13777 35332 13833 35334
rect 13857 35332 13913 35334
rect 9396 34842 9452 34844
rect 9476 34842 9532 34844
rect 9556 34842 9612 34844
rect 9636 34842 9692 34844
rect 9396 34790 9442 34842
rect 9442 34790 9452 34842
rect 9476 34790 9506 34842
rect 9506 34790 9518 34842
rect 9518 34790 9532 34842
rect 9556 34790 9570 34842
rect 9570 34790 9582 34842
rect 9582 34790 9612 34842
rect 9636 34790 9646 34842
rect 9646 34790 9692 34842
rect 9396 34788 9452 34790
rect 9476 34788 9532 34790
rect 9556 34788 9612 34790
rect 9636 34788 9692 34790
rect 5176 34298 5232 34300
rect 5256 34298 5312 34300
rect 5336 34298 5392 34300
rect 5416 34298 5472 34300
rect 5176 34246 5222 34298
rect 5222 34246 5232 34298
rect 5256 34246 5286 34298
rect 5286 34246 5298 34298
rect 5298 34246 5312 34298
rect 5336 34246 5350 34298
rect 5350 34246 5362 34298
rect 5362 34246 5392 34298
rect 5416 34246 5426 34298
rect 5426 34246 5472 34298
rect 5176 34244 5232 34246
rect 5256 34244 5312 34246
rect 5336 34244 5392 34246
rect 5416 34244 5472 34246
rect 13617 34298 13673 34300
rect 13697 34298 13753 34300
rect 13777 34298 13833 34300
rect 13857 34298 13913 34300
rect 13617 34246 13663 34298
rect 13663 34246 13673 34298
rect 13697 34246 13727 34298
rect 13727 34246 13739 34298
rect 13739 34246 13753 34298
rect 13777 34246 13791 34298
rect 13791 34246 13803 34298
rect 13803 34246 13833 34298
rect 13857 34246 13867 34298
rect 13867 34246 13913 34298
rect 13617 34244 13673 34246
rect 13697 34244 13753 34246
rect 13777 34244 13833 34246
rect 13857 34244 13913 34246
rect 9396 33754 9452 33756
rect 9476 33754 9532 33756
rect 9556 33754 9612 33756
rect 9636 33754 9692 33756
rect 9396 33702 9442 33754
rect 9442 33702 9452 33754
rect 9476 33702 9506 33754
rect 9506 33702 9518 33754
rect 9518 33702 9532 33754
rect 9556 33702 9570 33754
rect 9570 33702 9582 33754
rect 9582 33702 9612 33754
rect 9636 33702 9646 33754
rect 9646 33702 9692 33754
rect 9396 33700 9452 33702
rect 9476 33700 9532 33702
rect 9556 33700 9612 33702
rect 9636 33700 9692 33702
rect 5176 33210 5232 33212
rect 5256 33210 5312 33212
rect 5336 33210 5392 33212
rect 5416 33210 5472 33212
rect 5176 33158 5222 33210
rect 5222 33158 5232 33210
rect 5256 33158 5286 33210
rect 5286 33158 5298 33210
rect 5298 33158 5312 33210
rect 5336 33158 5350 33210
rect 5350 33158 5362 33210
rect 5362 33158 5392 33210
rect 5416 33158 5426 33210
rect 5426 33158 5472 33210
rect 5176 33156 5232 33158
rect 5256 33156 5312 33158
rect 5336 33156 5392 33158
rect 5416 33156 5472 33158
rect 13617 33210 13673 33212
rect 13697 33210 13753 33212
rect 13777 33210 13833 33212
rect 13857 33210 13913 33212
rect 13617 33158 13663 33210
rect 13663 33158 13673 33210
rect 13697 33158 13727 33210
rect 13727 33158 13739 33210
rect 13739 33158 13753 33210
rect 13777 33158 13791 33210
rect 13791 33158 13803 33210
rect 13803 33158 13833 33210
rect 13857 33158 13867 33210
rect 13867 33158 13913 33210
rect 13617 33156 13673 33158
rect 13697 33156 13753 33158
rect 13777 33156 13833 33158
rect 13857 33156 13913 33158
rect 9396 32666 9452 32668
rect 9476 32666 9532 32668
rect 9556 32666 9612 32668
rect 9636 32666 9692 32668
rect 9396 32614 9442 32666
rect 9442 32614 9452 32666
rect 9476 32614 9506 32666
rect 9506 32614 9518 32666
rect 9518 32614 9532 32666
rect 9556 32614 9570 32666
rect 9570 32614 9582 32666
rect 9582 32614 9612 32666
rect 9636 32614 9646 32666
rect 9646 32614 9692 32666
rect 9396 32612 9452 32614
rect 9476 32612 9532 32614
rect 9556 32612 9612 32614
rect 9636 32612 9692 32614
rect 5176 32122 5232 32124
rect 5256 32122 5312 32124
rect 5336 32122 5392 32124
rect 5416 32122 5472 32124
rect 5176 32070 5222 32122
rect 5222 32070 5232 32122
rect 5256 32070 5286 32122
rect 5286 32070 5298 32122
rect 5298 32070 5312 32122
rect 5336 32070 5350 32122
rect 5350 32070 5362 32122
rect 5362 32070 5392 32122
rect 5416 32070 5426 32122
rect 5426 32070 5472 32122
rect 5176 32068 5232 32070
rect 5256 32068 5312 32070
rect 5336 32068 5392 32070
rect 5416 32068 5472 32070
rect 13617 32122 13673 32124
rect 13697 32122 13753 32124
rect 13777 32122 13833 32124
rect 13857 32122 13913 32124
rect 13617 32070 13663 32122
rect 13663 32070 13673 32122
rect 13697 32070 13727 32122
rect 13727 32070 13739 32122
rect 13739 32070 13753 32122
rect 13777 32070 13791 32122
rect 13791 32070 13803 32122
rect 13803 32070 13833 32122
rect 13857 32070 13867 32122
rect 13867 32070 13913 32122
rect 13617 32068 13673 32070
rect 13697 32068 13753 32070
rect 13777 32068 13833 32070
rect 13857 32068 13913 32070
rect 9396 31578 9452 31580
rect 9476 31578 9532 31580
rect 9556 31578 9612 31580
rect 9636 31578 9692 31580
rect 9396 31526 9442 31578
rect 9442 31526 9452 31578
rect 9476 31526 9506 31578
rect 9506 31526 9518 31578
rect 9518 31526 9532 31578
rect 9556 31526 9570 31578
rect 9570 31526 9582 31578
rect 9582 31526 9612 31578
rect 9636 31526 9646 31578
rect 9646 31526 9692 31578
rect 9396 31524 9452 31526
rect 9476 31524 9532 31526
rect 9556 31524 9612 31526
rect 9636 31524 9692 31526
rect 5176 31034 5232 31036
rect 5256 31034 5312 31036
rect 5336 31034 5392 31036
rect 5416 31034 5472 31036
rect 5176 30982 5222 31034
rect 5222 30982 5232 31034
rect 5256 30982 5286 31034
rect 5286 30982 5298 31034
rect 5298 30982 5312 31034
rect 5336 30982 5350 31034
rect 5350 30982 5362 31034
rect 5362 30982 5392 31034
rect 5416 30982 5426 31034
rect 5426 30982 5472 31034
rect 5176 30980 5232 30982
rect 5256 30980 5312 30982
rect 5336 30980 5392 30982
rect 5416 30980 5472 30982
rect 13617 31034 13673 31036
rect 13697 31034 13753 31036
rect 13777 31034 13833 31036
rect 13857 31034 13913 31036
rect 13617 30982 13663 31034
rect 13663 30982 13673 31034
rect 13697 30982 13727 31034
rect 13727 30982 13739 31034
rect 13739 30982 13753 31034
rect 13777 30982 13791 31034
rect 13791 30982 13803 31034
rect 13803 30982 13833 31034
rect 13857 30982 13867 31034
rect 13867 30982 13913 31034
rect 13617 30980 13673 30982
rect 13697 30980 13753 30982
rect 13777 30980 13833 30982
rect 13857 30980 13913 30982
rect 9396 30490 9452 30492
rect 9476 30490 9532 30492
rect 9556 30490 9612 30492
rect 9636 30490 9692 30492
rect 9396 30438 9442 30490
rect 9442 30438 9452 30490
rect 9476 30438 9506 30490
rect 9506 30438 9518 30490
rect 9518 30438 9532 30490
rect 9556 30438 9570 30490
rect 9570 30438 9582 30490
rect 9582 30438 9612 30490
rect 9636 30438 9646 30490
rect 9646 30438 9692 30490
rect 9396 30436 9452 30438
rect 9476 30436 9532 30438
rect 9556 30436 9612 30438
rect 9636 30436 9692 30438
rect 938 29996 940 30016
rect 940 29996 992 30016
rect 992 29996 994 30016
rect 938 29960 994 29996
rect 5176 29946 5232 29948
rect 5256 29946 5312 29948
rect 5336 29946 5392 29948
rect 5416 29946 5472 29948
rect 5176 29894 5222 29946
rect 5222 29894 5232 29946
rect 5256 29894 5286 29946
rect 5286 29894 5298 29946
rect 5298 29894 5312 29946
rect 5336 29894 5350 29946
rect 5350 29894 5362 29946
rect 5362 29894 5392 29946
rect 5416 29894 5426 29946
rect 5426 29894 5472 29946
rect 5176 29892 5232 29894
rect 5256 29892 5312 29894
rect 5336 29892 5392 29894
rect 5416 29892 5472 29894
rect 13617 29946 13673 29948
rect 13697 29946 13753 29948
rect 13777 29946 13833 29948
rect 13857 29946 13913 29948
rect 13617 29894 13663 29946
rect 13663 29894 13673 29946
rect 13697 29894 13727 29946
rect 13727 29894 13739 29946
rect 13739 29894 13753 29946
rect 13777 29894 13791 29946
rect 13791 29894 13803 29946
rect 13803 29894 13833 29946
rect 13857 29894 13867 29946
rect 13867 29894 13913 29946
rect 13617 29892 13673 29894
rect 13697 29892 13753 29894
rect 13777 29892 13833 29894
rect 13857 29892 13913 29894
rect 9396 29402 9452 29404
rect 9476 29402 9532 29404
rect 9556 29402 9612 29404
rect 9636 29402 9692 29404
rect 9396 29350 9442 29402
rect 9442 29350 9452 29402
rect 9476 29350 9506 29402
rect 9506 29350 9518 29402
rect 9518 29350 9532 29402
rect 9556 29350 9570 29402
rect 9570 29350 9582 29402
rect 9582 29350 9612 29402
rect 9636 29350 9646 29402
rect 9646 29350 9692 29402
rect 9396 29348 9452 29350
rect 9476 29348 9532 29350
rect 9556 29348 9612 29350
rect 9636 29348 9692 29350
rect 5176 28858 5232 28860
rect 5256 28858 5312 28860
rect 5336 28858 5392 28860
rect 5416 28858 5472 28860
rect 5176 28806 5222 28858
rect 5222 28806 5232 28858
rect 5256 28806 5286 28858
rect 5286 28806 5298 28858
rect 5298 28806 5312 28858
rect 5336 28806 5350 28858
rect 5350 28806 5362 28858
rect 5362 28806 5392 28858
rect 5416 28806 5426 28858
rect 5426 28806 5472 28858
rect 5176 28804 5232 28806
rect 5256 28804 5312 28806
rect 5336 28804 5392 28806
rect 5416 28804 5472 28806
rect 13617 28858 13673 28860
rect 13697 28858 13753 28860
rect 13777 28858 13833 28860
rect 13857 28858 13913 28860
rect 13617 28806 13663 28858
rect 13663 28806 13673 28858
rect 13697 28806 13727 28858
rect 13727 28806 13739 28858
rect 13739 28806 13753 28858
rect 13777 28806 13791 28858
rect 13791 28806 13803 28858
rect 13803 28806 13833 28858
rect 13857 28806 13867 28858
rect 13867 28806 13913 28858
rect 13617 28804 13673 28806
rect 13697 28804 13753 28806
rect 13777 28804 13833 28806
rect 13857 28804 13913 28806
rect 9396 28314 9452 28316
rect 9476 28314 9532 28316
rect 9556 28314 9612 28316
rect 9636 28314 9692 28316
rect 9396 28262 9442 28314
rect 9442 28262 9452 28314
rect 9476 28262 9506 28314
rect 9506 28262 9518 28314
rect 9518 28262 9532 28314
rect 9556 28262 9570 28314
rect 9570 28262 9582 28314
rect 9582 28262 9612 28314
rect 9636 28262 9646 28314
rect 9646 28262 9692 28314
rect 9396 28260 9452 28262
rect 9476 28260 9532 28262
rect 9556 28260 9612 28262
rect 9636 28260 9692 28262
rect 5176 27770 5232 27772
rect 5256 27770 5312 27772
rect 5336 27770 5392 27772
rect 5416 27770 5472 27772
rect 5176 27718 5222 27770
rect 5222 27718 5232 27770
rect 5256 27718 5286 27770
rect 5286 27718 5298 27770
rect 5298 27718 5312 27770
rect 5336 27718 5350 27770
rect 5350 27718 5362 27770
rect 5362 27718 5392 27770
rect 5416 27718 5426 27770
rect 5426 27718 5472 27770
rect 5176 27716 5232 27718
rect 5256 27716 5312 27718
rect 5336 27716 5392 27718
rect 5416 27716 5472 27718
rect 13617 27770 13673 27772
rect 13697 27770 13753 27772
rect 13777 27770 13833 27772
rect 13857 27770 13913 27772
rect 13617 27718 13663 27770
rect 13663 27718 13673 27770
rect 13697 27718 13727 27770
rect 13727 27718 13739 27770
rect 13739 27718 13753 27770
rect 13777 27718 13791 27770
rect 13791 27718 13803 27770
rect 13803 27718 13833 27770
rect 13857 27718 13867 27770
rect 13867 27718 13913 27770
rect 13617 27716 13673 27718
rect 13697 27716 13753 27718
rect 13777 27716 13833 27718
rect 13857 27716 13913 27718
rect 9396 27226 9452 27228
rect 9476 27226 9532 27228
rect 9556 27226 9612 27228
rect 9636 27226 9692 27228
rect 9396 27174 9442 27226
rect 9442 27174 9452 27226
rect 9476 27174 9506 27226
rect 9506 27174 9518 27226
rect 9518 27174 9532 27226
rect 9556 27174 9570 27226
rect 9570 27174 9582 27226
rect 9582 27174 9612 27226
rect 9636 27174 9646 27226
rect 9646 27174 9692 27226
rect 9396 27172 9452 27174
rect 9476 27172 9532 27174
rect 9556 27172 9612 27174
rect 9636 27172 9692 27174
rect 5176 26682 5232 26684
rect 5256 26682 5312 26684
rect 5336 26682 5392 26684
rect 5416 26682 5472 26684
rect 5176 26630 5222 26682
rect 5222 26630 5232 26682
rect 5256 26630 5286 26682
rect 5286 26630 5298 26682
rect 5298 26630 5312 26682
rect 5336 26630 5350 26682
rect 5350 26630 5362 26682
rect 5362 26630 5392 26682
rect 5416 26630 5426 26682
rect 5426 26630 5472 26682
rect 5176 26628 5232 26630
rect 5256 26628 5312 26630
rect 5336 26628 5392 26630
rect 5416 26628 5472 26630
rect 13617 26682 13673 26684
rect 13697 26682 13753 26684
rect 13777 26682 13833 26684
rect 13857 26682 13913 26684
rect 13617 26630 13663 26682
rect 13663 26630 13673 26682
rect 13697 26630 13727 26682
rect 13727 26630 13739 26682
rect 13739 26630 13753 26682
rect 13777 26630 13791 26682
rect 13791 26630 13803 26682
rect 13803 26630 13833 26682
rect 13857 26630 13867 26682
rect 13867 26630 13913 26682
rect 13617 26628 13673 26630
rect 13697 26628 13753 26630
rect 13777 26628 13833 26630
rect 13857 26628 13913 26630
rect 9396 26138 9452 26140
rect 9476 26138 9532 26140
rect 9556 26138 9612 26140
rect 9636 26138 9692 26140
rect 9396 26086 9442 26138
rect 9442 26086 9452 26138
rect 9476 26086 9506 26138
rect 9506 26086 9518 26138
rect 9518 26086 9532 26138
rect 9556 26086 9570 26138
rect 9570 26086 9582 26138
rect 9582 26086 9612 26138
rect 9636 26086 9646 26138
rect 9646 26086 9692 26138
rect 9396 26084 9452 26086
rect 9476 26084 9532 26086
rect 9556 26084 9612 26086
rect 9636 26084 9692 26086
rect 5176 25594 5232 25596
rect 5256 25594 5312 25596
rect 5336 25594 5392 25596
rect 5416 25594 5472 25596
rect 5176 25542 5222 25594
rect 5222 25542 5232 25594
rect 5256 25542 5286 25594
rect 5286 25542 5298 25594
rect 5298 25542 5312 25594
rect 5336 25542 5350 25594
rect 5350 25542 5362 25594
rect 5362 25542 5392 25594
rect 5416 25542 5426 25594
rect 5426 25542 5472 25594
rect 5176 25540 5232 25542
rect 5256 25540 5312 25542
rect 5336 25540 5392 25542
rect 5416 25540 5472 25542
rect 13617 25594 13673 25596
rect 13697 25594 13753 25596
rect 13777 25594 13833 25596
rect 13857 25594 13913 25596
rect 13617 25542 13663 25594
rect 13663 25542 13673 25594
rect 13697 25542 13727 25594
rect 13727 25542 13739 25594
rect 13739 25542 13753 25594
rect 13777 25542 13791 25594
rect 13791 25542 13803 25594
rect 13803 25542 13833 25594
rect 13857 25542 13867 25594
rect 13867 25542 13913 25594
rect 13617 25540 13673 25542
rect 13697 25540 13753 25542
rect 13777 25540 13833 25542
rect 13857 25540 13913 25542
rect 9396 25050 9452 25052
rect 9476 25050 9532 25052
rect 9556 25050 9612 25052
rect 9636 25050 9692 25052
rect 9396 24998 9442 25050
rect 9442 24998 9452 25050
rect 9476 24998 9506 25050
rect 9506 24998 9518 25050
rect 9518 24998 9532 25050
rect 9556 24998 9570 25050
rect 9570 24998 9582 25050
rect 9582 24998 9612 25050
rect 9636 24998 9646 25050
rect 9646 24998 9692 25050
rect 9396 24996 9452 24998
rect 9476 24996 9532 24998
rect 9556 24996 9612 24998
rect 9636 24996 9692 24998
rect 5176 24506 5232 24508
rect 5256 24506 5312 24508
rect 5336 24506 5392 24508
rect 5416 24506 5472 24508
rect 5176 24454 5222 24506
rect 5222 24454 5232 24506
rect 5256 24454 5286 24506
rect 5286 24454 5298 24506
rect 5298 24454 5312 24506
rect 5336 24454 5350 24506
rect 5350 24454 5362 24506
rect 5362 24454 5392 24506
rect 5416 24454 5426 24506
rect 5426 24454 5472 24506
rect 5176 24452 5232 24454
rect 5256 24452 5312 24454
rect 5336 24452 5392 24454
rect 5416 24452 5472 24454
rect 13617 24506 13673 24508
rect 13697 24506 13753 24508
rect 13777 24506 13833 24508
rect 13857 24506 13913 24508
rect 13617 24454 13663 24506
rect 13663 24454 13673 24506
rect 13697 24454 13727 24506
rect 13727 24454 13739 24506
rect 13739 24454 13753 24506
rect 13777 24454 13791 24506
rect 13791 24454 13803 24506
rect 13803 24454 13833 24506
rect 13857 24454 13867 24506
rect 13867 24454 13913 24506
rect 13617 24452 13673 24454
rect 13697 24452 13753 24454
rect 13777 24452 13833 24454
rect 13857 24452 13913 24454
rect 9396 23962 9452 23964
rect 9476 23962 9532 23964
rect 9556 23962 9612 23964
rect 9636 23962 9692 23964
rect 9396 23910 9442 23962
rect 9442 23910 9452 23962
rect 9476 23910 9506 23962
rect 9506 23910 9518 23962
rect 9518 23910 9532 23962
rect 9556 23910 9570 23962
rect 9570 23910 9582 23962
rect 9582 23910 9612 23962
rect 9636 23910 9646 23962
rect 9646 23910 9692 23962
rect 9396 23908 9452 23910
rect 9476 23908 9532 23910
rect 9556 23908 9612 23910
rect 9636 23908 9692 23910
rect 5176 23418 5232 23420
rect 5256 23418 5312 23420
rect 5336 23418 5392 23420
rect 5416 23418 5472 23420
rect 5176 23366 5222 23418
rect 5222 23366 5232 23418
rect 5256 23366 5286 23418
rect 5286 23366 5298 23418
rect 5298 23366 5312 23418
rect 5336 23366 5350 23418
rect 5350 23366 5362 23418
rect 5362 23366 5392 23418
rect 5416 23366 5426 23418
rect 5426 23366 5472 23418
rect 5176 23364 5232 23366
rect 5256 23364 5312 23366
rect 5336 23364 5392 23366
rect 5416 23364 5472 23366
rect 13617 23418 13673 23420
rect 13697 23418 13753 23420
rect 13777 23418 13833 23420
rect 13857 23418 13913 23420
rect 13617 23366 13663 23418
rect 13663 23366 13673 23418
rect 13697 23366 13727 23418
rect 13727 23366 13739 23418
rect 13739 23366 13753 23418
rect 13777 23366 13791 23418
rect 13791 23366 13803 23418
rect 13803 23366 13833 23418
rect 13857 23366 13867 23418
rect 13867 23366 13913 23418
rect 13617 23364 13673 23366
rect 13697 23364 13753 23366
rect 13777 23364 13833 23366
rect 13857 23364 13913 23366
rect 9396 22874 9452 22876
rect 9476 22874 9532 22876
rect 9556 22874 9612 22876
rect 9636 22874 9692 22876
rect 9396 22822 9442 22874
rect 9442 22822 9452 22874
rect 9476 22822 9506 22874
rect 9506 22822 9518 22874
rect 9518 22822 9532 22874
rect 9556 22822 9570 22874
rect 9570 22822 9582 22874
rect 9582 22822 9612 22874
rect 9636 22822 9646 22874
rect 9646 22822 9692 22874
rect 9396 22820 9452 22822
rect 9476 22820 9532 22822
rect 9556 22820 9612 22822
rect 9636 22820 9692 22822
rect 5176 22330 5232 22332
rect 5256 22330 5312 22332
rect 5336 22330 5392 22332
rect 5416 22330 5472 22332
rect 5176 22278 5222 22330
rect 5222 22278 5232 22330
rect 5256 22278 5286 22330
rect 5286 22278 5298 22330
rect 5298 22278 5312 22330
rect 5336 22278 5350 22330
rect 5350 22278 5362 22330
rect 5362 22278 5392 22330
rect 5416 22278 5426 22330
rect 5426 22278 5472 22330
rect 5176 22276 5232 22278
rect 5256 22276 5312 22278
rect 5336 22276 5392 22278
rect 5416 22276 5472 22278
rect 13617 22330 13673 22332
rect 13697 22330 13753 22332
rect 13777 22330 13833 22332
rect 13857 22330 13913 22332
rect 13617 22278 13663 22330
rect 13663 22278 13673 22330
rect 13697 22278 13727 22330
rect 13727 22278 13739 22330
rect 13739 22278 13753 22330
rect 13777 22278 13791 22330
rect 13791 22278 13803 22330
rect 13803 22278 13833 22330
rect 13857 22278 13867 22330
rect 13867 22278 13913 22330
rect 13617 22276 13673 22278
rect 13697 22276 13753 22278
rect 13777 22276 13833 22278
rect 13857 22276 13913 22278
rect 17837 39194 17893 39196
rect 17917 39194 17973 39196
rect 17997 39194 18053 39196
rect 18077 39194 18133 39196
rect 17837 39142 17883 39194
rect 17883 39142 17893 39194
rect 17917 39142 17947 39194
rect 17947 39142 17959 39194
rect 17959 39142 17973 39194
rect 17997 39142 18011 39194
rect 18011 39142 18023 39194
rect 18023 39142 18053 39194
rect 18077 39142 18087 39194
rect 18087 39142 18133 39194
rect 17837 39140 17893 39142
rect 17917 39140 17973 39142
rect 17997 39140 18053 39142
rect 18077 39140 18133 39142
rect 26278 39194 26334 39196
rect 26358 39194 26414 39196
rect 26438 39194 26494 39196
rect 26518 39194 26574 39196
rect 26278 39142 26324 39194
rect 26324 39142 26334 39194
rect 26358 39142 26388 39194
rect 26388 39142 26400 39194
rect 26400 39142 26414 39194
rect 26438 39142 26452 39194
rect 26452 39142 26464 39194
rect 26464 39142 26494 39194
rect 26518 39142 26528 39194
rect 26528 39142 26574 39194
rect 26278 39140 26334 39142
rect 26358 39140 26414 39142
rect 26438 39140 26494 39142
rect 26518 39140 26574 39142
rect 22058 38650 22114 38652
rect 22138 38650 22194 38652
rect 22218 38650 22274 38652
rect 22298 38650 22354 38652
rect 22058 38598 22104 38650
rect 22104 38598 22114 38650
rect 22138 38598 22168 38650
rect 22168 38598 22180 38650
rect 22180 38598 22194 38650
rect 22218 38598 22232 38650
rect 22232 38598 22244 38650
rect 22244 38598 22274 38650
rect 22298 38598 22308 38650
rect 22308 38598 22354 38650
rect 22058 38596 22114 38598
rect 22138 38596 22194 38598
rect 22218 38596 22274 38598
rect 22298 38596 22354 38598
rect 30499 38650 30555 38652
rect 30579 38650 30635 38652
rect 30659 38650 30715 38652
rect 30739 38650 30795 38652
rect 30499 38598 30545 38650
rect 30545 38598 30555 38650
rect 30579 38598 30609 38650
rect 30609 38598 30621 38650
rect 30621 38598 30635 38650
rect 30659 38598 30673 38650
rect 30673 38598 30685 38650
rect 30685 38598 30715 38650
rect 30739 38598 30749 38650
rect 30749 38598 30795 38650
rect 30499 38596 30555 38598
rect 30579 38596 30635 38598
rect 30659 38596 30715 38598
rect 30739 38596 30795 38598
rect 17837 38106 17893 38108
rect 17917 38106 17973 38108
rect 17997 38106 18053 38108
rect 18077 38106 18133 38108
rect 17837 38054 17883 38106
rect 17883 38054 17893 38106
rect 17917 38054 17947 38106
rect 17947 38054 17959 38106
rect 17959 38054 17973 38106
rect 17997 38054 18011 38106
rect 18011 38054 18023 38106
rect 18023 38054 18053 38106
rect 18077 38054 18087 38106
rect 18087 38054 18133 38106
rect 17837 38052 17893 38054
rect 17917 38052 17973 38054
rect 17997 38052 18053 38054
rect 18077 38052 18133 38054
rect 26278 38106 26334 38108
rect 26358 38106 26414 38108
rect 26438 38106 26494 38108
rect 26518 38106 26574 38108
rect 26278 38054 26324 38106
rect 26324 38054 26334 38106
rect 26358 38054 26388 38106
rect 26388 38054 26400 38106
rect 26400 38054 26414 38106
rect 26438 38054 26452 38106
rect 26452 38054 26464 38106
rect 26464 38054 26494 38106
rect 26518 38054 26528 38106
rect 26528 38054 26574 38106
rect 26278 38052 26334 38054
rect 26358 38052 26414 38054
rect 26438 38052 26494 38054
rect 26518 38052 26574 38054
rect 22058 37562 22114 37564
rect 22138 37562 22194 37564
rect 22218 37562 22274 37564
rect 22298 37562 22354 37564
rect 22058 37510 22104 37562
rect 22104 37510 22114 37562
rect 22138 37510 22168 37562
rect 22168 37510 22180 37562
rect 22180 37510 22194 37562
rect 22218 37510 22232 37562
rect 22232 37510 22244 37562
rect 22244 37510 22274 37562
rect 22298 37510 22308 37562
rect 22308 37510 22354 37562
rect 22058 37508 22114 37510
rect 22138 37508 22194 37510
rect 22218 37508 22274 37510
rect 22298 37508 22354 37510
rect 30499 37562 30555 37564
rect 30579 37562 30635 37564
rect 30659 37562 30715 37564
rect 30739 37562 30795 37564
rect 30499 37510 30545 37562
rect 30545 37510 30555 37562
rect 30579 37510 30609 37562
rect 30609 37510 30621 37562
rect 30621 37510 30635 37562
rect 30659 37510 30673 37562
rect 30673 37510 30685 37562
rect 30685 37510 30715 37562
rect 30739 37510 30749 37562
rect 30749 37510 30795 37562
rect 30499 37508 30555 37510
rect 30579 37508 30635 37510
rect 30659 37508 30715 37510
rect 30739 37508 30795 37510
rect 17837 37018 17893 37020
rect 17917 37018 17973 37020
rect 17997 37018 18053 37020
rect 18077 37018 18133 37020
rect 17837 36966 17883 37018
rect 17883 36966 17893 37018
rect 17917 36966 17947 37018
rect 17947 36966 17959 37018
rect 17959 36966 17973 37018
rect 17997 36966 18011 37018
rect 18011 36966 18023 37018
rect 18023 36966 18053 37018
rect 18077 36966 18087 37018
rect 18087 36966 18133 37018
rect 17837 36964 17893 36966
rect 17917 36964 17973 36966
rect 17997 36964 18053 36966
rect 18077 36964 18133 36966
rect 26278 37018 26334 37020
rect 26358 37018 26414 37020
rect 26438 37018 26494 37020
rect 26518 37018 26574 37020
rect 26278 36966 26324 37018
rect 26324 36966 26334 37018
rect 26358 36966 26388 37018
rect 26388 36966 26400 37018
rect 26400 36966 26414 37018
rect 26438 36966 26452 37018
rect 26452 36966 26464 37018
rect 26464 36966 26494 37018
rect 26518 36966 26528 37018
rect 26528 36966 26574 37018
rect 26278 36964 26334 36966
rect 26358 36964 26414 36966
rect 26438 36964 26494 36966
rect 26518 36964 26574 36966
rect 22058 36474 22114 36476
rect 22138 36474 22194 36476
rect 22218 36474 22274 36476
rect 22298 36474 22354 36476
rect 22058 36422 22104 36474
rect 22104 36422 22114 36474
rect 22138 36422 22168 36474
rect 22168 36422 22180 36474
rect 22180 36422 22194 36474
rect 22218 36422 22232 36474
rect 22232 36422 22244 36474
rect 22244 36422 22274 36474
rect 22298 36422 22308 36474
rect 22308 36422 22354 36474
rect 22058 36420 22114 36422
rect 22138 36420 22194 36422
rect 22218 36420 22274 36422
rect 22298 36420 22354 36422
rect 30499 36474 30555 36476
rect 30579 36474 30635 36476
rect 30659 36474 30715 36476
rect 30739 36474 30795 36476
rect 30499 36422 30545 36474
rect 30545 36422 30555 36474
rect 30579 36422 30609 36474
rect 30609 36422 30621 36474
rect 30621 36422 30635 36474
rect 30659 36422 30673 36474
rect 30673 36422 30685 36474
rect 30685 36422 30715 36474
rect 30739 36422 30749 36474
rect 30749 36422 30795 36474
rect 30499 36420 30555 36422
rect 30579 36420 30635 36422
rect 30659 36420 30715 36422
rect 30739 36420 30795 36422
rect 17837 35930 17893 35932
rect 17917 35930 17973 35932
rect 17997 35930 18053 35932
rect 18077 35930 18133 35932
rect 17837 35878 17883 35930
rect 17883 35878 17893 35930
rect 17917 35878 17947 35930
rect 17947 35878 17959 35930
rect 17959 35878 17973 35930
rect 17997 35878 18011 35930
rect 18011 35878 18023 35930
rect 18023 35878 18053 35930
rect 18077 35878 18087 35930
rect 18087 35878 18133 35930
rect 17837 35876 17893 35878
rect 17917 35876 17973 35878
rect 17997 35876 18053 35878
rect 18077 35876 18133 35878
rect 26278 35930 26334 35932
rect 26358 35930 26414 35932
rect 26438 35930 26494 35932
rect 26518 35930 26574 35932
rect 26278 35878 26324 35930
rect 26324 35878 26334 35930
rect 26358 35878 26388 35930
rect 26388 35878 26400 35930
rect 26400 35878 26414 35930
rect 26438 35878 26452 35930
rect 26452 35878 26464 35930
rect 26464 35878 26494 35930
rect 26518 35878 26528 35930
rect 26528 35878 26574 35930
rect 26278 35876 26334 35878
rect 26358 35876 26414 35878
rect 26438 35876 26494 35878
rect 26518 35876 26574 35878
rect 22058 35386 22114 35388
rect 22138 35386 22194 35388
rect 22218 35386 22274 35388
rect 22298 35386 22354 35388
rect 22058 35334 22104 35386
rect 22104 35334 22114 35386
rect 22138 35334 22168 35386
rect 22168 35334 22180 35386
rect 22180 35334 22194 35386
rect 22218 35334 22232 35386
rect 22232 35334 22244 35386
rect 22244 35334 22274 35386
rect 22298 35334 22308 35386
rect 22308 35334 22354 35386
rect 22058 35332 22114 35334
rect 22138 35332 22194 35334
rect 22218 35332 22274 35334
rect 22298 35332 22354 35334
rect 30499 35386 30555 35388
rect 30579 35386 30635 35388
rect 30659 35386 30715 35388
rect 30739 35386 30795 35388
rect 30499 35334 30545 35386
rect 30545 35334 30555 35386
rect 30579 35334 30609 35386
rect 30609 35334 30621 35386
rect 30621 35334 30635 35386
rect 30659 35334 30673 35386
rect 30673 35334 30685 35386
rect 30685 35334 30715 35386
rect 30739 35334 30749 35386
rect 30749 35334 30795 35386
rect 30499 35332 30555 35334
rect 30579 35332 30635 35334
rect 30659 35332 30715 35334
rect 30739 35332 30795 35334
rect 17837 34842 17893 34844
rect 17917 34842 17973 34844
rect 17997 34842 18053 34844
rect 18077 34842 18133 34844
rect 17837 34790 17883 34842
rect 17883 34790 17893 34842
rect 17917 34790 17947 34842
rect 17947 34790 17959 34842
rect 17959 34790 17973 34842
rect 17997 34790 18011 34842
rect 18011 34790 18023 34842
rect 18023 34790 18053 34842
rect 18077 34790 18087 34842
rect 18087 34790 18133 34842
rect 17837 34788 17893 34790
rect 17917 34788 17973 34790
rect 17997 34788 18053 34790
rect 18077 34788 18133 34790
rect 26278 34842 26334 34844
rect 26358 34842 26414 34844
rect 26438 34842 26494 34844
rect 26518 34842 26574 34844
rect 26278 34790 26324 34842
rect 26324 34790 26334 34842
rect 26358 34790 26388 34842
rect 26388 34790 26400 34842
rect 26400 34790 26414 34842
rect 26438 34790 26452 34842
rect 26452 34790 26464 34842
rect 26464 34790 26494 34842
rect 26518 34790 26528 34842
rect 26528 34790 26574 34842
rect 26278 34788 26334 34790
rect 26358 34788 26414 34790
rect 26438 34788 26494 34790
rect 26518 34788 26574 34790
rect 22058 34298 22114 34300
rect 22138 34298 22194 34300
rect 22218 34298 22274 34300
rect 22298 34298 22354 34300
rect 22058 34246 22104 34298
rect 22104 34246 22114 34298
rect 22138 34246 22168 34298
rect 22168 34246 22180 34298
rect 22180 34246 22194 34298
rect 22218 34246 22232 34298
rect 22232 34246 22244 34298
rect 22244 34246 22274 34298
rect 22298 34246 22308 34298
rect 22308 34246 22354 34298
rect 22058 34244 22114 34246
rect 22138 34244 22194 34246
rect 22218 34244 22274 34246
rect 22298 34244 22354 34246
rect 30499 34298 30555 34300
rect 30579 34298 30635 34300
rect 30659 34298 30715 34300
rect 30739 34298 30795 34300
rect 30499 34246 30545 34298
rect 30545 34246 30555 34298
rect 30579 34246 30609 34298
rect 30609 34246 30621 34298
rect 30621 34246 30635 34298
rect 30659 34246 30673 34298
rect 30673 34246 30685 34298
rect 30685 34246 30715 34298
rect 30739 34246 30749 34298
rect 30749 34246 30795 34298
rect 30499 34244 30555 34246
rect 30579 34244 30635 34246
rect 30659 34244 30715 34246
rect 30739 34244 30795 34246
rect 17837 33754 17893 33756
rect 17917 33754 17973 33756
rect 17997 33754 18053 33756
rect 18077 33754 18133 33756
rect 17837 33702 17883 33754
rect 17883 33702 17893 33754
rect 17917 33702 17947 33754
rect 17947 33702 17959 33754
rect 17959 33702 17973 33754
rect 17997 33702 18011 33754
rect 18011 33702 18023 33754
rect 18023 33702 18053 33754
rect 18077 33702 18087 33754
rect 18087 33702 18133 33754
rect 17837 33700 17893 33702
rect 17917 33700 17973 33702
rect 17997 33700 18053 33702
rect 18077 33700 18133 33702
rect 22058 33210 22114 33212
rect 22138 33210 22194 33212
rect 22218 33210 22274 33212
rect 22298 33210 22354 33212
rect 22058 33158 22104 33210
rect 22104 33158 22114 33210
rect 22138 33158 22168 33210
rect 22168 33158 22180 33210
rect 22180 33158 22194 33210
rect 22218 33158 22232 33210
rect 22232 33158 22244 33210
rect 22244 33158 22274 33210
rect 22298 33158 22308 33210
rect 22308 33158 22354 33210
rect 22058 33156 22114 33158
rect 22138 33156 22194 33158
rect 22218 33156 22274 33158
rect 22298 33156 22354 33158
rect 17837 32666 17893 32668
rect 17917 32666 17973 32668
rect 17997 32666 18053 32668
rect 18077 32666 18133 32668
rect 17837 32614 17883 32666
rect 17883 32614 17893 32666
rect 17917 32614 17947 32666
rect 17947 32614 17959 32666
rect 17959 32614 17973 32666
rect 17997 32614 18011 32666
rect 18011 32614 18023 32666
rect 18023 32614 18053 32666
rect 18077 32614 18087 32666
rect 18087 32614 18133 32666
rect 17837 32612 17893 32614
rect 17917 32612 17973 32614
rect 17997 32612 18053 32614
rect 18077 32612 18133 32614
rect 17837 31578 17893 31580
rect 17917 31578 17973 31580
rect 17997 31578 18053 31580
rect 18077 31578 18133 31580
rect 17837 31526 17883 31578
rect 17883 31526 17893 31578
rect 17917 31526 17947 31578
rect 17947 31526 17959 31578
rect 17959 31526 17973 31578
rect 17997 31526 18011 31578
rect 18011 31526 18023 31578
rect 18023 31526 18053 31578
rect 18077 31526 18087 31578
rect 18087 31526 18133 31578
rect 17837 31524 17893 31526
rect 17917 31524 17973 31526
rect 17997 31524 18053 31526
rect 18077 31524 18133 31526
rect 17837 30490 17893 30492
rect 17917 30490 17973 30492
rect 17997 30490 18053 30492
rect 18077 30490 18133 30492
rect 17837 30438 17883 30490
rect 17883 30438 17893 30490
rect 17917 30438 17947 30490
rect 17947 30438 17959 30490
rect 17959 30438 17973 30490
rect 17997 30438 18011 30490
rect 18011 30438 18023 30490
rect 18023 30438 18053 30490
rect 18077 30438 18087 30490
rect 18087 30438 18133 30490
rect 17837 30436 17893 30438
rect 17917 30436 17973 30438
rect 17997 30436 18053 30438
rect 18077 30436 18133 30438
rect 17837 29402 17893 29404
rect 17917 29402 17973 29404
rect 17997 29402 18053 29404
rect 18077 29402 18133 29404
rect 17837 29350 17883 29402
rect 17883 29350 17893 29402
rect 17917 29350 17947 29402
rect 17947 29350 17959 29402
rect 17959 29350 17973 29402
rect 17997 29350 18011 29402
rect 18011 29350 18023 29402
rect 18023 29350 18053 29402
rect 18077 29350 18087 29402
rect 18087 29350 18133 29402
rect 17837 29348 17893 29350
rect 17917 29348 17973 29350
rect 17997 29348 18053 29350
rect 18077 29348 18133 29350
rect 18694 30676 18696 30696
rect 18696 30676 18748 30696
rect 18748 30676 18750 30696
rect 18694 30640 18750 30676
rect 19246 30640 19302 30696
rect 17837 28314 17893 28316
rect 17917 28314 17973 28316
rect 17997 28314 18053 28316
rect 18077 28314 18133 28316
rect 17837 28262 17883 28314
rect 17883 28262 17893 28314
rect 17917 28262 17947 28314
rect 17947 28262 17959 28314
rect 17959 28262 17973 28314
rect 17997 28262 18011 28314
rect 18011 28262 18023 28314
rect 18023 28262 18053 28314
rect 18077 28262 18087 28314
rect 18087 28262 18133 28314
rect 17837 28260 17893 28262
rect 17917 28260 17973 28262
rect 17997 28260 18053 28262
rect 18077 28260 18133 28262
rect 17837 27226 17893 27228
rect 17917 27226 17973 27228
rect 17997 27226 18053 27228
rect 18077 27226 18133 27228
rect 17837 27174 17883 27226
rect 17883 27174 17893 27226
rect 17917 27174 17947 27226
rect 17947 27174 17959 27226
rect 17959 27174 17973 27226
rect 17997 27174 18011 27226
rect 18011 27174 18023 27226
rect 18023 27174 18053 27226
rect 18077 27174 18087 27226
rect 18087 27174 18133 27226
rect 17837 27172 17893 27174
rect 17917 27172 17973 27174
rect 17997 27172 18053 27174
rect 18077 27172 18133 27174
rect 17837 26138 17893 26140
rect 17917 26138 17973 26140
rect 17997 26138 18053 26140
rect 18077 26138 18133 26140
rect 17837 26086 17883 26138
rect 17883 26086 17893 26138
rect 17917 26086 17947 26138
rect 17947 26086 17959 26138
rect 17959 26086 17973 26138
rect 17997 26086 18011 26138
rect 18011 26086 18023 26138
rect 18023 26086 18053 26138
rect 18077 26086 18087 26138
rect 18087 26086 18133 26138
rect 17837 26084 17893 26086
rect 17917 26084 17973 26086
rect 17997 26084 18053 26086
rect 18077 26084 18133 26086
rect 22058 32122 22114 32124
rect 22138 32122 22194 32124
rect 22218 32122 22274 32124
rect 22298 32122 22354 32124
rect 22058 32070 22104 32122
rect 22104 32070 22114 32122
rect 22138 32070 22168 32122
rect 22168 32070 22180 32122
rect 22180 32070 22194 32122
rect 22218 32070 22232 32122
rect 22232 32070 22244 32122
rect 22244 32070 22274 32122
rect 22298 32070 22308 32122
rect 22308 32070 22354 32122
rect 22058 32068 22114 32070
rect 22138 32068 22194 32070
rect 22218 32068 22274 32070
rect 22298 32068 22354 32070
rect 20350 29144 20406 29200
rect 20902 29144 20958 29200
rect 26278 33754 26334 33756
rect 26358 33754 26414 33756
rect 26438 33754 26494 33756
rect 26518 33754 26574 33756
rect 26278 33702 26324 33754
rect 26324 33702 26334 33754
rect 26358 33702 26388 33754
rect 26388 33702 26400 33754
rect 26400 33702 26414 33754
rect 26438 33702 26452 33754
rect 26452 33702 26464 33754
rect 26464 33702 26494 33754
rect 26518 33702 26528 33754
rect 26528 33702 26574 33754
rect 26278 33700 26334 33702
rect 26358 33700 26414 33702
rect 26438 33700 26494 33702
rect 26518 33700 26574 33702
rect 22058 31034 22114 31036
rect 22138 31034 22194 31036
rect 22218 31034 22274 31036
rect 22298 31034 22354 31036
rect 22058 30982 22104 31034
rect 22104 30982 22114 31034
rect 22138 30982 22168 31034
rect 22168 30982 22180 31034
rect 22180 30982 22194 31034
rect 22218 30982 22232 31034
rect 22232 30982 22244 31034
rect 22244 30982 22274 31034
rect 22298 30982 22308 31034
rect 22308 30982 22354 31034
rect 22058 30980 22114 30982
rect 22138 30980 22194 30982
rect 22218 30980 22274 30982
rect 22298 30980 22354 30982
rect 22058 29946 22114 29948
rect 22138 29946 22194 29948
rect 22218 29946 22274 29948
rect 22298 29946 22354 29948
rect 22058 29894 22104 29946
rect 22104 29894 22114 29946
rect 22138 29894 22168 29946
rect 22168 29894 22180 29946
rect 22180 29894 22194 29946
rect 22218 29894 22232 29946
rect 22232 29894 22244 29946
rect 22244 29894 22274 29946
rect 22298 29894 22308 29946
rect 22308 29894 22354 29946
rect 22058 29892 22114 29894
rect 22138 29892 22194 29894
rect 22218 29892 22274 29894
rect 22298 29892 22354 29894
rect 20442 27396 20498 27432
rect 20442 27376 20444 27396
rect 20444 27376 20496 27396
rect 20496 27376 20498 27396
rect 20074 26868 20076 26888
rect 20076 26868 20128 26888
rect 20128 26868 20130 26888
rect 17837 25050 17893 25052
rect 17917 25050 17973 25052
rect 17997 25050 18053 25052
rect 18077 25050 18133 25052
rect 17837 24998 17883 25050
rect 17883 24998 17893 25050
rect 17917 24998 17947 25050
rect 17947 24998 17959 25050
rect 17959 24998 17973 25050
rect 17997 24998 18011 25050
rect 18011 24998 18023 25050
rect 18023 24998 18053 25050
rect 18077 24998 18087 25050
rect 18087 24998 18133 25050
rect 17837 24996 17893 24998
rect 17917 24996 17973 24998
rect 17997 24996 18053 24998
rect 18077 24996 18133 24998
rect 20074 26832 20130 26868
rect 20810 27376 20866 27432
rect 22058 28858 22114 28860
rect 22138 28858 22194 28860
rect 22218 28858 22274 28860
rect 22298 28858 22354 28860
rect 22058 28806 22104 28858
rect 22104 28806 22114 28858
rect 22138 28806 22168 28858
rect 22168 28806 22180 28858
rect 22180 28806 22194 28858
rect 22218 28806 22232 28858
rect 22232 28806 22244 28858
rect 22244 28806 22274 28858
rect 22298 28806 22308 28858
rect 22308 28806 22354 28858
rect 22058 28804 22114 28806
rect 22138 28804 22194 28806
rect 22218 28804 22274 28806
rect 22298 28804 22354 28806
rect 22058 27770 22114 27772
rect 22138 27770 22194 27772
rect 22218 27770 22274 27772
rect 22298 27770 22354 27772
rect 22058 27718 22104 27770
rect 22104 27718 22114 27770
rect 22138 27718 22168 27770
rect 22168 27718 22180 27770
rect 22180 27718 22194 27770
rect 22218 27718 22232 27770
rect 22232 27718 22244 27770
rect 22244 27718 22274 27770
rect 22298 27718 22308 27770
rect 22308 27718 22354 27770
rect 22058 27716 22114 27718
rect 22138 27716 22194 27718
rect 22218 27716 22274 27718
rect 22298 27716 22354 27718
rect 20810 26968 20866 27024
rect 20902 26424 20958 26480
rect 17837 23962 17893 23964
rect 17917 23962 17973 23964
rect 17997 23962 18053 23964
rect 18077 23962 18133 23964
rect 17837 23910 17883 23962
rect 17883 23910 17893 23962
rect 17917 23910 17947 23962
rect 17947 23910 17959 23962
rect 17959 23910 17973 23962
rect 17997 23910 18011 23962
rect 18011 23910 18023 23962
rect 18023 23910 18053 23962
rect 18077 23910 18087 23962
rect 18087 23910 18133 23962
rect 17837 23908 17893 23910
rect 17917 23908 17973 23910
rect 17997 23908 18053 23910
rect 18077 23908 18133 23910
rect 17837 22874 17893 22876
rect 17917 22874 17973 22876
rect 17997 22874 18053 22876
rect 18077 22874 18133 22876
rect 17837 22822 17883 22874
rect 17883 22822 17893 22874
rect 17917 22822 17947 22874
rect 17947 22822 17959 22874
rect 17959 22822 17973 22874
rect 17997 22822 18011 22874
rect 18011 22822 18023 22874
rect 18023 22822 18053 22874
rect 18077 22822 18087 22874
rect 18087 22822 18133 22874
rect 17837 22820 17893 22822
rect 17917 22820 17973 22822
rect 17997 22820 18053 22822
rect 18077 22820 18133 22822
rect 9396 21786 9452 21788
rect 9476 21786 9532 21788
rect 9556 21786 9612 21788
rect 9636 21786 9692 21788
rect 9396 21734 9442 21786
rect 9442 21734 9452 21786
rect 9476 21734 9506 21786
rect 9506 21734 9518 21786
rect 9518 21734 9532 21786
rect 9556 21734 9570 21786
rect 9570 21734 9582 21786
rect 9582 21734 9612 21786
rect 9636 21734 9646 21786
rect 9646 21734 9692 21786
rect 9396 21732 9452 21734
rect 9476 21732 9532 21734
rect 9556 21732 9612 21734
rect 9636 21732 9692 21734
rect 5176 21242 5232 21244
rect 5256 21242 5312 21244
rect 5336 21242 5392 21244
rect 5416 21242 5472 21244
rect 5176 21190 5222 21242
rect 5222 21190 5232 21242
rect 5256 21190 5286 21242
rect 5286 21190 5298 21242
rect 5298 21190 5312 21242
rect 5336 21190 5350 21242
rect 5350 21190 5362 21242
rect 5362 21190 5392 21242
rect 5416 21190 5426 21242
rect 5426 21190 5472 21242
rect 5176 21188 5232 21190
rect 5256 21188 5312 21190
rect 5336 21188 5392 21190
rect 5416 21188 5472 21190
rect 13617 21242 13673 21244
rect 13697 21242 13753 21244
rect 13777 21242 13833 21244
rect 13857 21242 13913 21244
rect 13617 21190 13663 21242
rect 13663 21190 13673 21242
rect 13697 21190 13727 21242
rect 13727 21190 13739 21242
rect 13739 21190 13753 21242
rect 13777 21190 13791 21242
rect 13791 21190 13803 21242
rect 13803 21190 13833 21242
rect 13857 21190 13867 21242
rect 13867 21190 13913 21242
rect 13617 21188 13673 21190
rect 13697 21188 13753 21190
rect 13777 21188 13833 21190
rect 13857 21188 13913 21190
rect 9396 20698 9452 20700
rect 9476 20698 9532 20700
rect 9556 20698 9612 20700
rect 9636 20698 9692 20700
rect 9396 20646 9442 20698
rect 9442 20646 9452 20698
rect 9476 20646 9506 20698
rect 9506 20646 9518 20698
rect 9518 20646 9532 20698
rect 9556 20646 9570 20698
rect 9570 20646 9582 20698
rect 9582 20646 9612 20698
rect 9636 20646 9646 20698
rect 9646 20646 9692 20698
rect 9396 20644 9452 20646
rect 9476 20644 9532 20646
rect 9556 20644 9612 20646
rect 9636 20644 9692 20646
rect 5176 20154 5232 20156
rect 5256 20154 5312 20156
rect 5336 20154 5392 20156
rect 5416 20154 5472 20156
rect 5176 20102 5222 20154
rect 5222 20102 5232 20154
rect 5256 20102 5286 20154
rect 5286 20102 5298 20154
rect 5298 20102 5312 20154
rect 5336 20102 5350 20154
rect 5350 20102 5362 20154
rect 5362 20102 5392 20154
rect 5416 20102 5426 20154
rect 5426 20102 5472 20154
rect 5176 20100 5232 20102
rect 5256 20100 5312 20102
rect 5336 20100 5392 20102
rect 5416 20100 5472 20102
rect 13617 20154 13673 20156
rect 13697 20154 13753 20156
rect 13777 20154 13833 20156
rect 13857 20154 13913 20156
rect 13617 20102 13663 20154
rect 13663 20102 13673 20154
rect 13697 20102 13727 20154
rect 13727 20102 13739 20154
rect 13739 20102 13753 20154
rect 13777 20102 13791 20154
rect 13791 20102 13803 20154
rect 13803 20102 13833 20154
rect 13857 20102 13867 20154
rect 13867 20102 13913 20154
rect 13617 20100 13673 20102
rect 13697 20100 13753 20102
rect 13777 20100 13833 20102
rect 13857 20100 13913 20102
rect 938 19796 940 19816
rect 940 19796 992 19816
rect 992 19796 994 19816
rect 938 19760 994 19796
rect 9396 19610 9452 19612
rect 9476 19610 9532 19612
rect 9556 19610 9612 19612
rect 9636 19610 9692 19612
rect 9396 19558 9442 19610
rect 9442 19558 9452 19610
rect 9476 19558 9506 19610
rect 9506 19558 9518 19610
rect 9518 19558 9532 19610
rect 9556 19558 9570 19610
rect 9570 19558 9582 19610
rect 9582 19558 9612 19610
rect 9636 19558 9646 19610
rect 9646 19558 9692 19610
rect 9396 19556 9452 19558
rect 9476 19556 9532 19558
rect 9556 19556 9612 19558
rect 9636 19556 9692 19558
rect 5176 19066 5232 19068
rect 5256 19066 5312 19068
rect 5336 19066 5392 19068
rect 5416 19066 5472 19068
rect 5176 19014 5222 19066
rect 5222 19014 5232 19066
rect 5256 19014 5286 19066
rect 5286 19014 5298 19066
rect 5298 19014 5312 19066
rect 5336 19014 5350 19066
rect 5350 19014 5362 19066
rect 5362 19014 5392 19066
rect 5416 19014 5426 19066
rect 5426 19014 5472 19066
rect 5176 19012 5232 19014
rect 5256 19012 5312 19014
rect 5336 19012 5392 19014
rect 5416 19012 5472 19014
rect 13617 19066 13673 19068
rect 13697 19066 13753 19068
rect 13777 19066 13833 19068
rect 13857 19066 13913 19068
rect 13617 19014 13663 19066
rect 13663 19014 13673 19066
rect 13697 19014 13727 19066
rect 13727 19014 13739 19066
rect 13739 19014 13753 19066
rect 13777 19014 13791 19066
rect 13791 19014 13803 19066
rect 13803 19014 13833 19066
rect 13857 19014 13867 19066
rect 13867 19014 13913 19066
rect 13617 19012 13673 19014
rect 13697 19012 13753 19014
rect 13777 19012 13833 19014
rect 13857 19012 13913 19014
rect 9396 18522 9452 18524
rect 9476 18522 9532 18524
rect 9556 18522 9612 18524
rect 9636 18522 9692 18524
rect 9396 18470 9442 18522
rect 9442 18470 9452 18522
rect 9476 18470 9506 18522
rect 9506 18470 9518 18522
rect 9518 18470 9532 18522
rect 9556 18470 9570 18522
rect 9570 18470 9582 18522
rect 9582 18470 9612 18522
rect 9636 18470 9646 18522
rect 9646 18470 9692 18522
rect 9396 18468 9452 18470
rect 9476 18468 9532 18470
rect 9556 18468 9612 18470
rect 9636 18468 9692 18470
rect 5176 17978 5232 17980
rect 5256 17978 5312 17980
rect 5336 17978 5392 17980
rect 5416 17978 5472 17980
rect 5176 17926 5222 17978
rect 5222 17926 5232 17978
rect 5256 17926 5286 17978
rect 5286 17926 5298 17978
rect 5298 17926 5312 17978
rect 5336 17926 5350 17978
rect 5350 17926 5362 17978
rect 5362 17926 5392 17978
rect 5416 17926 5426 17978
rect 5426 17926 5472 17978
rect 5176 17924 5232 17926
rect 5256 17924 5312 17926
rect 5336 17924 5392 17926
rect 5416 17924 5472 17926
rect 13617 17978 13673 17980
rect 13697 17978 13753 17980
rect 13777 17978 13833 17980
rect 13857 17978 13913 17980
rect 13617 17926 13663 17978
rect 13663 17926 13673 17978
rect 13697 17926 13727 17978
rect 13727 17926 13739 17978
rect 13739 17926 13753 17978
rect 13777 17926 13791 17978
rect 13791 17926 13803 17978
rect 13803 17926 13833 17978
rect 13857 17926 13867 17978
rect 13867 17926 13913 17978
rect 13617 17924 13673 17926
rect 13697 17924 13753 17926
rect 13777 17924 13833 17926
rect 13857 17924 13913 17926
rect 9396 17434 9452 17436
rect 9476 17434 9532 17436
rect 9556 17434 9612 17436
rect 9636 17434 9692 17436
rect 9396 17382 9442 17434
rect 9442 17382 9452 17434
rect 9476 17382 9506 17434
rect 9506 17382 9518 17434
rect 9518 17382 9532 17434
rect 9556 17382 9570 17434
rect 9570 17382 9582 17434
rect 9582 17382 9612 17434
rect 9636 17382 9646 17434
rect 9646 17382 9692 17434
rect 9396 17380 9452 17382
rect 9476 17380 9532 17382
rect 9556 17380 9612 17382
rect 9636 17380 9692 17382
rect 17837 21786 17893 21788
rect 17917 21786 17973 21788
rect 17997 21786 18053 21788
rect 18077 21786 18133 21788
rect 17837 21734 17883 21786
rect 17883 21734 17893 21786
rect 17917 21734 17947 21786
rect 17947 21734 17959 21786
rect 17959 21734 17973 21786
rect 17997 21734 18011 21786
rect 18011 21734 18023 21786
rect 18023 21734 18053 21786
rect 18077 21734 18087 21786
rect 18087 21734 18133 21786
rect 17837 21732 17893 21734
rect 17917 21732 17973 21734
rect 17997 21732 18053 21734
rect 18077 21732 18133 21734
rect 17837 20698 17893 20700
rect 17917 20698 17973 20700
rect 17997 20698 18053 20700
rect 18077 20698 18133 20700
rect 17837 20646 17883 20698
rect 17883 20646 17893 20698
rect 17917 20646 17947 20698
rect 17947 20646 17959 20698
rect 17959 20646 17973 20698
rect 17997 20646 18011 20698
rect 18011 20646 18023 20698
rect 18023 20646 18053 20698
rect 18077 20646 18087 20698
rect 18087 20646 18133 20698
rect 17837 20644 17893 20646
rect 17917 20644 17973 20646
rect 17997 20644 18053 20646
rect 18077 20644 18133 20646
rect 17837 19610 17893 19612
rect 17917 19610 17973 19612
rect 17997 19610 18053 19612
rect 18077 19610 18133 19612
rect 17837 19558 17883 19610
rect 17883 19558 17893 19610
rect 17917 19558 17947 19610
rect 17947 19558 17959 19610
rect 17959 19558 17973 19610
rect 17997 19558 18011 19610
rect 18011 19558 18023 19610
rect 18023 19558 18053 19610
rect 18077 19558 18087 19610
rect 18087 19558 18133 19610
rect 17837 19556 17893 19558
rect 17917 19556 17973 19558
rect 17997 19556 18053 19558
rect 18077 19556 18133 19558
rect 17837 18522 17893 18524
rect 17917 18522 17973 18524
rect 17997 18522 18053 18524
rect 18077 18522 18133 18524
rect 17837 18470 17883 18522
rect 17883 18470 17893 18522
rect 17917 18470 17947 18522
rect 17947 18470 17959 18522
rect 17959 18470 17973 18522
rect 17997 18470 18011 18522
rect 18011 18470 18023 18522
rect 18023 18470 18053 18522
rect 18077 18470 18087 18522
rect 18087 18470 18133 18522
rect 17837 18468 17893 18470
rect 17917 18468 17973 18470
rect 17997 18468 18053 18470
rect 18077 18468 18133 18470
rect 20626 26288 20682 26344
rect 21270 26968 21326 27024
rect 21362 26832 21418 26888
rect 21362 26324 21364 26344
rect 21364 26324 21416 26344
rect 21416 26324 21418 26344
rect 21362 26288 21418 26324
rect 22058 26682 22114 26684
rect 22138 26682 22194 26684
rect 22218 26682 22274 26684
rect 22298 26682 22354 26684
rect 22058 26630 22104 26682
rect 22104 26630 22114 26682
rect 22138 26630 22168 26682
rect 22168 26630 22180 26682
rect 22180 26630 22194 26682
rect 22218 26630 22232 26682
rect 22232 26630 22244 26682
rect 22244 26630 22274 26682
rect 22298 26630 22308 26682
rect 22308 26630 22354 26682
rect 22058 26628 22114 26630
rect 22138 26628 22194 26630
rect 22218 26628 22274 26630
rect 22298 26628 22354 26630
rect 21914 26460 21916 26480
rect 21916 26460 21968 26480
rect 21968 26460 21970 26480
rect 21914 26424 21970 26460
rect 22058 25594 22114 25596
rect 22138 25594 22194 25596
rect 22218 25594 22274 25596
rect 22298 25594 22354 25596
rect 22058 25542 22104 25594
rect 22104 25542 22114 25594
rect 22138 25542 22168 25594
rect 22168 25542 22180 25594
rect 22180 25542 22194 25594
rect 22218 25542 22232 25594
rect 22232 25542 22244 25594
rect 22244 25542 22274 25594
rect 22298 25542 22308 25594
rect 22308 25542 22354 25594
rect 22058 25540 22114 25542
rect 22138 25540 22194 25542
rect 22218 25540 22274 25542
rect 22298 25540 22354 25542
rect 22058 24506 22114 24508
rect 22138 24506 22194 24508
rect 22218 24506 22274 24508
rect 22298 24506 22354 24508
rect 22058 24454 22104 24506
rect 22104 24454 22114 24506
rect 22138 24454 22168 24506
rect 22168 24454 22180 24506
rect 22180 24454 22194 24506
rect 22218 24454 22232 24506
rect 22232 24454 22244 24506
rect 22244 24454 22274 24506
rect 22298 24454 22308 24506
rect 22308 24454 22354 24506
rect 22058 24452 22114 24454
rect 22138 24452 22194 24454
rect 22218 24452 22274 24454
rect 22298 24452 22354 24454
rect 22058 23418 22114 23420
rect 22138 23418 22194 23420
rect 22218 23418 22274 23420
rect 22298 23418 22354 23420
rect 22058 23366 22104 23418
rect 22104 23366 22114 23418
rect 22138 23366 22168 23418
rect 22168 23366 22180 23418
rect 22180 23366 22194 23418
rect 22218 23366 22232 23418
rect 22232 23366 22244 23418
rect 22244 23366 22274 23418
rect 22298 23366 22308 23418
rect 22308 23366 22354 23418
rect 22058 23364 22114 23366
rect 22138 23364 22194 23366
rect 22218 23364 22274 23366
rect 22298 23364 22354 23366
rect 26278 32666 26334 32668
rect 26358 32666 26414 32668
rect 26438 32666 26494 32668
rect 26518 32666 26574 32668
rect 26278 32614 26324 32666
rect 26324 32614 26334 32666
rect 26358 32614 26388 32666
rect 26388 32614 26400 32666
rect 26400 32614 26414 32666
rect 26438 32614 26452 32666
rect 26452 32614 26464 32666
rect 26464 32614 26494 32666
rect 26518 32614 26528 32666
rect 26528 32614 26574 32666
rect 26278 32612 26334 32614
rect 26358 32612 26414 32614
rect 26438 32612 26494 32614
rect 26518 32612 26574 32614
rect 26278 31578 26334 31580
rect 26358 31578 26414 31580
rect 26438 31578 26494 31580
rect 26518 31578 26574 31580
rect 26278 31526 26324 31578
rect 26324 31526 26334 31578
rect 26358 31526 26388 31578
rect 26388 31526 26400 31578
rect 26400 31526 26414 31578
rect 26438 31526 26452 31578
rect 26452 31526 26464 31578
rect 26464 31526 26494 31578
rect 26518 31526 26528 31578
rect 26528 31526 26574 31578
rect 26278 31524 26334 31526
rect 26358 31524 26414 31526
rect 26438 31524 26494 31526
rect 26518 31524 26574 31526
rect 26278 30490 26334 30492
rect 26358 30490 26414 30492
rect 26438 30490 26494 30492
rect 26518 30490 26574 30492
rect 26278 30438 26324 30490
rect 26324 30438 26334 30490
rect 26358 30438 26388 30490
rect 26388 30438 26400 30490
rect 26400 30438 26414 30490
rect 26438 30438 26452 30490
rect 26452 30438 26464 30490
rect 26464 30438 26494 30490
rect 26518 30438 26528 30490
rect 26528 30438 26574 30490
rect 26278 30436 26334 30438
rect 26358 30436 26414 30438
rect 26438 30436 26494 30438
rect 26518 30436 26574 30438
rect 26278 29402 26334 29404
rect 26358 29402 26414 29404
rect 26438 29402 26494 29404
rect 26518 29402 26574 29404
rect 26278 29350 26324 29402
rect 26324 29350 26334 29402
rect 26358 29350 26388 29402
rect 26388 29350 26400 29402
rect 26400 29350 26414 29402
rect 26438 29350 26452 29402
rect 26452 29350 26464 29402
rect 26464 29350 26494 29402
rect 26518 29350 26528 29402
rect 26528 29350 26574 29402
rect 26278 29348 26334 29350
rect 26358 29348 26414 29350
rect 26438 29348 26494 29350
rect 26518 29348 26574 29350
rect 26278 28314 26334 28316
rect 26358 28314 26414 28316
rect 26438 28314 26494 28316
rect 26518 28314 26574 28316
rect 26278 28262 26324 28314
rect 26324 28262 26334 28314
rect 26358 28262 26388 28314
rect 26388 28262 26400 28314
rect 26400 28262 26414 28314
rect 26438 28262 26452 28314
rect 26452 28262 26464 28314
rect 26464 28262 26494 28314
rect 26518 28262 26528 28314
rect 26528 28262 26574 28314
rect 26278 28260 26334 28262
rect 26358 28260 26414 28262
rect 26438 28260 26494 28262
rect 26518 28260 26574 28262
rect 30499 33210 30555 33212
rect 30579 33210 30635 33212
rect 30659 33210 30715 33212
rect 30739 33210 30795 33212
rect 30499 33158 30545 33210
rect 30545 33158 30555 33210
rect 30579 33158 30609 33210
rect 30609 33158 30621 33210
rect 30621 33158 30635 33210
rect 30659 33158 30673 33210
rect 30673 33158 30685 33210
rect 30685 33158 30715 33210
rect 30739 33158 30749 33210
rect 30749 33158 30795 33210
rect 30499 33156 30555 33158
rect 30579 33156 30635 33158
rect 30659 33156 30715 33158
rect 30739 33156 30795 33158
rect 30499 32122 30555 32124
rect 30579 32122 30635 32124
rect 30659 32122 30715 32124
rect 30739 32122 30795 32124
rect 30499 32070 30545 32122
rect 30545 32070 30555 32122
rect 30579 32070 30609 32122
rect 30609 32070 30621 32122
rect 30621 32070 30635 32122
rect 30659 32070 30673 32122
rect 30673 32070 30685 32122
rect 30685 32070 30715 32122
rect 30739 32070 30749 32122
rect 30749 32070 30795 32122
rect 30499 32068 30555 32070
rect 30579 32068 30635 32070
rect 30659 32068 30715 32070
rect 30739 32068 30795 32070
rect 26278 27226 26334 27228
rect 26358 27226 26414 27228
rect 26438 27226 26494 27228
rect 26518 27226 26574 27228
rect 26278 27174 26324 27226
rect 26324 27174 26334 27226
rect 26358 27174 26388 27226
rect 26388 27174 26400 27226
rect 26400 27174 26414 27226
rect 26438 27174 26452 27226
rect 26452 27174 26464 27226
rect 26464 27174 26494 27226
rect 26518 27174 26528 27226
rect 26528 27174 26574 27226
rect 26278 27172 26334 27174
rect 26358 27172 26414 27174
rect 26438 27172 26494 27174
rect 26518 27172 26574 27174
rect 25594 26288 25650 26344
rect 5176 16890 5232 16892
rect 5256 16890 5312 16892
rect 5336 16890 5392 16892
rect 5416 16890 5472 16892
rect 5176 16838 5222 16890
rect 5222 16838 5232 16890
rect 5256 16838 5286 16890
rect 5286 16838 5298 16890
rect 5298 16838 5312 16890
rect 5336 16838 5350 16890
rect 5350 16838 5362 16890
rect 5362 16838 5392 16890
rect 5416 16838 5426 16890
rect 5426 16838 5472 16890
rect 5176 16836 5232 16838
rect 5256 16836 5312 16838
rect 5336 16836 5392 16838
rect 5416 16836 5472 16838
rect 13617 16890 13673 16892
rect 13697 16890 13753 16892
rect 13777 16890 13833 16892
rect 13857 16890 13913 16892
rect 13617 16838 13663 16890
rect 13663 16838 13673 16890
rect 13697 16838 13727 16890
rect 13727 16838 13739 16890
rect 13739 16838 13753 16890
rect 13777 16838 13791 16890
rect 13791 16838 13803 16890
rect 13803 16838 13833 16890
rect 13857 16838 13867 16890
rect 13867 16838 13913 16890
rect 13617 16836 13673 16838
rect 13697 16836 13753 16838
rect 13777 16836 13833 16838
rect 13857 16836 13913 16838
rect 9396 16346 9452 16348
rect 9476 16346 9532 16348
rect 9556 16346 9612 16348
rect 9636 16346 9692 16348
rect 9396 16294 9442 16346
rect 9442 16294 9452 16346
rect 9476 16294 9506 16346
rect 9506 16294 9518 16346
rect 9518 16294 9532 16346
rect 9556 16294 9570 16346
rect 9570 16294 9582 16346
rect 9582 16294 9612 16346
rect 9636 16294 9646 16346
rect 9646 16294 9692 16346
rect 9396 16292 9452 16294
rect 9476 16292 9532 16294
rect 9556 16292 9612 16294
rect 9636 16292 9692 16294
rect 5176 15802 5232 15804
rect 5256 15802 5312 15804
rect 5336 15802 5392 15804
rect 5416 15802 5472 15804
rect 5176 15750 5222 15802
rect 5222 15750 5232 15802
rect 5256 15750 5286 15802
rect 5286 15750 5298 15802
rect 5298 15750 5312 15802
rect 5336 15750 5350 15802
rect 5350 15750 5362 15802
rect 5362 15750 5392 15802
rect 5416 15750 5426 15802
rect 5426 15750 5472 15802
rect 5176 15748 5232 15750
rect 5256 15748 5312 15750
rect 5336 15748 5392 15750
rect 5416 15748 5472 15750
rect 13617 15802 13673 15804
rect 13697 15802 13753 15804
rect 13777 15802 13833 15804
rect 13857 15802 13913 15804
rect 13617 15750 13663 15802
rect 13663 15750 13673 15802
rect 13697 15750 13727 15802
rect 13727 15750 13739 15802
rect 13739 15750 13753 15802
rect 13777 15750 13791 15802
rect 13791 15750 13803 15802
rect 13803 15750 13833 15802
rect 13857 15750 13867 15802
rect 13867 15750 13913 15802
rect 13617 15748 13673 15750
rect 13697 15748 13753 15750
rect 13777 15748 13833 15750
rect 13857 15748 13913 15750
rect 9396 15258 9452 15260
rect 9476 15258 9532 15260
rect 9556 15258 9612 15260
rect 9636 15258 9692 15260
rect 9396 15206 9442 15258
rect 9442 15206 9452 15258
rect 9476 15206 9506 15258
rect 9506 15206 9518 15258
rect 9518 15206 9532 15258
rect 9556 15206 9570 15258
rect 9570 15206 9582 15258
rect 9582 15206 9612 15258
rect 9636 15206 9646 15258
rect 9646 15206 9692 15258
rect 9396 15204 9452 15206
rect 9476 15204 9532 15206
rect 9556 15204 9612 15206
rect 9636 15204 9692 15206
rect 5176 14714 5232 14716
rect 5256 14714 5312 14716
rect 5336 14714 5392 14716
rect 5416 14714 5472 14716
rect 5176 14662 5222 14714
rect 5222 14662 5232 14714
rect 5256 14662 5286 14714
rect 5286 14662 5298 14714
rect 5298 14662 5312 14714
rect 5336 14662 5350 14714
rect 5350 14662 5362 14714
rect 5362 14662 5392 14714
rect 5416 14662 5426 14714
rect 5426 14662 5472 14714
rect 5176 14660 5232 14662
rect 5256 14660 5312 14662
rect 5336 14660 5392 14662
rect 5416 14660 5472 14662
rect 13617 14714 13673 14716
rect 13697 14714 13753 14716
rect 13777 14714 13833 14716
rect 13857 14714 13913 14716
rect 13617 14662 13663 14714
rect 13663 14662 13673 14714
rect 13697 14662 13727 14714
rect 13727 14662 13739 14714
rect 13739 14662 13753 14714
rect 13777 14662 13791 14714
rect 13791 14662 13803 14714
rect 13803 14662 13833 14714
rect 13857 14662 13867 14714
rect 13867 14662 13913 14714
rect 13617 14660 13673 14662
rect 13697 14660 13753 14662
rect 13777 14660 13833 14662
rect 13857 14660 13913 14662
rect 1398 9560 1454 9616
rect 9396 14170 9452 14172
rect 9476 14170 9532 14172
rect 9556 14170 9612 14172
rect 9636 14170 9692 14172
rect 9396 14118 9442 14170
rect 9442 14118 9452 14170
rect 9476 14118 9506 14170
rect 9506 14118 9518 14170
rect 9518 14118 9532 14170
rect 9556 14118 9570 14170
rect 9570 14118 9582 14170
rect 9582 14118 9612 14170
rect 9636 14118 9646 14170
rect 9646 14118 9692 14170
rect 9396 14116 9452 14118
rect 9476 14116 9532 14118
rect 9556 14116 9612 14118
rect 9636 14116 9692 14118
rect 5176 13626 5232 13628
rect 5256 13626 5312 13628
rect 5336 13626 5392 13628
rect 5416 13626 5472 13628
rect 5176 13574 5222 13626
rect 5222 13574 5232 13626
rect 5256 13574 5286 13626
rect 5286 13574 5298 13626
rect 5298 13574 5312 13626
rect 5336 13574 5350 13626
rect 5350 13574 5362 13626
rect 5362 13574 5392 13626
rect 5416 13574 5426 13626
rect 5426 13574 5472 13626
rect 5176 13572 5232 13574
rect 5256 13572 5312 13574
rect 5336 13572 5392 13574
rect 5416 13572 5472 13574
rect 13617 13626 13673 13628
rect 13697 13626 13753 13628
rect 13777 13626 13833 13628
rect 13857 13626 13913 13628
rect 13617 13574 13663 13626
rect 13663 13574 13673 13626
rect 13697 13574 13727 13626
rect 13727 13574 13739 13626
rect 13739 13574 13753 13626
rect 13777 13574 13791 13626
rect 13791 13574 13803 13626
rect 13803 13574 13833 13626
rect 13857 13574 13867 13626
rect 13867 13574 13913 13626
rect 13617 13572 13673 13574
rect 13697 13572 13753 13574
rect 13777 13572 13833 13574
rect 13857 13572 13913 13574
rect 9396 13082 9452 13084
rect 9476 13082 9532 13084
rect 9556 13082 9612 13084
rect 9636 13082 9692 13084
rect 9396 13030 9442 13082
rect 9442 13030 9452 13082
rect 9476 13030 9506 13082
rect 9506 13030 9518 13082
rect 9518 13030 9532 13082
rect 9556 13030 9570 13082
rect 9570 13030 9582 13082
rect 9582 13030 9612 13082
rect 9636 13030 9646 13082
rect 9646 13030 9692 13082
rect 9396 13028 9452 13030
rect 9476 13028 9532 13030
rect 9556 13028 9612 13030
rect 9636 13028 9692 13030
rect 5176 12538 5232 12540
rect 5256 12538 5312 12540
rect 5336 12538 5392 12540
rect 5416 12538 5472 12540
rect 5176 12486 5222 12538
rect 5222 12486 5232 12538
rect 5256 12486 5286 12538
rect 5286 12486 5298 12538
rect 5298 12486 5312 12538
rect 5336 12486 5350 12538
rect 5350 12486 5362 12538
rect 5362 12486 5392 12538
rect 5416 12486 5426 12538
rect 5426 12486 5472 12538
rect 5176 12484 5232 12486
rect 5256 12484 5312 12486
rect 5336 12484 5392 12486
rect 5416 12484 5472 12486
rect 13617 12538 13673 12540
rect 13697 12538 13753 12540
rect 13777 12538 13833 12540
rect 13857 12538 13913 12540
rect 13617 12486 13663 12538
rect 13663 12486 13673 12538
rect 13697 12486 13727 12538
rect 13727 12486 13739 12538
rect 13739 12486 13753 12538
rect 13777 12486 13791 12538
rect 13791 12486 13803 12538
rect 13803 12486 13833 12538
rect 13857 12486 13867 12538
rect 13867 12486 13913 12538
rect 13617 12484 13673 12486
rect 13697 12484 13753 12486
rect 13777 12484 13833 12486
rect 13857 12484 13913 12486
rect 17837 17434 17893 17436
rect 17917 17434 17973 17436
rect 17997 17434 18053 17436
rect 18077 17434 18133 17436
rect 17837 17382 17883 17434
rect 17883 17382 17893 17434
rect 17917 17382 17947 17434
rect 17947 17382 17959 17434
rect 17959 17382 17973 17434
rect 17997 17382 18011 17434
rect 18011 17382 18023 17434
rect 18023 17382 18053 17434
rect 18077 17382 18087 17434
rect 18087 17382 18133 17434
rect 17837 17380 17893 17382
rect 17917 17380 17973 17382
rect 17997 17380 18053 17382
rect 18077 17380 18133 17382
rect 17837 16346 17893 16348
rect 17917 16346 17973 16348
rect 17997 16346 18053 16348
rect 18077 16346 18133 16348
rect 17837 16294 17883 16346
rect 17883 16294 17893 16346
rect 17917 16294 17947 16346
rect 17947 16294 17959 16346
rect 17959 16294 17973 16346
rect 17997 16294 18011 16346
rect 18011 16294 18023 16346
rect 18023 16294 18053 16346
rect 18077 16294 18087 16346
rect 18087 16294 18133 16346
rect 17837 16292 17893 16294
rect 17917 16292 17973 16294
rect 17997 16292 18053 16294
rect 18077 16292 18133 16294
rect 17837 15258 17893 15260
rect 17917 15258 17973 15260
rect 17997 15258 18053 15260
rect 18077 15258 18133 15260
rect 17837 15206 17883 15258
rect 17883 15206 17893 15258
rect 17917 15206 17947 15258
rect 17947 15206 17959 15258
rect 17959 15206 17973 15258
rect 17997 15206 18011 15258
rect 18011 15206 18023 15258
rect 18023 15206 18053 15258
rect 18077 15206 18087 15258
rect 18087 15206 18133 15258
rect 17837 15204 17893 15206
rect 17917 15204 17973 15206
rect 17997 15204 18053 15206
rect 18077 15204 18133 15206
rect 17837 14170 17893 14172
rect 17917 14170 17973 14172
rect 17997 14170 18053 14172
rect 18077 14170 18133 14172
rect 17837 14118 17883 14170
rect 17883 14118 17893 14170
rect 17917 14118 17947 14170
rect 17947 14118 17959 14170
rect 17959 14118 17973 14170
rect 17997 14118 18011 14170
rect 18011 14118 18023 14170
rect 18023 14118 18053 14170
rect 18077 14118 18087 14170
rect 18087 14118 18133 14170
rect 17837 14116 17893 14118
rect 17917 14116 17973 14118
rect 17997 14116 18053 14118
rect 18077 14116 18133 14118
rect 17837 13082 17893 13084
rect 17917 13082 17973 13084
rect 17997 13082 18053 13084
rect 18077 13082 18133 13084
rect 17837 13030 17883 13082
rect 17883 13030 17893 13082
rect 17917 13030 17947 13082
rect 17947 13030 17959 13082
rect 17959 13030 17973 13082
rect 17997 13030 18011 13082
rect 18011 13030 18023 13082
rect 18023 13030 18053 13082
rect 18077 13030 18087 13082
rect 18087 13030 18133 13082
rect 17837 13028 17893 13030
rect 17917 13028 17973 13030
rect 17997 13028 18053 13030
rect 18077 13028 18133 13030
rect 9396 11994 9452 11996
rect 9476 11994 9532 11996
rect 9556 11994 9612 11996
rect 9636 11994 9692 11996
rect 9396 11942 9442 11994
rect 9442 11942 9452 11994
rect 9476 11942 9506 11994
rect 9506 11942 9518 11994
rect 9518 11942 9532 11994
rect 9556 11942 9570 11994
rect 9570 11942 9582 11994
rect 9582 11942 9612 11994
rect 9636 11942 9646 11994
rect 9646 11942 9692 11994
rect 9396 11940 9452 11942
rect 9476 11940 9532 11942
rect 9556 11940 9612 11942
rect 9636 11940 9692 11942
rect 17837 11994 17893 11996
rect 17917 11994 17973 11996
rect 17997 11994 18053 11996
rect 18077 11994 18133 11996
rect 17837 11942 17883 11994
rect 17883 11942 17893 11994
rect 17917 11942 17947 11994
rect 17947 11942 17959 11994
rect 17959 11942 17973 11994
rect 17997 11942 18011 11994
rect 18011 11942 18023 11994
rect 18023 11942 18053 11994
rect 18077 11942 18087 11994
rect 18087 11942 18133 11994
rect 17837 11940 17893 11942
rect 17917 11940 17973 11942
rect 17997 11940 18053 11942
rect 18077 11940 18133 11942
rect 5176 11450 5232 11452
rect 5256 11450 5312 11452
rect 5336 11450 5392 11452
rect 5416 11450 5472 11452
rect 5176 11398 5222 11450
rect 5222 11398 5232 11450
rect 5256 11398 5286 11450
rect 5286 11398 5298 11450
rect 5298 11398 5312 11450
rect 5336 11398 5350 11450
rect 5350 11398 5362 11450
rect 5362 11398 5392 11450
rect 5416 11398 5426 11450
rect 5426 11398 5472 11450
rect 5176 11396 5232 11398
rect 5256 11396 5312 11398
rect 5336 11396 5392 11398
rect 5416 11396 5472 11398
rect 13617 11450 13673 11452
rect 13697 11450 13753 11452
rect 13777 11450 13833 11452
rect 13857 11450 13913 11452
rect 13617 11398 13663 11450
rect 13663 11398 13673 11450
rect 13697 11398 13727 11450
rect 13727 11398 13739 11450
rect 13739 11398 13753 11450
rect 13777 11398 13791 11450
rect 13791 11398 13803 11450
rect 13803 11398 13833 11450
rect 13857 11398 13867 11450
rect 13867 11398 13913 11450
rect 13617 11396 13673 11398
rect 13697 11396 13753 11398
rect 13777 11396 13833 11398
rect 13857 11396 13913 11398
rect 9396 10906 9452 10908
rect 9476 10906 9532 10908
rect 9556 10906 9612 10908
rect 9636 10906 9692 10908
rect 9396 10854 9442 10906
rect 9442 10854 9452 10906
rect 9476 10854 9506 10906
rect 9506 10854 9518 10906
rect 9518 10854 9532 10906
rect 9556 10854 9570 10906
rect 9570 10854 9582 10906
rect 9582 10854 9612 10906
rect 9636 10854 9646 10906
rect 9646 10854 9692 10906
rect 9396 10852 9452 10854
rect 9476 10852 9532 10854
rect 9556 10852 9612 10854
rect 9636 10852 9692 10854
rect 17837 10906 17893 10908
rect 17917 10906 17973 10908
rect 17997 10906 18053 10908
rect 18077 10906 18133 10908
rect 17837 10854 17883 10906
rect 17883 10854 17893 10906
rect 17917 10854 17947 10906
rect 17947 10854 17959 10906
rect 17959 10854 17973 10906
rect 17997 10854 18011 10906
rect 18011 10854 18023 10906
rect 18023 10854 18053 10906
rect 18077 10854 18087 10906
rect 18087 10854 18133 10906
rect 17837 10852 17893 10854
rect 17917 10852 17973 10854
rect 17997 10852 18053 10854
rect 18077 10852 18133 10854
rect 5176 10362 5232 10364
rect 5256 10362 5312 10364
rect 5336 10362 5392 10364
rect 5416 10362 5472 10364
rect 5176 10310 5222 10362
rect 5222 10310 5232 10362
rect 5256 10310 5286 10362
rect 5286 10310 5298 10362
rect 5298 10310 5312 10362
rect 5336 10310 5350 10362
rect 5350 10310 5362 10362
rect 5362 10310 5392 10362
rect 5416 10310 5426 10362
rect 5426 10310 5472 10362
rect 5176 10308 5232 10310
rect 5256 10308 5312 10310
rect 5336 10308 5392 10310
rect 5416 10308 5472 10310
rect 13617 10362 13673 10364
rect 13697 10362 13753 10364
rect 13777 10362 13833 10364
rect 13857 10362 13913 10364
rect 13617 10310 13663 10362
rect 13663 10310 13673 10362
rect 13697 10310 13727 10362
rect 13727 10310 13739 10362
rect 13739 10310 13753 10362
rect 13777 10310 13791 10362
rect 13791 10310 13803 10362
rect 13803 10310 13833 10362
rect 13857 10310 13867 10362
rect 13867 10310 13913 10362
rect 13617 10308 13673 10310
rect 13697 10308 13753 10310
rect 13777 10308 13833 10310
rect 13857 10308 13913 10310
rect 9396 9818 9452 9820
rect 9476 9818 9532 9820
rect 9556 9818 9612 9820
rect 9636 9818 9692 9820
rect 9396 9766 9442 9818
rect 9442 9766 9452 9818
rect 9476 9766 9506 9818
rect 9506 9766 9518 9818
rect 9518 9766 9532 9818
rect 9556 9766 9570 9818
rect 9570 9766 9582 9818
rect 9582 9766 9612 9818
rect 9636 9766 9646 9818
rect 9646 9766 9692 9818
rect 9396 9764 9452 9766
rect 9476 9764 9532 9766
rect 9556 9764 9612 9766
rect 9636 9764 9692 9766
rect 17837 9818 17893 9820
rect 17917 9818 17973 9820
rect 17997 9818 18053 9820
rect 18077 9818 18133 9820
rect 17837 9766 17883 9818
rect 17883 9766 17893 9818
rect 17917 9766 17947 9818
rect 17947 9766 17959 9818
rect 17959 9766 17973 9818
rect 17997 9766 18011 9818
rect 18011 9766 18023 9818
rect 18023 9766 18053 9818
rect 18077 9766 18087 9818
rect 18087 9766 18133 9818
rect 17837 9764 17893 9766
rect 17917 9764 17973 9766
rect 17997 9764 18053 9766
rect 18077 9764 18133 9766
rect 5176 9274 5232 9276
rect 5256 9274 5312 9276
rect 5336 9274 5392 9276
rect 5416 9274 5472 9276
rect 5176 9222 5222 9274
rect 5222 9222 5232 9274
rect 5256 9222 5286 9274
rect 5286 9222 5298 9274
rect 5298 9222 5312 9274
rect 5336 9222 5350 9274
rect 5350 9222 5362 9274
rect 5362 9222 5392 9274
rect 5416 9222 5426 9274
rect 5426 9222 5472 9274
rect 5176 9220 5232 9222
rect 5256 9220 5312 9222
rect 5336 9220 5392 9222
rect 5416 9220 5472 9222
rect 13617 9274 13673 9276
rect 13697 9274 13753 9276
rect 13777 9274 13833 9276
rect 13857 9274 13913 9276
rect 13617 9222 13663 9274
rect 13663 9222 13673 9274
rect 13697 9222 13727 9274
rect 13727 9222 13739 9274
rect 13739 9222 13753 9274
rect 13777 9222 13791 9274
rect 13791 9222 13803 9274
rect 13803 9222 13833 9274
rect 13857 9222 13867 9274
rect 13867 9222 13913 9274
rect 13617 9220 13673 9222
rect 13697 9220 13753 9222
rect 13777 9220 13833 9222
rect 13857 9220 13913 9222
rect 9396 8730 9452 8732
rect 9476 8730 9532 8732
rect 9556 8730 9612 8732
rect 9636 8730 9692 8732
rect 9396 8678 9442 8730
rect 9442 8678 9452 8730
rect 9476 8678 9506 8730
rect 9506 8678 9518 8730
rect 9518 8678 9532 8730
rect 9556 8678 9570 8730
rect 9570 8678 9582 8730
rect 9582 8678 9612 8730
rect 9636 8678 9646 8730
rect 9646 8678 9692 8730
rect 9396 8676 9452 8678
rect 9476 8676 9532 8678
rect 9556 8676 9612 8678
rect 9636 8676 9692 8678
rect 17837 8730 17893 8732
rect 17917 8730 17973 8732
rect 17997 8730 18053 8732
rect 18077 8730 18133 8732
rect 17837 8678 17883 8730
rect 17883 8678 17893 8730
rect 17917 8678 17947 8730
rect 17947 8678 17959 8730
rect 17959 8678 17973 8730
rect 17997 8678 18011 8730
rect 18011 8678 18023 8730
rect 18023 8678 18053 8730
rect 18077 8678 18087 8730
rect 18087 8678 18133 8730
rect 17837 8676 17893 8678
rect 17917 8676 17973 8678
rect 17997 8676 18053 8678
rect 18077 8676 18133 8678
rect 5176 8186 5232 8188
rect 5256 8186 5312 8188
rect 5336 8186 5392 8188
rect 5416 8186 5472 8188
rect 5176 8134 5222 8186
rect 5222 8134 5232 8186
rect 5256 8134 5286 8186
rect 5286 8134 5298 8186
rect 5298 8134 5312 8186
rect 5336 8134 5350 8186
rect 5350 8134 5362 8186
rect 5362 8134 5392 8186
rect 5416 8134 5426 8186
rect 5426 8134 5472 8186
rect 5176 8132 5232 8134
rect 5256 8132 5312 8134
rect 5336 8132 5392 8134
rect 5416 8132 5472 8134
rect 13617 8186 13673 8188
rect 13697 8186 13753 8188
rect 13777 8186 13833 8188
rect 13857 8186 13913 8188
rect 13617 8134 13663 8186
rect 13663 8134 13673 8186
rect 13697 8134 13727 8186
rect 13727 8134 13739 8186
rect 13739 8134 13753 8186
rect 13777 8134 13791 8186
rect 13791 8134 13803 8186
rect 13803 8134 13833 8186
rect 13857 8134 13867 8186
rect 13867 8134 13913 8186
rect 13617 8132 13673 8134
rect 13697 8132 13753 8134
rect 13777 8132 13833 8134
rect 13857 8132 13913 8134
rect 9396 7642 9452 7644
rect 9476 7642 9532 7644
rect 9556 7642 9612 7644
rect 9636 7642 9692 7644
rect 9396 7590 9442 7642
rect 9442 7590 9452 7642
rect 9476 7590 9506 7642
rect 9506 7590 9518 7642
rect 9518 7590 9532 7642
rect 9556 7590 9570 7642
rect 9570 7590 9582 7642
rect 9582 7590 9612 7642
rect 9636 7590 9646 7642
rect 9646 7590 9692 7642
rect 9396 7588 9452 7590
rect 9476 7588 9532 7590
rect 9556 7588 9612 7590
rect 9636 7588 9692 7590
rect 17837 7642 17893 7644
rect 17917 7642 17973 7644
rect 17997 7642 18053 7644
rect 18077 7642 18133 7644
rect 17837 7590 17883 7642
rect 17883 7590 17893 7642
rect 17917 7590 17947 7642
rect 17947 7590 17959 7642
rect 17959 7590 17973 7642
rect 17997 7590 18011 7642
rect 18011 7590 18023 7642
rect 18023 7590 18053 7642
rect 18077 7590 18087 7642
rect 18087 7590 18133 7642
rect 17837 7588 17893 7590
rect 17917 7588 17973 7590
rect 17997 7588 18053 7590
rect 18077 7588 18133 7590
rect 5176 7098 5232 7100
rect 5256 7098 5312 7100
rect 5336 7098 5392 7100
rect 5416 7098 5472 7100
rect 5176 7046 5222 7098
rect 5222 7046 5232 7098
rect 5256 7046 5286 7098
rect 5286 7046 5298 7098
rect 5298 7046 5312 7098
rect 5336 7046 5350 7098
rect 5350 7046 5362 7098
rect 5362 7046 5392 7098
rect 5416 7046 5426 7098
rect 5426 7046 5472 7098
rect 5176 7044 5232 7046
rect 5256 7044 5312 7046
rect 5336 7044 5392 7046
rect 5416 7044 5472 7046
rect 13617 7098 13673 7100
rect 13697 7098 13753 7100
rect 13777 7098 13833 7100
rect 13857 7098 13913 7100
rect 13617 7046 13663 7098
rect 13663 7046 13673 7098
rect 13697 7046 13727 7098
rect 13727 7046 13739 7098
rect 13739 7046 13753 7098
rect 13777 7046 13791 7098
rect 13791 7046 13803 7098
rect 13803 7046 13833 7098
rect 13857 7046 13867 7098
rect 13867 7046 13913 7098
rect 13617 7044 13673 7046
rect 13697 7044 13753 7046
rect 13777 7044 13833 7046
rect 13857 7044 13913 7046
rect 22058 22330 22114 22332
rect 22138 22330 22194 22332
rect 22218 22330 22274 22332
rect 22298 22330 22354 22332
rect 22058 22278 22104 22330
rect 22104 22278 22114 22330
rect 22138 22278 22168 22330
rect 22168 22278 22180 22330
rect 22180 22278 22194 22330
rect 22218 22278 22232 22330
rect 22232 22278 22244 22330
rect 22244 22278 22274 22330
rect 22298 22278 22308 22330
rect 22308 22278 22354 22330
rect 22058 22276 22114 22278
rect 22138 22276 22194 22278
rect 22218 22276 22274 22278
rect 22298 22276 22354 22278
rect 22058 21242 22114 21244
rect 22138 21242 22194 21244
rect 22218 21242 22274 21244
rect 22298 21242 22354 21244
rect 22058 21190 22104 21242
rect 22104 21190 22114 21242
rect 22138 21190 22168 21242
rect 22168 21190 22180 21242
rect 22180 21190 22194 21242
rect 22218 21190 22232 21242
rect 22232 21190 22244 21242
rect 22244 21190 22274 21242
rect 22298 21190 22308 21242
rect 22308 21190 22354 21242
rect 22058 21188 22114 21190
rect 22138 21188 22194 21190
rect 22218 21188 22274 21190
rect 22298 21188 22354 21190
rect 22058 20154 22114 20156
rect 22138 20154 22194 20156
rect 22218 20154 22274 20156
rect 22298 20154 22354 20156
rect 22058 20102 22104 20154
rect 22104 20102 22114 20154
rect 22138 20102 22168 20154
rect 22168 20102 22180 20154
rect 22180 20102 22194 20154
rect 22218 20102 22232 20154
rect 22232 20102 22244 20154
rect 22244 20102 22274 20154
rect 22298 20102 22308 20154
rect 22308 20102 22354 20154
rect 22058 20100 22114 20102
rect 22138 20100 22194 20102
rect 22218 20100 22274 20102
rect 22298 20100 22354 20102
rect 22058 19066 22114 19068
rect 22138 19066 22194 19068
rect 22218 19066 22274 19068
rect 22298 19066 22354 19068
rect 22058 19014 22104 19066
rect 22104 19014 22114 19066
rect 22138 19014 22168 19066
rect 22168 19014 22180 19066
rect 22180 19014 22194 19066
rect 22218 19014 22232 19066
rect 22232 19014 22244 19066
rect 22244 19014 22274 19066
rect 22298 19014 22308 19066
rect 22308 19014 22354 19066
rect 22058 19012 22114 19014
rect 22138 19012 22194 19014
rect 22218 19012 22274 19014
rect 22298 19012 22354 19014
rect 22058 17978 22114 17980
rect 22138 17978 22194 17980
rect 22218 17978 22274 17980
rect 22298 17978 22354 17980
rect 22058 17926 22104 17978
rect 22104 17926 22114 17978
rect 22138 17926 22168 17978
rect 22168 17926 22180 17978
rect 22180 17926 22194 17978
rect 22218 17926 22232 17978
rect 22232 17926 22244 17978
rect 22244 17926 22274 17978
rect 22298 17926 22308 17978
rect 22308 17926 22354 17978
rect 22058 17924 22114 17926
rect 22138 17924 22194 17926
rect 22218 17924 22274 17926
rect 22298 17924 22354 17926
rect 22058 16890 22114 16892
rect 22138 16890 22194 16892
rect 22218 16890 22274 16892
rect 22298 16890 22354 16892
rect 22058 16838 22104 16890
rect 22104 16838 22114 16890
rect 22138 16838 22168 16890
rect 22168 16838 22180 16890
rect 22180 16838 22194 16890
rect 22218 16838 22232 16890
rect 22232 16838 22244 16890
rect 22244 16838 22274 16890
rect 22298 16838 22308 16890
rect 22308 16838 22354 16890
rect 22058 16836 22114 16838
rect 22138 16836 22194 16838
rect 22218 16836 22274 16838
rect 22298 16836 22354 16838
rect 22058 15802 22114 15804
rect 22138 15802 22194 15804
rect 22218 15802 22274 15804
rect 22298 15802 22354 15804
rect 22058 15750 22104 15802
rect 22104 15750 22114 15802
rect 22138 15750 22168 15802
rect 22168 15750 22180 15802
rect 22180 15750 22194 15802
rect 22218 15750 22232 15802
rect 22232 15750 22244 15802
rect 22244 15750 22274 15802
rect 22298 15750 22308 15802
rect 22308 15750 22354 15802
rect 22058 15748 22114 15750
rect 22138 15748 22194 15750
rect 22218 15748 22274 15750
rect 22298 15748 22354 15750
rect 26278 26138 26334 26140
rect 26358 26138 26414 26140
rect 26438 26138 26494 26140
rect 26518 26138 26574 26140
rect 26278 26086 26324 26138
rect 26324 26086 26334 26138
rect 26358 26086 26388 26138
rect 26388 26086 26400 26138
rect 26400 26086 26414 26138
rect 26438 26086 26452 26138
rect 26452 26086 26464 26138
rect 26464 26086 26494 26138
rect 26518 26086 26528 26138
rect 26528 26086 26574 26138
rect 26278 26084 26334 26086
rect 26358 26084 26414 26086
rect 26438 26084 26494 26086
rect 26518 26084 26574 26086
rect 30499 31034 30555 31036
rect 30579 31034 30635 31036
rect 30659 31034 30715 31036
rect 30739 31034 30795 31036
rect 30499 30982 30545 31034
rect 30545 30982 30555 31034
rect 30579 30982 30609 31034
rect 30609 30982 30621 31034
rect 30621 30982 30635 31034
rect 30659 30982 30673 31034
rect 30673 30982 30685 31034
rect 30685 30982 30715 31034
rect 30739 30982 30749 31034
rect 30749 30982 30795 31034
rect 30499 30980 30555 30982
rect 30579 30980 30635 30982
rect 30659 30980 30715 30982
rect 30739 30980 30795 30982
rect 30499 29946 30555 29948
rect 30579 29946 30635 29948
rect 30659 29946 30715 29948
rect 30739 29946 30795 29948
rect 30499 29894 30545 29946
rect 30545 29894 30555 29946
rect 30579 29894 30609 29946
rect 30609 29894 30621 29946
rect 30621 29894 30635 29946
rect 30659 29894 30673 29946
rect 30673 29894 30685 29946
rect 30685 29894 30715 29946
rect 30739 29894 30749 29946
rect 30749 29894 30795 29946
rect 30499 29892 30555 29894
rect 30579 29892 30635 29894
rect 30659 29892 30715 29894
rect 30739 29892 30795 29894
rect 30499 28858 30555 28860
rect 30579 28858 30635 28860
rect 30659 28858 30715 28860
rect 30739 28858 30795 28860
rect 30499 28806 30545 28858
rect 30545 28806 30555 28858
rect 30579 28806 30609 28858
rect 30609 28806 30621 28858
rect 30621 28806 30635 28858
rect 30659 28806 30673 28858
rect 30673 28806 30685 28858
rect 30685 28806 30715 28858
rect 30739 28806 30749 28858
rect 30749 28806 30795 28858
rect 30499 28804 30555 28806
rect 30579 28804 30635 28806
rect 30659 28804 30715 28806
rect 30739 28804 30795 28806
rect 30499 27770 30555 27772
rect 30579 27770 30635 27772
rect 30659 27770 30715 27772
rect 30739 27770 30795 27772
rect 30499 27718 30545 27770
rect 30545 27718 30555 27770
rect 30579 27718 30609 27770
rect 30609 27718 30621 27770
rect 30621 27718 30635 27770
rect 30659 27718 30673 27770
rect 30673 27718 30685 27770
rect 30685 27718 30715 27770
rect 30739 27718 30749 27770
rect 30749 27718 30795 27770
rect 30499 27716 30555 27718
rect 30579 27716 30635 27718
rect 30659 27716 30715 27718
rect 30739 27716 30795 27718
rect 26278 25050 26334 25052
rect 26358 25050 26414 25052
rect 26438 25050 26494 25052
rect 26518 25050 26574 25052
rect 26278 24998 26324 25050
rect 26324 24998 26334 25050
rect 26358 24998 26388 25050
rect 26388 24998 26400 25050
rect 26400 24998 26414 25050
rect 26438 24998 26452 25050
rect 26452 24998 26464 25050
rect 26464 24998 26494 25050
rect 26518 24998 26528 25050
rect 26528 24998 26574 25050
rect 26278 24996 26334 24998
rect 26358 24996 26414 24998
rect 26438 24996 26494 24998
rect 26518 24996 26574 24998
rect 26278 23962 26334 23964
rect 26358 23962 26414 23964
rect 26438 23962 26494 23964
rect 26518 23962 26574 23964
rect 26278 23910 26324 23962
rect 26324 23910 26334 23962
rect 26358 23910 26388 23962
rect 26388 23910 26400 23962
rect 26400 23910 26414 23962
rect 26438 23910 26452 23962
rect 26452 23910 26464 23962
rect 26464 23910 26494 23962
rect 26518 23910 26528 23962
rect 26528 23910 26574 23962
rect 26278 23908 26334 23910
rect 26358 23908 26414 23910
rect 26438 23908 26494 23910
rect 26518 23908 26574 23910
rect 26278 22874 26334 22876
rect 26358 22874 26414 22876
rect 26438 22874 26494 22876
rect 26518 22874 26574 22876
rect 26278 22822 26324 22874
rect 26324 22822 26334 22874
rect 26358 22822 26388 22874
rect 26388 22822 26400 22874
rect 26400 22822 26414 22874
rect 26438 22822 26452 22874
rect 26452 22822 26464 22874
rect 26464 22822 26494 22874
rect 26518 22822 26528 22874
rect 26528 22822 26574 22874
rect 26278 22820 26334 22822
rect 26358 22820 26414 22822
rect 26438 22820 26494 22822
rect 26518 22820 26574 22822
rect 22058 14714 22114 14716
rect 22138 14714 22194 14716
rect 22218 14714 22274 14716
rect 22298 14714 22354 14716
rect 22058 14662 22104 14714
rect 22104 14662 22114 14714
rect 22138 14662 22168 14714
rect 22168 14662 22180 14714
rect 22180 14662 22194 14714
rect 22218 14662 22232 14714
rect 22232 14662 22244 14714
rect 22244 14662 22274 14714
rect 22298 14662 22308 14714
rect 22308 14662 22354 14714
rect 22058 14660 22114 14662
rect 22138 14660 22194 14662
rect 22218 14660 22274 14662
rect 22298 14660 22354 14662
rect 26278 21786 26334 21788
rect 26358 21786 26414 21788
rect 26438 21786 26494 21788
rect 26518 21786 26574 21788
rect 26278 21734 26324 21786
rect 26324 21734 26334 21786
rect 26358 21734 26388 21786
rect 26388 21734 26400 21786
rect 26400 21734 26414 21786
rect 26438 21734 26452 21786
rect 26452 21734 26464 21786
rect 26464 21734 26494 21786
rect 26518 21734 26528 21786
rect 26528 21734 26574 21786
rect 26278 21732 26334 21734
rect 26358 21732 26414 21734
rect 26438 21732 26494 21734
rect 26518 21732 26574 21734
rect 26278 20698 26334 20700
rect 26358 20698 26414 20700
rect 26438 20698 26494 20700
rect 26518 20698 26574 20700
rect 26278 20646 26324 20698
rect 26324 20646 26334 20698
rect 26358 20646 26388 20698
rect 26388 20646 26400 20698
rect 26400 20646 26414 20698
rect 26438 20646 26452 20698
rect 26452 20646 26464 20698
rect 26464 20646 26494 20698
rect 26518 20646 26528 20698
rect 26528 20646 26574 20698
rect 26278 20644 26334 20646
rect 26358 20644 26414 20646
rect 26438 20644 26494 20646
rect 26518 20644 26574 20646
rect 26278 19610 26334 19612
rect 26358 19610 26414 19612
rect 26438 19610 26494 19612
rect 26518 19610 26574 19612
rect 26278 19558 26324 19610
rect 26324 19558 26334 19610
rect 26358 19558 26388 19610
rect 26388 19558 26400 19610
rect 26400 19558 26414 19610
rect 26438 19558 26452 19610
rect 26452 19558 26464 19610
rect 26464 19558 26494 19610
rect 26518 19558 26528 19610
rect 26528 19558 26574 19610
rect 26278 19556 26334 19558
rect 26358 19556 26414 19558
rect 26438 19556 26494 19558
rect 26518 19556 26574 19558
rect 26278 18522 26334 18524
rect 26358 18522 26414 18524
rect 26438 18522 26494 18524
rect 26518 18522 26574 18524
rect 26278 18470 26324 18522
rect 26324 18470 26334 18522
rect 26358 18470 26388 18522
rect 26388 18470 26400 18522
rect 26400 18470 26414 18522
rect 26438 18470 26452 18522
rect 26452 18470 26464 18522
rect 26464 18470 26494 18522
rect 26518 18470 26528 18522
rect 26528 18470 26574 18522
rect 26278 18468 26334 18470
rect 26358 18468 26414 18470
rect 26438 18468 26494 18470
rect 26518 18468 26574 18470
rect 30499 26682 30555 26684
rect 30579 26682 30635 26684
rect 30659 26682 30715 26684
rect 30739 26682 30795 26684
rect 30499 26630 30545 26682
rect 30545 26630 30555 26682
rect 30579 26630 30609 26682
rect 30609 26630 30621 26682
rect 30621 26630 30635 26682
rect 30659 26630 30673 26682
rect 30673 26630 30685 26682
rect 30685 26630 30715 26682
rect 30739 26630 30749 26682
rect 30749 26630 30795 26682
rect 30499 26628 30555 26630
rect 30579 26628 30635 26630
rect 30659 26628 30715 26630
rect 30739 26628 30795 26630
rect 34719 39194 34775 39196
rect 34799 39194 34855 39196
rect 34879 39194 34935 39196
rect 34959 39194 35015 39196
rect 34719 39142 34765 39194
rect 34765 39142 34775 39194
rect 34799 39142 34829 39194
rect 34829 39142 34841 39194
rect 34841 39142 34855 39194
rect 34879 39142 34893 39194
rect 34893 39142 34905 39194
rect 34905 39142 34935 39194
rect 34959 39142 34969 39194
rect 34969 39142 35015 39194
rect 34719 39140 34775 39142
rect 34799 39140 34855 39142
rect 34879 39140 34935 39142
rect 34959 39140 35015 39142
rect 34719 38106 34775 38108
rect 34799 38106 34855 38108
rect 34879 38106 34935 38108
rect 34959 38106 35015 38108
rect 34719 38054 34765 38106
rect 34765 38054 34775 38106
rect 34799 38054 34829 38106
rect 34829 38054 34841 38106
rect 34841 38054 34855 38106
rect 34879 38054 34893 38106
rect 34893 38054 34905 38106
rect 34905 38054 34935 38106
rect 34959 38054 34969 38106
rect 34969 38054 35015 38106
rect 34719 38052 34775 38054
rect 34799 38052 34855 38054
rect 34879 38052 34935 38054
rect 34959 38052 35015 38054
rect 34719 37018 34775 37020
rect 34799 37018 34855 37020
rect 34879 37018 34935 37020
rect 34959 37018 35015 37020
rect 34719 36966 34765 37018
rect 34765 36966 34775 37018
rect 34799 36966 34829 37018
rect 34829 36966 34841 37018
rect 34841 36966 34855 37018
rect 34879 36966 34893 37018
rect 34893 36966 34905 37018
rect 34905 36966 34935 37018
rect 34959 36966 34969 37018
rect 34969 36966 35015 37018
rect 34719 36964 34775 36966
rect 34799 36964 34855 36966
rect 34879 36964 34935 36966
rect 34959 36964 35015 36966
rect 34719 35930 34775 35932
rect 34799 35930 34855 35932
rect 34879 35930 34935 35932
rect 34959 35930 35015 35932
rect 34719 35878 34765 35930
rect 34765 35878 34775 35930
rect 34799 35878 34829 35930
rect 34829 35878 34841 35930
rect 34841 35878 34855 35930
rect 34879 35878 34893 35930
rect 34893 35878 34905 35930
rect 34905 35878 34935 35930
rect 34959 35878 34969 35930
rect 34969 35878 35015 35930
rect 34719 35876 34775 35878
rect 34799 35876 34855 35878
rect 34879 35876 34935 35878
rect 34959 35876 35015 35878
rect 34719 34842 34775 34844
rect 34799 34842 34855 34844
rect 34879 34842 34935 34844
rect 34959 34842 35015 34844
rect 34719 34790 34765 34842
rect 34765 34790 34775 34842
rect 34799 34790 34829 34842
rect 34829 34790 34841 34842
rect 34841 34790 34855 34842
rect 34879 34790 34893 34842
rect 34893 34790 34905 34842
rect 34905 34790 34935 34842
rect 34959 34790 34969 34842
rect 34969 34790 35015 34842
rect 34719 34788 34775 34790
rect 34799 34788 34855 34790
rect 34879 34788 34935 34790
rect 34959 34788 35015 34790
rect 34719 33754 34775 33756
rect 34799 33754 34855 33756
rect 34879 33754 34935 33756
rect 34959 33754 35015 33756
rect 34719 33702 34765 33754
rect 34765 33702 34775 33754
rect 34799 33702 34829 33754
rect 34829 33702 34841 33754
rect 34841 33702 34855 33754
rect 34879 33702 34893 33754
rect 34893 33702 34905 33754
rect 34905 33702 34935 33754
rect 34959 33702 34969 33754
rect 34969 33702 35015 33754
rect 34719 33700 34775 33702
rect 34799 33700 34855 33702
rect 34879 33700 34935 33702
rect 34959 33700 35015 33702
rect 34719 32666 34775 32668
rect 34799 32666 34855 32668
rect 34879 32666 34935 32668
rect 34959 32666 35015 32668
rect 34719 32614 34765 32666
rect 34765 32614 34775 32666
rect 34799 32614 34829 32666
rect 34829 32614 34841 32666
rect 34841 32614 34855 32666
rect 34879 32614 34893 32666
rect 34893 32614 34905 32666
rect 34905 32614 34935 32666
rect 34959 32614 34969 32666
rect 34969 32614 35015 32666
rect 34719 32612 34775 32614
rect 34799 32612 34855 32614
rect 34879 32612 34935 32614
rect 34959 32612 35015 32614
rect 34886 32000 34942 32056
rect 34719 31578 34775 31580
rect 34799 31578 34855 31580
rect 34879 31578 34935 31580
rect 34959 31578 35015 31580
rect 34719 31526 34765 31578
rect 34765 31526 34775 31578
rect 34799 31526 34829 31578
rect 34829 31526 34841 31578
rect 34841 31526 34855 31578
rect 34879 31526 34893 31578
rect 34893 31526 34905 31578
rect 34905 31526 34935 31578
rect 34959 31526 34969 31578
rect 34969 31526 35015 31578
rect 34719 31524 34775 31526
rect 34799 31524 34855 31526
rect 34879 31524 34935 31526
rect 34959 31524 35015 31526
rect 34719 30490 34775 30492
rect 34799 30490 34855 30492
rect 34879 30490 34935 30492
rect 34959 30490 35015 30492
rect 34719 30438 34765 30490
rect 34765 30438 34775 30490
rect 34799 30438 34829 30490
rect 34829 30438 34841 30490
rect 34841 30438 34855 30490
rect 34879 30438 34893 30490
rect 34893 30438 34905 30490
rect 34905 30438 34935 30490
rect 34959 30438 34969 30490
rect 34969 30438 35015 30490
rect 34719 30436 34775 30438
rect 34799 30436 34855 30438
rect 34879 30436 34935 30438
rect 34959 30436 35015 30438
rect 34719 29402 34775 29404
rect 34799 29402 34855 29404
rect 34879 29402 34935 29404
rect 34959 29402 35015 29404
rect 34719 29350 34765 29402
rect 34765 29350 34775 29402
rect 34799 29350 34829 29402
rect 34829 29350 34841 29402
rect 34841 29350 34855 29402
rect 34879 29350 34893 29402
rect 34893 29350 34905 29402
rect 34905 29350 34935 29402
rect 34959 29350 34969 29402
rect 34969 29350 35015 29402
rect 34719 29348 34775 29350
rect 34799 29348 34855 29350
rect 34879 29348 34935 29350
rect 34959 29348 35015 29350
rect 34719 28314 34775 28316
rect 34799 28314 34855 28316
rect 34879 28314 34935 28316
rect 34959 28314 35015 28316
rect 34719 28262 34765 28314
rect 34765 28262 34775 28314
rect 34799 28262 34829 28314
rect 34829 28262 34841 28314
rect 34841 28262 34855 28314
rect 34879 28262 34893 28314
rect 34893 28262 34905 28314
rect 34905 28262 34935 28314
rect 34959 28262 34969 28314
rect 34969 28262 35015 28314
rect 34719 28260 34775 28262
rect 34799 28260 34855 28262
rect 34879 28260 34935 28262
rect 34959 28260 35015 28262
rect 29090 25220 29146 25256
rect 29090 25200 29092 25220
rect 29092 25200 29144 25220
rect 29144 25200 29146 25220
rect 30102 25236 30104 25256
rect 30104 25236 30156 25256
rect 30156 25236 30158 25256
rect 30102 25200 30158 25236
rect 30499 25594 30555 25596
rect 30579 25594 30635 25596
rect 30659 25594 30715 25596
rect 30739 25594 30795 25596
rect 30499 25542 30545 25594
rect 30545 25542 30555 25594
rect 30579 25542 30609 25594
rect 30609 25542 30621 25594
rect 30621 25542 30635 25594
rect 30659 25542 30673 25594
rect 30673 25542 30685 25594
rect 30685 25542 30715 25594
rect 30739 25542 30749 25594
rect 30749 25542 30795 25594
rect 30499 25540 30555 25542
rect 30579 25540 30635 25542
rect 30659 25540 30715 25542
rect 30739 25540 30795 25542
rect 30499 24506 30555 24508
rect 30579 24506 30635 24508
rect 30659 24506 30715 24508
rect 30739 24506 30795 24508
rect 30499 24454 30545 24506
rect 30545 24454 30555 24506
rect 30579 24454 30609 24506
rect 30609 24454 30621 24506
rect 30621 24454 30635 24506
rect 30659 24454 30673 24506
rect 30673 24454 30685 24506
rect 30685 24454 30715 24506
rect 30739 24454 30749 24506
rect 30749 24454 30795 24506
rect 30499 24452 30555 24454
rect 30579 24452 30635 24454
rect 30659 24452 30715 24454
rect 30739 24452 30795 24454
rect 30499 23418 30555 23420
rect 30579 23418 30635 23420
rect 30659 23418 30715 23420
rect 30739 23418 30795 23420
rect 30499 23366 30545 23418
rect 30545 23366 30555 23418
rect 30579 23366 30609 23418
rect 30609 23366 30621 23418
rect 30621 23366 30635 23418
rect 30659 23366 30673 23418
rect 30673 23366 30685 23418
rect 30685 23366 30715 23418
rect 30739 23366 30749 23418
rect 30749 23366 30795 23418
rect 30499 23364 30555 23366
rect 30579 23364 30635 23366
rect 30659 23364 30715 23366
rect 30739 23364 30795 23366
rect 30499 22330 30555 22332
rect 30579 22330 30635 22332
rect 30659 22330 30715 22332
rect 30739 22330 30795 22332
rect 30499 22278 30545 22330
rect 30545 22278 30555 22330
rect 30579 22278 30609 22330
rect 30609 22278 30621 22330
rect 30621 22278 30635 22330
rect 30659 22278 30673 22330
rect 30673 22278 30685 22330
rect 30685 22278 30715 22330
rect 30739 22278 30749 22330
rect 30749 22278 30795 22330
rect 30499 22276 30555 22278
rect 30579 22276 30635 22278
rect 30659 22276 30715 22278
rect 30739 22276 30795 22278
rect 30499 21242 30555 21244
rect 30579 21242 30635 21244
rect 30659 21242 30715 21244
rect 30739 21242 30795 21244
rect 30499 21190 30545 21242
rect 30545 21190 30555 21242
rect 30579 21190 30609 21242
rect 30609 21190 30621 21242
rect 30621 21190 30635 21242
rect 30659 21190 30673 21242
rect 30673 21190 30685 21242
rect 30685 21190 30715 21242
rect 30739 21190 30749 21242
rect 30749 21190 30795 21242
rect 30499 21188 30555 21190
rect 30579 21188 30635 21190
rect 30659 21188 30715 21190
rect 30739 21188 30795 21190
rect 34719 27226 34775 27228
rect 34799 27226 34855 27228
rect 34879 27226 34935 27228
rect 34959 27226 35015 27228
rect 34719 27174 34765 27226
rect 34765 27174 34775 27226
rect 34799 27174 34829 27226
rect 34829 27174 34841 27226
rect 34841 27174 34855 27226
rect 34879 27174 34893 27226
rect 34893 27174 34905 27226
rect 34905 27174 34935 27226
rect 34959 27174 34969 27226
rect 34969 27174 35015 27226
rect 34719 27172 34775 27174
rect 34799 27172 34855 27174
rect 34879 27172 34935 27174
rect 34959 27172 35015 27174
rect 34719 26138 34775 26140
rect 34799 26138 34855 26140
rect 34879 26138 34935 26140
rect 34959 26138 35015 26140
rect 34719 26086 34765 26138
rect 34765 26086 34775 26138
rect 34799 26086 34829 26138
rect 34829 26086 34841 26138
rect 34841 26086 34855 26138
rect 34879 26086 34893 26138
rect 34893 26086 34905 26138
rect 34905 26086 34935 26138
rect 34959 26086 34969 26138
rect 34969 26086 35015 26138
rect 34719 26084 34775 26086
rect 34799 26084 34855 26086
rect 34879 26084 34935 26086
rect 34959 26084 35015 26086
rect 34719 25050 34775 25052
rect 34799 25050 34855 25052
rect 34879 25050 34935 25052
rect 34959 25050 35015 25052
rect 34719 24998 34765 25050
rect 34765 24998 34775 25050
rect 34799 24998 34829 25050
rect 34829 24998 34841 25050
rect 34841 24998 34855 25050
rect 34879 24998 34893 25050
rect 34893 24998 34905 25050
rect 34905 24998 34935 25050
rect 34959 24998 34969 25050
rect 34969 24998 35015 25050
rect 34719 24996 34775 24998
rect 34799 24996 34855 24998
rect 34879 24996 34935 24998
rect 34959 24996 35015 24998
rect 34719 23962 34775 23964
rect 34799 23962 34855 23964
rect 34879 23962 34935 23964
rect 34959 23962 35015 23964
rect 34719 23910 34765 23962
rect 34765 23910 34775 23962
rect 34799 23910 34829 23962
rect 34829 23910 34841 23962
rect 34841 23910 34855 23962
rect 34879 23910 34893 23962
rect 34893 23910 34905 23962
rect 34905 23910 34935 23962
rect 34959 23910 34969 23962
rect 34969 23910 35015 23962
rect 34719 23908 34775 23910
rect 34799 23908 34855 23910
rect 34879 23908 34935 23910
rect 34959 23908 35015 23910
rect 34719 22874 34775 22876
rect 34799 22874 34855 22876
rect 34879 22874 34935 22876
rect 34959 22874 35015 22876
rect 34719 22822 34765 22874
rect 34765 22822 34775 22874
rect 34799 22822 34829 22874
rect 34829 22822 34841 22874
rect 34841 22822 34855 22874
rect 34879 22822 34893 22874
rect 34893 22822 34905 22874
rect 34905 22822 34935 22874
rect 34959 22822 34969 22874
rect 34969 22822 35015 22874
rect 34719 22820 34775 22822
rect 34799 22820 34855 22822
rect 34879 22820 34935 22822
rect 34959 22820 35015 22822
rect 30499 20154 30555 20156
rect 30579 20154 30635 20156
rect 30659 20154 30715 20156
rect 30739 20154 30795 20156
rect 30499 20102 30545 20154
rect 30545 20102 30555 20154
rect 30579 20102 30609 20154
rect 30609 20102 30621 20154
rect 30621 20102 30635 20154
rect 30659 20102 30673 20154
rect 30673 20102 30685 20154
rect 30685 20102 30715 20154
rect 30739 20102 30749 20154
rect 30749 20102 30795 20154
rect 30499 20100 30555 20102
rect 30579 20100 30635 20102
rect 30659 20100 30715 20102
rect 30739 20100 30795 20102
rect 26278 17434 26334 17436
rect 26358 17434 26414 17436
rect 26438 17434 26494 17436
rect 26518 17434 26574 17436
rect 26278 17382 26324 17434
rect 26324 17382 26334 17434
rect 26358 17382 26388 17434
rect 26388 17382 26400 17434
rect 26400 17382 26414 17434
rect 26438 17382 26452 17434
rect 26452 17382 26464 17434
rect 26464 17382 26494 17434
rect 26518 17382 26528 17434
rect 26528 17382 26574 17434
rect 26278 17380 26334 17382
rect 26358 17380 26414 17382
rect 26438 17380 26494 17382
rect 26518 17380 26574 17382
rect 26278 16346 26334 16348
rect 26358 16346 26414 16348
rect 26438 16346 26494 16348
rect 26518 16346 26574 16348
rect 26278 16294 26324 16346
rect 26324 16294 26334 16346
rect 26358 16294 26388 16346
rect 26388 16294 26400 16346
rect 26400 16294 26414 16346
rect 26438 16294 26452 16346
rect 26452 16294 26464 16346
rect 26464 16294 26494 16346
rect 26518 16294 26528 16346
rect 26528 16294 26574 16346
rect 26278 16292 26334 16294
rect 26358 16292 26414 16294
rect 26438 16292 26494 16294
rect 26518 16292 26574 16294
rect 26278 15258 26334 15260
rect 26358 15258 26414 15260
rect 26438 15258 26494 15260
rect 26518 15258 26574 15260
rect 26278 15206 26324 15258
rect 26324 15206 26334 15258
rect 26358 15206 26388 15258
rect 26388 15206 26400 15258
rect 26400 15206 26414 15258
rect 26438 15206 26452 15258
rect 26452 15206 26464 15258
rect 26464 15206 26494 15258
rect 26518 15206 26528 15258
rect 26528 15206 26574 15258
rect 26278 15204 26334 15206
rect 26358 15204 26414 15206
rect 26438 15204 26494 15206
rect 26518 15204 26574 15206
rect 34886 21972 34888 21992
rect 34888 21972 34940 21992
rect 34940 21972 34942 21992
rect 34886 21936 34942 21972
rect 34719 21786 34775 21788
rect 34799 21786 34855 21788
rect 34879 21786 34935 21788
rect 34959 21786 35015 21788
rect 34719 21734 34765 21786
rect 34765 21734 34775 21786
rect 34799 21734 34829 21786
rect 34829 21734 34841 21786
rect 34841 21734 34855 21786
rect 34879 21734 34893 21786
rect 34893 21734 34905 21786
rect 34905 21734 34935 21786
rect 34959 21734 34969 21786
rect 34969 21734 35015 21786
rect 34719 21732 34775 21734
rect 34799 21732 34855 21734
rect 34879 21732 34935 21734
rect 34959 21732 35015 21734
rect 30499 19066 30555 19068
rect 30579 19066 30635 19068
rect 30659 19066 30715 19068
rect 30739 19066 30795 19068
rect 30499 19014 30545 19066
rect 30545 19014 30555 19066
rect 30579 19014 30609 19066
rect 30609 19014 30621 19066
rect 30621 19014 30635 19066
rect 30659 19014 30673 19066
rect 30673 19014 30685 19066
rect 30685 19014 30715 19066
rect 30739 19014 30749 19066
rect 30749 19014 30795 19066
rect 30499 19012 30555 19014
rect 30579 19012 30635 19014
rect 30659 19012 30715 19014
rect 30739 19012 30795 19014
rect 30499 17978 30555 17980
rect 30579 17978 30635 17980
rect 30659 17978 30715 17980
rect 30739 17978 30795 17980
rect 30499 17926 30545 17978
rect 30545 17926 30555 17978
rect 30579 17926 30609 17978
rect 30609 17926 30621 17978
rect 30621 17926 30635 17978
rect 30659 17926 30673 17978
rect 30673 17926 30685 17978
rect 30685 17926 30715 17978
rect 30739 17926 30749 17978
rect 30749 17926 30795 17978
rect 30499 17924 30555 17926
rect 30579 17924 30635 17926
rect 30659 17924 30715 17926
rect 30739 17924 30795 17926
rect 30499 16890 30555 16892
rect 30579 16890 30635 16892
rect 30659 16890 30715 16892
rect 30739 16890 30795 16892
rect 30499 16838 30545 16890
rect 30545 16838 30555 16890
rect 30579 16838 30609 16890
rect 30609 16838 30621 16890
rect 30621 16838 30635 16890
rect 30659 16838 30673 16890
rect 30673 16838 30685 16890
rect 30685 16838 30715 16890
rect 30739 16838 30749 16890
rect 30749 16838 30795 16890
rect 30499 16836 30555 16838
rect 30579 16836 30635 16838
rect 30659 16836 30715 16838
rect 30739 16836 30795 16838
rect 34719 20698 34775 20700
rect 34799 20698 34855 20700
rect 34879 20698 34935 20700
rect 34959 20698 35015 20700
rect 34719 20646 34765 20698
rect 34765 20646 34775 20698
rect 34799 20646 34829 20698
rect 34829 20646 34841 20698
rect 34841 20646 34855 20698
rect 34879 20646 34893 20698
rect 34893 20646 34905 20698
rect 34905 20646 34935 20698
rect 34959 20646 34969 20698
rect 34969 20646 35015 20698
rect 34719 20644 34775 20646
rect 34799 20644 34855 20646
rect 34879 20644 34935 20646
rect 34959 20644 35015 20646
rect 34719 19610 34775 19612
rect 34799 19610 34855 19612
rect 34879 19610 34935 19612
rect 34959 19610 35015 19612
rect 34719 19558 34765 19610
rect 34765 19558 34775 19610
rect 34799 19558 34829 19610
rect 34829 19558 34841 19610
rect 34841 19558 34855 19610
rect 34879 19558 34893 19610
rect 34893 19558 34905 19610
rect 34905 19558 34935 19610
rect 34959 19558 34969 19610
rect 34969 19558 35015 19610
rect 34719 19556 34775 19558
rect 34799 19556 34855 19558
rect 34879 19556 34935 19558
rect 34959 19556 35015 19558
rect 34719 18522 34775 18524
rect 34799 18522 34855 18524
rect 34879 18522 34935 18524
rect 34959 18522 35015 18524
rect 34719 18470 34765 18522
rect 34765 18470 34775 18522
rect 34799 18470 34829 18522
rect 34829 18470 34841 18522
rect 34841 18470 34855 18522
rect 34879 18470 34893 18522
rect 34893 18470 34905 18522
rect 34905 18470 34935 18522
rect 34959 18470 34969 18522
rect 34969 18470 35015 18522
rect 34719 18468 34775 18470
rect 34799 18468 34855 18470
rect 34879 18468 34935 18470
rect 34959 18468 35015 18470
rect 30499 15802 30555 15804
rect 30579 15802 30635 15804
rect 30659 15802 30715 15804
rect 30739 15802 30795 15804
rect 30499 15750 30545 15802
rect 30545 15750 30555 15802
rect 30579 15750 30609 15802
rect 30609 15750 30621 15802
rect 30621 15750 30635 15802
rect 30659 15750 30673 15802
rect 30673 15750 30685 15802
rect 30685 15750 30715 15802
rect 30739 15750 30749 15802
rect 30749 15750 30795 15802
rect 30499 15748 30555 15750
rect 30579 15748 30635 15750
rect 30659 15748 30715 15750
rect 30739 15748 30795 15750
rect 34719 17434 34775 17436
rect 34799 17434 34855 17436
rect 34879 17434 34935 17436
rect 34959 17434 35015 17436
rect 34719 17382 34765 17434
rect 34765 17382 34775 17434
rect 34799 17382 34829 17434
rect 34829 17382 34841 17434
rect 34841 17382 34855 17434
rect 34879 17382 34893 17434
rect 34893 17382 34905 17434
rect 34905 17382 34935 17434
rect 34959 17382 34969 17434
rect 34969 17382 35015 17434
rect 34719 17380 34775 17382
rect 34799 17380 34855 17382
rect 34879 17380 34935 17382
rect 34959 17380 35015 17382
rect 34719 16346 34775 16348
rect 34799 16346 34855 16348
rect 34879 16346 34935 16348
rect 34959 16346 35015 16348
rect 34719 16294 34765 16346
rect 34765 16294 34775 16346
rect 34799 16294 34829 16346
rect 34829 16294 34841 16346
rect 34841 16294 34855 16346
rect 34879 16294 34893 16346
rect 34893 16294 34905 16346
rect 34905 16294 34935 16346
rect 34959 16294 34969 16346
rect 34969 16294 35015 16346
rect 34719 16292 34775 16294
rect 34799 16292 34855 16294
rect 34879 16292 34935 16294
rect 34959 16292 35015 16294
rect 34719 15258 34775 15260
rect 34799 15258 34855 15260
rect 34879 15258 34935 15260
rect 34959 15258 35015 15260
rect 34719 15206 34765 15258
rect 34765 15206 34775 15258
rect 34799 15206 34829 15258
rect 34829 15206 34841 15258
rect 34841 15206 34855 15258
rect 34879 15206 34893 15258
rect 34893 15206 34905 15258
rect 34905 15206 34935 15258
rect 34959 15206 34969 15258
rect 34969 15206 35015 15258
rect 34719 15204 34775 15206
rect 34799 15204 34855 15206
rect 34879 15204 34935 15206
rect 34959 15204 35015 15206
rect 30499 14714 30555 14716
rect 30579 14714 30635 14716
rect 30659 14714 30715 14716
rect 30739 14714 30795 14716
rect 30499 14662 30545 14714
rect 30545 14662 30555 14714
rect 30579 14662 30609 14714
rect 30609 14662 30621 14714
rect 30621 14662 30635 14714
rect 30659 14662 30673 14714
rect 30673 14662 30685 14714
rect 30685 14662 30715 14714
rect 30739 14662 30749 14714
rect 30749 14662 30795 14714
rect 30499 14660 30555 14662
rect 30579 14660 30635 14662
rect 30659 14660 30715 14662
rect 30739 14660 30795 14662
rect 26278 14170 26334 14172
rect 26358 14170 26414 14172
rect 26438 14170 26494 14172
rect 26518 14170 26574 14172
rect 26278 14118 26324 14170
rect 26324 14118 26334 14170
rect 26358 14118 26388 14170
rect 26388 14118 26400 14170
rect 26400 14118 26414 14170
rect 26438 14118 26452 14170
rect 26452 14118 26464 14170
rect 26464 14118 26494 14170
rect 26518 14118 26528 14170
rect 26528 14118 26574 14170
rect 26278 14116 26334 14118
rect 26358 14116 26414 14118
rect 26438 14116 26494 14118
rect 26518 14116 26574 14118
rect 22058 13626 22114 13628
rect 22138 13626 22194 13628
rect 22218 13626 22274 13628
rect 22298 13626 22354 13628
rect 22058 13574 22104 13626
rect 22104 13574 22114 13626
rect 22138 13574 22168 13626
rect 22168 13574 22180 13626
rect 22180 13574 22194 13626
rect 22218 13574 22232 13626
rect 22232 13574 22244 13626
rect 22244 13574 22274 13626
rect 22298 13574 22308 13626
rect 22308 13574 22354 13626
rect 22058 13572 22114 13574
rect 22138 13572 22194 13574
rect 22218 13572 22274 13574
rect 22298 13572 22354 13574
rect 26278 13082 26334 13084
rect 26358 13082 26414 13084
rect 26438 13082 26494 13084
rect 26518 13082 26574 13084
rect 26278 13030 26324 13082
rect 26324 13030 26334 13082
rect 26358 13030 26388 13082
rect 26388 13030 26400 13082
rect 26400 13030 26414 13082
rect 26438 13030 26452 13082
rect 26452 13030 26464 13082
rect 26464 13030 26494 13082
rect 26518 13030 26528 13082
rect 26528 13030 26574 13082
rect 26278 13028 26334 13030
rect 26358 13028 26414 13030
rect 26438 13028 26494 13030
rect 26518 13028 26574 13030
rect 22058 12538 22114 12540
rect 22138 12538 22194 12540
rect 22218 12538 22274 12540
rect 22298 12538 22354 12540
rect 22058 12486 22104 12538
rect 22104 12486 22114 12538
rect 22138 12486 22168 12538
rect 22168 12486 22180 12538
rect 22180 12486 22194 12538
rect 22218 12486 22232 12538
rect 22232 12486 22244 12538
rect 22244 12486 22274 12538
rect 22298 12486 22308 12538
rect 22308 12486 22354 12538
rect 22058 12484 22114 12486
rect 22138 12484 22194 12486
rect 22218 12484 22274 12486
rect 22298 12484 22354 12486
rect 26278 11994 26334 11996
rect 26358 11994 26414 11996
rect 26438 11994 26494 11996
rect 26518 11994 26574 11996
rect 26278 11942 26324 11994
rect 26324 11942 26334 11994
rect 26358 11942 26388 11994
rect 26388 11942 26400 11994
rect 26400 11942 26414 11994
rect 26438 11942 26452 11994
rect 26452 11942 26464 11994
rect 26464 11942 26494 11994
rect 26518 11942 26528 11994
rect 26528 11942 26574 11994
rect 26278 11940 26334 11942
rect 26358 11940 26414 11942
rect 26438 11940 26494 11942
rect 26518 11940 26574 11942
rect 22058 11450 22114 11452
rect 22138 11450 22194 11452
rect 22218 11450 22274 11452
rect 22298 11450 22354 11452
rect 22058 11398 22104 11450
rect 22104 11398 22114 11450
rect 22138 11398 22168 11450
rect 22168 11398 22180 11450
rect 22180 11398 22194 11450
rect 22218 11398 22232 11450
rect 22232 11398 22244 11450
rect 22244 11398 22274 11450
rect 22298 11398 22308 11450
rect 22308 11398 22354 11450
rect 22058 11396 22114 11398
rect 22138 11396 22194 11398
rect 22218 11396 22274 11398
rect 22298 11396 22354 11398
rect 26278 10906 26334 10908
rect 26358 10906 26414 10908
rect 26438 10906 26494 10908
rect 26518 10906 26574 10908
rect 26278 10854 26324 10906
rect 26324 10854 26334 10906
rect 26358 10854 26388 10906
rect 26388 10854 26400 10906
rect 26400 10854 26414 10906
rect 26438 10854 26452 10906
rect 26452 10854 26464 10906
rect 26464 10854 26494 10906
rect 26518 10854 26528 10906
rect 26528 10854 26574 10906
rect 26278 10852 26334 10854
rect 26358 10852 26414 10854
rect 26438 10852 26494 10854
rect 26518 10852 26574 10854
rect 22058 10362 22114 10364
rect 22138 10362 22194 10364
rect 22218 10362 22274 10364
rect 22298 10362 22354 10364
rect 22058 10310 22104 10362
rect 22104 10310 22114 10362
rect 22138 10310 22168 10362
rect 22168 10310 22180 10362
rect 22180 10310 22194 10362
rect 22218 10310 22232 10362
rect 22232 10310 22244 10362
rect 22244 10310 22274 10362
rect 22298 10310 22308 10362
rect 22308 10310 22354 10362
rect 22058 10308 22114 10310
rect 22138 10308 22194 10310
rect 22218 10308 22274 10310
rect 22298 10308 22354 10310
rect 26278 9818 26334 9820
rect 26358 9818 26414 9820
rect 26438 9818 26494 9820
rect 26518 9818 26574 9820
rect 26278 9766 26324 9818
rect 26324 9766 26334 9818
rect 26358 9766 26388 9818
rect 26388 9766 26400 9818
rect 26400 9766 26414 9818
rect 26438 9766 26452 9818
rect 26452 9766 26464 9818
rect 26464 9766 26494 9818
rect 26518 9766 26528 9818
rect 26528 9766 26574 9818
rect 26278 9764 26334 9766
rect 26358 9764 26414 9766
rect 26438 9764 26494 9766
rect 26518 9764 26574 9766
rect 22058 9274 22114 9276
rect 22138 9274 22194 9276
rect 22218 9274 22274 9276
rect 22298 9274 22354 9276
rect 22058 9222 22104 9274
rect 22104 9222 22114 9274
rect 22138 9222 22168 9274
rect 22168 9222 22180 9274
rect 22180 9222 22194 9274
rect 22218 9222 22232 9274
rect 22232 9222 22244 9274
rect 22244 9222 22274 9274
rect 22298 9222 22308 9274
rect 22308 9222 22354 9274
rect 22058 9220 22114 9222
rect 22138 9220 22194 9222
rect 22218 9220 22274 9222
rect 22298 9220 22354 9222
rect 26278 8730 26334 8732
rect 26358 8730 26414 8732
rect 26438 8730 26494 8732
rect 26518 8730 26574 8732
rect 26278 8678 26324 8730
rect 26324 8678 26334 8730
rect 26358 8678 26388 8730
rect 26388 8678 26400 8730
rect 26400 8678 26414 8730
rect 26438 8678 26452 8730
rect 26452 8678 26464 8730
rect 26464 8678 26494 8730
rect 26518 8678 26528 8730
rect 26528 8678 26574 8730
rect 26278 8676 26334 8678
rect 26358 8676 26414 8678
rect 26438 8676 26494 8678
rect 26518 8676 26574 8678
rect 22058 8186 22114 8188
rect 22138 8186 22194 8188
rect 22218 8186 22274 8188
rect 22298 8186 22354 8188
rect 22058 8134 22104 8186
rect 22104 8134 22114 8186
rect 22138 8134 22168 8186
rect 22168 8134 22180 8186
rect 22180 8134 22194 8186
rect 22218 8134 22232 8186
rect 22232 8134 22244 8186
rect 22244 8134 22274 8186
rect 22298 8134 22308 8186
rect 22308 8134 22354 8186
rect 22058 8132 22114 8134
rect 22138 8132 22194 8134
rect 22218 8132 22274 8134
rect 22298 8132 22354 8134
rect 26278 7642 26334 7644
rect 26358 7642 26414 7644
rect 26438 7642 26494 7644
rect 26518 7642 26574 7644
rect 26278 7590 26324 7642
rect 26324 7590 26334 7642
rect 26358 7590 26388 7642
rect 26388 7590 26400 7642
rect 26400 7590 26414 7642
rect 26438 7590 26452 7642
rect 26452 7590 26464 7642
rect 26464 7590 26494 7642
rect 26518 7590 26528 7642
rect 26528 7590 26574 7642
rect 26278 7588 26334 7590
rect 26358 7588 26414 7590
rect 26438 7588 26494 7590
rect 26518 7588 26574 7590
rect 22058 7098 22114 7100
rect 22138 7098 22194 7100
rect 22218 7098 22274 7100
rect 22298 7098 22354 7100
rect 22058 7046 22104 7098
rect 22104 7046 22114 7098
rect 22138 7046 22168 7098
rect 22168 7046 22180 7098
rect 22180 7046 22194 7098
rect 22218 7046 22232 7098
rect 22232 7046 22244 7098
rect 22244 7046 22274 7098
rect 22298 7046 22308 7098
rect 22308 7046 22354 7098
rect 22058 7044 22114 7046
rect 22138 7044 22194 7046
rect 22218 7044 22274 7046
rect 22298 7044 22354 7046
rect 9396 6554 9452 6556
rect 9476 6554 9532 6556
rect 9556 6554 9612 6556
rect 9636 6554 9692 6556
rect 9396 6502 9442 6554
rect 9442 6502 9452 6554
rect 9476 6502 9506 6554
rect 9506 6502 9518 6554
rect 9518 6502 9532 6554
rect 9556 6502 9570 6554
rect 9570 6502 9582 6554
rect 9582 6502 9612 6554
rect 9636 6502 9646 6554
rect 9646 6502 9692 6554
rect 9396 6500 9452 6502
rect 9476 6500 9532 6502
rect 9556 6500 9612 6502
rect 9636 6500 9692 6502
rect 17837 6554 17893 6556
rect 17917 6554 17973 6556
rect 17997 6554 18053 6556
rect 18077 6554 18133 6556
rect 17837 6502 17883 6554
rect 17883 6502 17893 6554
rect 17917 6502 17947 6554
rect 17947 6502 17959 6554
rect 17959 6502 17973 6554
rect 17997 6502 18011 6554
rect 18011 6502 18023 6554
rect 18023 6502 18053 6554
rect 18077 6502 18087 6554
rect 18087 6502 18133 6554
rect 17837 6500 17893 6502
rect 17917 6500 17973 6502
rect 17997 6500 18053 6502
rect 18077 6500 18133 6502
rect 5176 6010 5232 6012
rect 5256 6010 5312 6012
rect 5336 6010 5392 6012
rect 5416 6010 5472 6012
rect 5176 5958 5222 6010
rect 5222 5958 5232 6010
rect 5256 5958 5286 6010
rect 5286 5958 5298 6010
rect 5298 5958 5312 6010
rect 5336 5958 5350 6010
rect 5350 5958 5362 6010
rect 5362 5958 5392 6010
rect 5416 5958 5426 6010
rect 5426 5958 5472 6010
rect 5176 5956 5232 5958
rect 5256 5956 5312 5958
rect 5336 5956 5392 5958
rect 5416 5956 5472 5958
rect 13617 6010 13673 6012
rect 13697 6010 13753 6012
rect 13777 6010 13833 6012
rect 13857 6010 13913 6012
rect 13617 5958 13663 6010
rect 13663 5958 13673 6010
rect 13697 5958 13727 6010
rect 13727 5958 13739 6010
rect 13739 5958 13753 6010
rect 13777 5958 13791 6010
rect 13791 5958 13803 6010
rect 13803 5958 13833 6010
rect 13857 5958 13867 6010
rect 13867 5958 13913 6010
rect 13617 5956 13673 5958
rect 13697 5956 13753 5958
rect 13777 5956 13833 5958
rect 13857 5956 13913 5958
rect 9396 5466 9452 5468
rect 9476 5466 9532 5468
rect 9556 5466 9612 5468
rect 9636 5466 9692 5468
rect 9396 5414 9442 5466
rect 9442 5414 9452 5466
rect 9476 5414 9506 5466
rect 9506 5414 9518 5466
rect 9518 5414 9532 5466
rect 9556 5414 9570 5466
rect 9570 5414 9582 5466
rect 9582 5414 9612 5466
rect 9636 5414 9646 5466
rect 9646 5414 9692 5466
rect 9396 5412 9452 5414
rect 9476 5412 9532 5414
rect 9556 5412 9612 5414
rect 9636 5412 9692 5414
rect 17837 5466 17893 5468
rect 17917 5466 17973 5468
rect 17997 5466 18053 5468
rect 18077 5466 18133 5468
rect 17837 5414 17883 5466
rect 17883 5414 17893 5466
rect 17917 5414 17947 5466
rect 17947 5414 17959 5466
rect 17959 5414 17973 5466
rect 17997 5414 18011 5466
rect 18011 5414 18023 5466
rect 18023 5414 18053 5466
rect 18077 5414 18087 5466
rect 18087 5414 18133 5466
rect 17837 5412 17893 5414
rect 17917 5412 17973 5414
rect 17997 5412 18053 5414
rect 18077 5412 18133 5414
rect 5176 4922 5232 4924
rect 5256 4922 5312 4924
rect 5336 4922 5392 4924
rect 5416 4922 5472 4924
rect 5176 4870 5222 4922
rect 5222 4870 5232 4922
rect 5256 4870 5286 4922
rect 5286 4870 5298 4922
rect 5298 4870 5312 4922
rect 5336 4870 5350 4922
rect 5350 4870 5362 4922
rect 5362 4870 5392 4922
rect 5416 4870 5426 4922
rect 5426 4870 5472 4922
rect 5176 4868 5232 4870
rect 5256 4868 5312 4870
rect 5336 4868 5392 4870
rect 5416 4868 5472 4870
rect 13617 4922 13673 4924
rect 13697 4922 13753 4924
rect 13777 4922 13833 4924
rect 13857 4922 13913 4924
rect 13617 4870 13663 4922
rect 13663 4870 13673 4922
rect 13697 4870 13727 4922
rect 13727 4870 13739 4922
rect 13739 4870 13753 4922
rect 13777 4870 13791 4922
rect 13791 4870 13803 4922
rect 13803 4870 13833 4922
rect 13857 4870 13867 4922
rect 13867 4870 13913 4922
rect 13617 4868 13673 4870
rect 13697 4868 13753 4870
rect 13777 4868 13833 4870
rect 13857 4868 13913 4870
rect 9396 4378 9452 4380
rect 9476 4378 9532 4380
rect 9556 4378 9612 4380
rect 9636 4378 9692 4380
rect 9396 4326 9442 4378
rect 9442 4326 9452 4378
rect 9476 4326 9506 4378
rect 9506 4326 9518 4378
rect 9518 4326 9532 4378
rect 9556 4326 9570 4378
rect 9570 4326 9582 4378
rect 9582 4326 9612 4378
rect 9636 4326 9646 4378
rect 9646 4326 9692 4378
rect 9396 4324 9452 4326
rect 9476 4324 9532 4326
rect 9556 4324 9612 4326
rect 9636 4324 9692 4326
rect 17837 4378 17893 4380
rect 17917 4378 17973 4380
rect 17997 4378 18053 4380
rect 18077 4378 18133 4380
rect 17837 4326 17883 4378
rect 17883 4326 17893 4378
rect 17917 4326 17947 4378
rect 17947 4326 17959 4378
rect 17959 4326 17973 4378
rect 17997 4326 18011 4378
rect 18011 4326 18023 4378
rect 18023 4326 18053 4378
rect 18077 4326 18087 4378
rect 18087 4326 18133 4378
rect 17837 4324 17893 4326
rect 17917 4324 17973 4326
rect 17997 4324 18053 4326
rect 18077 4324 18133 4326
rect 5176 3834 5232 3836
rect 5256 3834 5312 3836
rect 5336 3834 5392 3836
rect 5416 3834 5472 3836
rect 5176 3782 5222 3834
rect 5222 3782 5232 3834
rect 5256 3782 5286 3834
rect 5286 3782 5298 3834
rect 5298 3782 5312 3834
rect 5336 3782 5350 3834
rect 5350 3782 5362 3834
rect 5362 3782 5392 3834
rect 5416 3782 5426 3834
rect 5426 3782 5472 3834
rect 5176 3780 5232 3782
rect 5256 3780 5312 3782
rect 5336 3780 5392 3782
rect 5416 3780 5472 3782
rect 13617 3834 13673 3836
rect 13697 3834 13753 3836
rect 13777 3834 13833 3836
rect 13857 3834 13913 3836
rect 13617 3782 13663 3834
rect 13663 3782 13673 3834
rect 13697 3782 13727 3834
rect 13727 3782 13739 3834
rect 13739 3782 13753 3834
rect 13777 3782 13791 3834
rect 13791 3782 13803 3834
rect 13803 3782 13833 3834
rect 13857 3782 13867 3834
rect 13867 3782 13913 3834
rect 13617 3780 13673 3782
rect 13697 3780 13753 3782
rect 13777 3780 13833 3782
rect 13857 3780 13913 3782
rect 9396 3290 9452 3292
rect 9476 3290 9532 3292
rect 9556 3290 9612 3292
rect 9636 3290 9692 3292
rect 9396 3238 9442 3290
rect 9442 3238 9452 3290
rect 9476 3238 9506 3290
rect 9506 3238 9518 3290
rect 9518 3238 9532 3290
rect 9556 3238 9570 3290
rect 9570 3238 9582 3290
rect 9582 3238 9612 3290
rect 9636 3238 9646 3290
rect 9646 3238 9692 3290
rect 9396 3236 9452 3238
rect 9476 3236 9532 3238
rect 9556 3236 9612 3238
rect 9636 3236 9692 3238
rect 17837 3290 17893 3292
rect 17917 3290 17973 3292
rect 17997 3290 18053 3292
rect 18077 3290 18133 3292
rect 17837 3238 17883 3290
rect 17883 3238 17893 3290
rect 17917 3238 17947 3290
rect 17947 3238 17959 3290
rect 17959 3238 17973 3290
rect 17997 3238 18011 3290
rect 18011 3238 18023 3290
rect 18023 3238 18053 3290
rect 18077 3238 18087 3290
rect 18087 3238 18133 3290
rect 17837 3236 17893 3238
rect 17917 3236 17973 3238
rect 17997 3236 18053 3238
rect 18077 3236 18133 3238
rect 5176 2746 5232 2748
rect 5256 2746 5312 2748
rect 5336 2746 5392 2748
rect 5416 2746 5472 2748
rect 5176 2694 5222 2746
rect 5222 2694 5232 2746
rect 5256 2694 5286 2746
rect 5286 2694 5298 2746
rect 5298 2694 5312 2746
rect 5336 2694 5350 2746
rect 5350 2694 5362 2746
rect 5362 2694 5392 2746
rect 5416 2694 5426 2746
rect 5426 2694 5472 2746
rect 5176 2692 5232 2694
rect 5256 2692 5312 2694
rect 5336 2692 5392 2694
rect 5416 2692 5472 2694
rect 13617 2746 13673 2748
rect 13697 2746 13753 2748
rect 13777 2746 13833 2748
rect 13857 2746 13913 2748
rect 13617 2694 13663 2746
rect 13663 2694 13673 2746
rect 13697 2694 13727 2746
rect 13727 2694 13739 2746
rect 13739 2694 13753 2746
rect 13777 2694 13791 2746
rect 13791 2694 13803 2746
rect 13803 2694 13833 2746
rect 13857 2694 13867 2746
rect 13867 2694 13913 2746
rect 13617 2692 13673 2694
rect 13697 2692 13753 2694
rect 13777 2692 13833 2694
rect 13857 2692 13913 2694
rect 26278 6554 26334 6556
rect 26358 6554 26414 6556
rect 26438 6554 26494 6556
rect 26518 6554 26574 6556
rect 26278 6502 26324 6554
rect 26324 6502 26334 6554
rect 26358 6502 26388 6554
rect 26388 6502 26400 6554
rect 26400 6502 26414 6554
rect 26438 6502 26452 6554
rect 26452 6502 26464 6554
rect 26464 6502 26494 6554
rect 26518 6502 26528 6554
rect 26528 6502 26574 6554
rect 26278 6500 26334 6502
rect 26358 6500 26414 6502
rect 26438 6500 26494 6502
rect 26518 6500 26574 6502
rect 22058 6010 22114 6012
rect 22138 6010 22194 6012
rect 22218 6010 22274 6012
rect 22298 6010 22354 6012
rect 22058 5958 22104 6010
rect 22104 5958 22114 6010
rect 22138 5958 22168 6010
rect 22168 5958 22180 6010
rect 22180 5958 22194 6010
rect 22218 5958 22232 6010
rect 22232 5958 22244 6010
rect 22244 5958 22274 6010
rect 22298 5958 22308 6010
rect 22308 5958 22354 6010
rect 22058 5956 22114 5958
rect 22138 5956 22194 5958
rect 22218 5956 22274 5958
rect 22298 5956 22354 5958
rect 26278 5466 26334 5468
rect 26358 5466 26414 5468
rect 26438 5466 26494 5468
rect 26518 5466 26574 5468
rect 26278 5414 26324 5466
rect 26324 5414 26334 5466
rect 26358 5414 26388 5466
rect 26388 5414 26400 5466
rect 26400 5414 26414 5466
rect 26438 5414 26452 5466
rect 26452 5414 26464 5466
rect 26464 5414 26494 5466
rect 26518 5414 26528 5466
rect 26528 5414 26574 5466
rect 26278 5412 26334 5414
rect 26358 5412 26414 5414
rect 26438 5412 26494 5414
rect 26518 5412 26574 5414
rect 22058 4922 22114 4924
rect 22138 4922 22194 4924
rect 22218 4922 22274 4924
rect 22298 4922 22354 4924
rect 22058 4870 22104 4922
rect 22104 4870 22114 4922
rect 22138 4870 22168 4922
rect 22168 4870 22180 4922
rect 22180 4870 22194 4922
rect 22218 4870 22232 4922
rect 22232 4870 22244 4922
rect 22244 4870 22274 4922
rect 22298 4870 22308 4922
rect 22308 4870 22354 4922
rect 22058 4868 22114 4870
rect 22138 4868 22194 4870
rect 22218 4868 22274 4870
rect 22298 4868 22354 4870
rect 26278 4378 26334 4380
rect 26358 4378 26414 4380
rect 26438 4378 26494 4380
rect 26518 4378 26574 4380
rect 26278 4326 26324 4378
rect 26324 4326 26334 4378
rect 26358 4326 26388 4378
rect 26388 4326 26400 4378
rect 26400 4326 26414 4378
rect 26438 4326 26452 4378
rect 26452 4326 26464 4378
rect 26464 4326 26494 4378
rect 26518 4326 26528 4378
rect 26528 4326 26574 4378
rect 26278 4324 26334 4326
rect 26358 4324 26414 4326
rect 26438 4324 26494 4326
rect 26518 4324 26574 4326
rect 22058 3834 22114 3836
rect 22138 3834 22194 3836
rect 22218 3834 22274 3836
rect 22298 3834 22354 3836
rect 22058 3782 22104 3834
rect 22104 3782 22114 3834
rect 22138 3782 22168 3834
rect 22168 3782 22180 3834
rect 22180 3782 22194 3834
rect 22218 3782 22232 3834
rect 22232 3782 22244 3834
rect 22244 3782 22274 3834
rect 22298 3782 22308 3834
rect 22308 3782 22354 3834
rect 22058 3780 22114 3782
rect 22138 3780 22194 3782
rect 22218 3780 22274 3782
rect 22298 3780 22354 3782
rect 26278 3290 26334 3292
rect 26358 3290 26414 3292
rect 26438 3290 26494 3292
rect 26518 3290 26574 3292
rect 26278 3238 26324 3290
rect 26324 3238 26334 3290
rect 26358 3238 26388 3290
rect 26388 3238 26400 3290
rect 26400 3238 26414 3290
rect 26438 3238 26452 3290
rect 26452 3238 26464 3290
rect 26464 3238 26494 3290
rect 26518 3238 26528 3290
rect 26528 3238 26574 3290
rect 26278 3236 26334 3238
rect 26358 3236 26414 3238
rect 26438 3236 26494 3238
rect 26518 3236 26574 3238
rect 22058 2746 22114 2748
rect 22138 2746 22194 2748
rect 22218 2746 22274 2748
rect 22298 2746 22354 2748
rect 22058 2694 22104 2746
rect 22104 2694 22114 2746
rect 22138 2694 22168 2746
rect 22168 2694 22180 2746
rect 22180 2694 22194 2746
rect 22218 2694 22232 2746
rect 22232 2694 22244 2746
rect 22244 2694 22274 2746
rect 22298 2694 22308 2746
rect 22308 2694 22354 2746
rect 22058 2692 22114 2694
rect 22138 2692 22194 2694
rect 22218 2692 22274 2694
rect 22298 2692 22354 2694
rect 30499 13626 30555 13628
rect 30579 13626 30635 13628
rect 30659 13626 30715 13628
rect 30739 13626 30795 13628
rect 30499 13574 30545 13626
rect 30545 13574 30555 13626
rect 30579 13574 30609 13626
rect 30609 13574 30621 13626
rect 30621 13574 30635 13626
rect 30659 13574 30673 13626
rect 30673 13574 30685 13626
rect 30685 13574 30715 13626
rect 30739 13574 30749 13626
rect 30749 13574 30795 13626
rect 30499 13572 30555 13574
rect 30579 13572 30635 13574
rect 30659 13572 30715 13574
rect 30739 13572 30795 13574
rect 30499 12538 30555 12540
rect 30579 12538 30635 12540
rect 30659 12538 30715 12540
rect 30739 12538 30795 12540
rect 30499 12486 30545 12538
rect 30545 12486 30555 12538
rect 30579 12486 30609 12538
rect 30609 12486 30621 12538
rect 30621 12486 30635 12538
rect 30659 12486 30673 12538
rect 30673 12486 30685 12538
rect 30685 12486 30715 12538
rect 30739 12486 30749 12538
rect 30749 12486 30795 12538
rect 30499 12484 30555 12486
rect 30579 12484 30635 12486
rect 30659 12484 30715 12486
rect 30739 12484 30795 12486
rect 30499 11450 30555 11452
rect 30579 11450 30635 11452
rect 30659 11450 30715 11452
rect 30739 11450 30795 11452
rect 30499 11398 30545 11450
rect 30545 11398 30555 11450
rect 30579 11398 30609 11450
rect 30609 11398 30621 11450
rect 30621 11398 30635 11450
rect 30659 11398 30673 11450
rect 30673 11398 30685 11450
rect 30685 11398 30715 11450
rect 30739 11398 30749 11450
rect 30749 11398 30795 11450
rect 30499 11396 30555 11398
rect 30579 11396 30635 11398
rect 30659 11396 30715 11398
rect 30739 11396 30795 11398
rect 30499 10362 30555 10364
rect 30579 10362 30635 10364
rect 30659 10362 30715 10364
rect 30739 10362 30795 10364
rect 30499 10310 30545 10362
rect 30545 10310 30555 10362
rect 30579 10310 30609 10362
rect 30609 10310 30621 10362
rect 30621 10310 30635 10362
rect 30659 10310 30673 10362
rect 30673 10310 30685 10362
rect 30685 10310 30715 10362
rect 30739 10310 30749 10362
rect 30749 10310 30795 10362
rect 30499 10308 30555 10310
rect 30579 10308 30635 10310
rect 30659 10308 30715 10310
rect 30739 10308 30795 10310
rect 30499 9274 30555 9276
rect 30579 9274 30635 9276
rect 30659 9274 30715 9276
rect 30739 9274 30795 9276
rect 30499 9222 30545 9274
rect 30545 9222 30555 9274
rect 30579 9222 30609 9274
rect 30609 9222 30621 9274
rect 30621 9222 30635 9274
rect 30659 9222 30673 9274
rect 30673 9222 30685 9274
rect 30685 9222 30715 9274
rect 30739 9222 30749 9274
rect 30749 9222 30795 9274
rect 30499 9220 30555 9222
rect 30579 9220 30635 9222
rect 30659 9220 30715 9222
rect 30739 9220 30795 9222
rect 30499 8186 30555 8188
rect 30579 8186 30635 8188
rect 30659 8186 30715 8188
rect 30739 8186 30795 8188
rect 30499 8134 30545 8186
rect 30545 8134 30555 8186
rect 30579 8134 30609 8186
rect 30609 8134 30621 8186
rect 30621 8134 30635 8186
rect 30659 8134 30673 8186
rect 30673 8134 30685 8186
rect 30685 8134 30715 8186
rect 30739 8134 30749 8186
rect 30749 8134 30795 8186
rect 30499 8132 30555 8134
rect 30579 8132 30635 8134
rect 30659 8132 30715 8134
rect 30739 8132 30795 8134
rect 30499 7098 30555 7100
rect 30579 7098 30635 7100
rect 30659 7098 30715 7100
rect 30739 7098 30795 7100
rect 30499 7046 30545 7098
rect 30545 7046 30555 7098
rect 30579 7046 30609 7098
rect 30609 7046 30621 7098
rect 30621 7046 30635 7098
rect 30659 7046 30673 7098
rect 30673 7046 30685 7098
rect 30685 7046 30715 7098
rect 30739 7046 30749 7098
rect 30749 7046 30795 7098
rect 30499 7044 30555 7046
rect 30579 7044 30635 7046
rect 30659 7044 30715 7046
rect 30739 7044 30795 7046
rect 30499 6010 30555 6012
rect 30579 6010 30635 6012
rect 30659 6010 30715 6012
rect 30739 6010 30795 6012
rect 30499 5958 30545 6010
rect 30545 5958 30555 6010
rect 30579 5958 30609 6010
rect 30609 5958 30621 6010
rect 30621 5958 30635 6010
rect 30659 5958 30673 6010
rect 30673 5958 30685 6010
rect 30685 5958 30715 6010
rect 30739 5958 30749 6010
rect 30749 5958 30795 6010
rect 30499 5956 30555 5958
rect 30579 5956 30635 5958
rect 30659 5956 30715 5958
rect 30739 5956 30795 5958
rect 30499 4922 30555 4924
rect 30579 4922 30635 4924
rect 30659 4922 30715 4924
rect 30739 4922 30795 4924
rect 30499 4870 30545 4922
rect 30545 4870 30555 4922
rect 30579 4870 30609 4922
rect 30609 4870 30621 4922
rect 30621 4870 30635 4922
rect 30659 4870 30673 4922
rect 30673 4870 30685 4922
rect 30685 4870 30715 4922
rect 30739 4870 30749 4922
rect 30749 4870 30795 4922
rect 30499 4868 30555 4870
rect 30579 4868 30635 4870
rect 30659 4868 30715 4870
rect 30739 4868 30795 4870
rect 30499 3834 30555 3836
rect 30579 3834 30635 3836
rect 30659 3834 30715 3836
rect 30739 3834 30795 3836
rect 30499 3782 30545 3834
rect 30545 3782 30555 3834
rect 30579 3782 30609 3834
rect 30609 3782 30621 3834
rect 30621 3782 30635 3834
rect 30659 3782 30673 3834
rect 30673 3782 30685 3834
rect 30685 3782 30715 3834
rect 30739 3782 30749 3834
rect 30749 3782 30795 3834
rect 30499 3780 30555 3782
rect 30579 3780 30635 3782
rect 30659 3780 30715 3782
rect 30739 3780 30795 3782
rect 30499 2746 30555 2748
rect 30579 2746 30635 2748
rect 30659 2746 30715 2748
rect 30739 2746 30795 2748
rect 30499 2694 30545 2746
rect 30545 2694 30555 2746
rect 30579 2694 30609 2746
rect 30609 2694 30621 2746
rect 30621 2694 30635 2746
rect 30659 2694 30673 2746
rect 30673 2694 30685 2746
rect 30685 2694 30715 2746
rect 30739 2694 30749 2746
rect 30749 2694 30795 2746
rect 30499 2692 30555 2694
rect 30579 2692 30635 2694
rect 30659 2692 30715 2694
rect 30739 2692 30795 2694
rect 34719 14170 34775 14172
rect 34799 14170 34855 14172
rect 34879 14170 34935 14172
rect 34959 14170 35015 14172
rect 34719 14118 34765 14170
rect 34765 14118 34775 14170
rect 34799 14118 34829 14170
rect 34829 14118 34841 14170
rect 34841 14118 34855 14170
rect 34879 14118 34893 14170
rect 34893 14118 34905 14170
rect 34905 14118 34935 14170
rect 34959 14118 34969 14170
rect 34969 14118 35015 14170
rect 34719 14116 34775 14118
rect 34799 14116 34855 14118
rect 34879 14116 34935 14118
rect 34959 14116 35015 14118
rect 34719 13082 34775 13084
rect 34799 13082 34855 13084
rect 34879 13082 34935 13084
rect 34959 13082 35015 13084
rect 34719 13030 34765 13082
rect 34765 13030 34775 13082
rect 34799 13030 34829 13082
rect 34829 13030 34841 13082
rect 34841 13030 34855 13082
rect 34879 13030 34893 13082
rect 34893 13030 34905 13082
rect 34905 13030 34935 13082
rect 34959 13030 34969 13082
rect 34969 13030 35015 13082
rect 34719 13028 34775 13030
rect 34799 13028 34855 13030
rect 34879 13028 34935 13030
rect 34959 13028 35015 13030
rect 34719 11994 34775 11996
rect 34799 11994 34855 11996
rect 34879 11994 34935 11996
rect 34959 11994 35015 11996
rect 34719 11942 34765 11994
rect 34765 11942 34775 11994
rect 34799 11942 34829 11994
rect 34829 11942 34841 11994
rect 34841 11942 34855 11994
rect 34879 11942 34893 11994
rect 34893 11942 34905 11994
rect 34905 11942 34935 11994
rect 34959 11942 34969 11994
rect 34969 11942 35015 11994
rect 34719 11940 34775 11942
rect 34799 11940 34855 11942
rect 34879 11940 34935 11942
rect 34959 11940 35015 11942
rect 34518 11620 34574 11656
rect 34518 11600 34520 11620
rect 34520 11600 34572 11620
rect 34572 11600 34574 11620
rect 34719 10906 34775 10908
rect 34799 10906 34855 10908
rect 34879 10906 34935 10908
rect 34959 10906 35015 10908
rect 34719 10854 34765 10906
rect 34765 10854 34775 10906
rect 34799 10854 34829 10906
rect 34829 10854 34841 10906
rect 34841 10854 34855 10906
rect 34879 10854 34893 10906
rect 34893 10854 34905 10906
rect 34905 10854 34935 10906
rect 34959 10854 34969 10906
rect 34969 10854 35015 10906
rect 34719 10852 34775 10854
rect 34799 10852 34855 10854
rect 34879 10852 34935 10854
rect 34959 10852 35015 10854
rect 34719 9818 34775 9820
rect 34799 9818 34855 9820
rect 34879 9818 34935 9820
rect 34959 9818 35015 9820
rect 34719 9766 34765 9818
rect 34765 9766 34775 9818
rect 34799 9766 34829 9818
rect 34829 9766 34841 9818
rect 34841 9766 34855 9818
rect 34879 9766 34893 9818
rect 34893 9766 34905 9818
rect 34905 9766 34935 9818
rect 34959 9766 34969 9818
rect 34969 9766 35015 9818
rect 34719 9764 34775 9766
rect 34799 9764 34855 9766
rect 34879 9764 34935 9766
rect 34959 9764 35015 9766
rect 34719 8730 34775 8732
rect 34799 8730 34855 8732
rect 34879 8730 34935 8732
rect 34959 8730 35015 8732
rect 34719 8678 34765 8730
rect 34765 8678 34775 8730
rect 34799 8678 34829 8730
rect 34829 8678 34841 8730
rect 34841 8678 34855 8730
rect 34879 8678 34893 8730
rect 34893 8678 34905 8730
rect 34905 8678 34935 8730
rect 34959 8678 34969 8730
rect 34969 8678 35015 8730
rect 34719 8676 34775 8678
rect 34799 8676 34855 8678
rect 34879 8676 34935 8678
rect 34959 8676 35015 8678
rect 34719 7642 34775 7644
rect 34799 7642 34855 7644
rect 34879 7642 34935 7644
rect 34959 7642 35015 7644
rect 34719 7590 34765 7642
rect 34765 7590 34775 7642
rect 34799 7590 34829 7642
rect 34829 7590 34841 7642
rect 34841 7590 34855 7642
rect 34879 7590 34893 7642
rect 34893 7590 34905 7642
rect 34905 7590 34935 7642
rect 34959 7590 34969 7642
rect 34969 7590 35015 7642
rect 34719 7588 34775 7590
rect 34799 7588 34855 7590
rect 34879 7588 34935 7590
rect 34959 7588 35015 7590
rect 34719 6554 34775 6556
rect 34799 6554 34855 6556
rect 34879 6554 34935 6556
rect 34959 6554 35015 6556
rect 34719 6502 34765 6554
rect 34765 6502 34775 6554
rect 34799 6502 34829 6554
rect 34829 6502 34841 6554
rect 34841 6502 34855 6554
rect 34879 6502 34893 6554
rect 34893 6502 34905 6554
rect 34905 6502 34935 6554
rect 34959 6502 34969 6554
rect 34969 6502 35015 6554
rect 34719 6500 34775 6502
rect 34799 6500 34855 6502
rect 34879 6500 34935 6502
rect 34959 6500 35015 6502
rect 34719 5466 34775 5468
rect 34799 5466 34855 5468
rect 34879 5466 34935 5468
rect 34959 5466 35015 5468
rect 34719 5414 34765 5466
rect 34765 5414 34775 5466
rect 34799 5414 34829 5466
rect 34829 5414 34841 5466
rect 34841 5414 34855 5466
rect 34879 5414 34893 5466
rect 34893 5414 34905 5466
rect 34905 5414 34935 5466
rect 34959 5414 34969 5466
rect 34969 5414 35015 5466
rect 34719 5412 34775 5414
rect 34799 5412 34855 5414
rect 34879 5412 34935 5414
rect 34959 5412 35015 5414
rect 34719 4378 34775 4380
rect 34799 4378 34855 4380
rect 34879 4378 34935 4380
rect 34959 4378 35015 4380
rect 34719 4326 34765 4378
rect 34765 4326 34775 4378
rect 34799 4326 34829 4378
rect 34829 4326 34841 4378
rect 34841 4326 34855 4378
rect 34879 4326 34893 4378
rect 34893 4326 34905 4378
rect 34905 4326 34935 4378
rect 34959 4326 34969 4378
rect 34969 4326 35015 4378
rect 34719 4324 34775 4326
rect 34799 4324 34855 4326
rect 34879 4324 34935 4326
rect 34959 4324 35015 4326
rect 34719 3290 34775 3292
rect 34799 3290 34855 3292
rect 34879 3290 34935 3292
rect 34959 3290 35015 3292
rect 34719 3238 34765 3290
rect 34765 3238 34775 3290
rect 34799 3238 34829 3290
rect 34829 3238 34841 3290
rect 34841 3238 34855 3290
rect 34879 3238 34893 3290
rect 34893 3238 34905 3290
rect 34905 3238 34935 3290
rect 34959 3238 34969 3290
rect 34969 3238 35015 3290
rect 34719 3236 34775 3238
rect 34799 3236 34855 3238
rect 34879 3236 34935 3238
rect 34959 3236 35015 3238
rect 9396 2202 9452 2204
rect 9476 2202 9532 2204
rect 9556 2202 9612 2204
rect 9636 2202 9692 2204
rect 9396 2150 9442 2202
rect 9442 2150 9452 2202
rect 9476 2150 9506 2202
rect 9506 2150 9518 2202
rect 9518 2150 9532 2202
rect 9556 2150 9570 2202
rect 9570 2150 9582 2202
rect 9582 2150 9612 2202
rect 9636 2150 9646 2202
rect 9646 2150 9692 2202
rect 9396 2148 9452 2150
rect 9476 2148 9532 2150
rect 9556 2148 9612 2150
rect 9636 2148 9692 2150
rect 17837 2202 17893 2204
rect 17917 2202 17973 2204
rect 17997 2202 18053 2204
rect 18077 2202 18133 2204
rect 17837 2150 17883 2202
rect 17883 2150 17893 2202
rect 17917 2150 17947 2202
rect 17947 2150 17959 2202
rect 17959 2150 17973 2202
rect 17997 2150 18011 2202
rect 18011 2150 18023 2202
rect 18023 2150 18053 2202
rect 18077 2150 18087 2202
rect 18087 2150 18133 2202
rect 17837 2148 17893 2150
rect 17917 2148 17973 2150
rect 17997 2148 18053 2150
rect 18077 2148 18133 2150
rect 26278 2202 26334 2204
rect 26358 2202 26414 2204
rect 26438 2202 26494 2204
rect 26518 2202 26574 2204
rect 26278 2150 26324 2202
rect 26324 2150 26334 2202
rect 26358 2150 26388 2202
rect 26388 2150 26400 2202
rect 26400 2150 26414 2202
rect 26438 2150 26452 2202
rect 26452 2150 26464 2202
rect 26464 2150 26494 2202
rect 26518 2150 26528 2202
rect 26528 2150 26574 2202
rect 26278 2148 26334 2150
rect 26358 2148 26414 2150
rect 26438 2148 26494 2150
rect 26518 2148 26574 2150
rect 34719 2202 34775 2204
rect 34799 2202 34855 2204
rect 34879 2202 34935 2204
rect 34959 2202 35015 2204
rect 34719 2150 34765 2202
rect 34765 2150 34775 2202
rect 34799 2150 34829 2202
rect 34829 2150 34841 2202
rect 34841 2150 34855 2202
rect 34879 2150 34893 2202
rect 34893 2150 34905 2202
rect 34905 2150 34935 2202
rect 34959 2150 34969 2202
rect 34969 2150 35015 2202
rect 34719 2148 34775 2150
rect 34799 2148 34855 2150
rect 34879 2148 34935 2150
rect 34959 2148 35015 2150
rect 35162 2080 35218 2136
<< metal3 >>
rect 5166 39744 5482 39745
rect 5166 39680 5172 39744
rect 5236 39680 5252 39744
rect 5316 39680 5332 39744
rect 5396 39680 5412 39744
rect 5476 39680 5482 39744
rect 5166 39679 5482 39680
rect 13607 39744 13923 39745
rect 13607 39680 13613 39744
rect 13677 39680 13693 39744
rect 13757 39680 13773 39744
rect 13837 39680 13853 39744
rect 13917 39680 13923 39744
rect 13607 39679 13923 39680
rect 22048 39744 22364 39745
rect 22048 39680 22054 39744
rect 22118 39680 22134 39744
rect 22198 39680 22214 39744
rect 22278 39680 22294 39744
rect 22358 39680 22364 39744
rect 22048 39679 22364 39680
rect 30489 39744 30805 39745
rect 30489 39680 30495 39744
rect 30559 39680 30575 39744
rect 30639 39680 30655 39744
rect 30719 39680 30735 39744
rect 30799 39680 30805 39744
rect 30489 39679 30805 39680
rect 0 39538 800 39628
rect 933 39538 999 39541
rect 0 39536 999 39538
rect 0 39480 938 39536
rect 994 39480 999 39536
rect 0 39478 999 39480
rect 0 39388 800 39478
rect 933 39475 999 39478
rect 9386 39200 9702 39201
rect 9386 39136 9392 39200
rect 9456 39136 9472 39200
rect 9536 39136 9552 39200
rect 9616 39136 9632 39200
rect 9696 39136 9702 39200
rect 9386 39135 9702 39136
rect 17827 39200 18143 39201
rect 17827 39136 17833 39200
rect 17897 39136 17913 39200
rect 17977 39136 17993 39200
rect 18057 39136 18073 39200
rect 18137 39136 18143 39200
rect 17827 39135 18143 39136
rect 26268 39200 26584 39201
rect 26268 39136 26274 39200
rect 26338 39136 26354 39200
rect 26418 39136 26434 39200
rect 26498 39136 26514 39200
rect 26578 39136 26584 39200
rect 26268 39135 26584 39136
rect 34709 39200 35025 39201
rect 34709 39136 34715 39200
rect 34779 39136 34795 39200
rect 34859 39136 34875 39200
rect 34939 39136 34955 39200
rect 35019 39136 35025 39200
rect 34709 39135 35025 39136
rect 5166 38656 5482 38657
rect 5166 38592 5172 38656
rect 5236 38592 5252 38656
rect 5316 38592 5332 38656
rect 5396 38592 5412 38656
rect 5476 38592 5482 38656
rect 5166 38591 5482 38592
rect 13607 38656 13923 38657
rect 13607 38592 13613 38656
rect 13677 38592 13693 38656
rect 13757 38592 13773 38656
rect 13837 38592 13853 38656
rect 13917 38592 13923 38656
rect 13607 38591 13923 38592
rect 22048 38656 22364 38657
rect 22048 38592 22054 38656
rect 22118 38592 22134 38656
rect 22198 38592 22214 38656
rect 22278 38592 22294 38656
rect 22358 38592 22364 38656
rect 22048 38591 22364 38592
rect 30489 38656 30805 38657
rect 30489 38592 30495 38656
rect 30559 38592 30575 38656
rect 30639 38592 30655 38656
rect 30719 38592 30735 38656
rect 30799 38592 30805 38656
rect 30489 38591 30805 38592
rect 9386 38112 9702 38113
rect 9386 38048 9392 38112
rect 9456 38048 9472 38112
rect 9536 38048 9552 38112
rect 9616 38048 9632 38112
rect 9696 38048 9702 38112
rect 9386 38047 9702 38048
rect 17827 38112 18143 38113
rect 17827 38048 17833 38112
rect 17897 38048 17913 38112
rect 17977 38048 17993 38112
rect 18057 38048 18073 38112
rect 18137 38048 18143 38112
rect 17827 38047 18143 38048
rect 26268 38112 26584 38113
rect 26268 38048 26274 38112
rect 26338 38048 26354 38112
rect 26418 38048 26434 38112
rect 26498 38048 26514 38112
rect 26578 38048 26584 38112
rect 26268 38047 26584 38048
rect 34709 38112 35025 38113
rect 34709 38048 34715 38112
rect 34779 38048 34795 38112
rect 34859 38048 34875 38112
rect 34939 38048 34955 38112
rect 35019 38048 35025 38112
rect 34709 38047 35025 38048
rect 5166 37568 5482 37569
rect 5166 37504 5172 37568
rect 5236 37504 5252 37568
rect 5316 37504 5332 37568
rect 5396 37504 5412 37568
rect 5476 37504 5482 37568
rect 5166 37503 5482 37504
rect 13607 37568 13923 37569
rect 13607 37504 13613 37568
rect 13677 37504 13693 37568
rect 13757 37504 13773 37568
rect 13837 37504 13853 37568
rect 13917 37504 13923 37568
rect 13607 37503 13923 37504
rect 22048 37568 22364 37569
rect 22048 37504 22054 37568
rect 22118 37504 22134 37568
rect 22198 37504 22214 37568
rect 22278 37504 22294 37568
rect 22358 37504 22364 37568
rect 22048 37503 22364 37504
rect 30489 37568 30805 37569
rect 30489 37504 30495 37568
rect 30559 37504 30575 37568
rect 30639 37504 30655 37568
rect 30719 37504 30735 37568
rect 30799 37504 30805 37568
rect 30489 37503 30805 37504
rect 9386 37024 9702 37025
rect 9386 36960 9392 37024
rect 9456 36960 9472 37024
rect 9536 36960 9552 37024
rect 9616 36960 9632 37024
rect 9696 36960 9702 37024
rect 9386 36959 9702 36960
rect 17827 37024 18143 37025
rect 17827 36960 17833 37024
rect 17897 36960 17913 37024
rect 17977 36960 17993 37024
rect 18057 36960 18073 37024
rect 18137 36960 18143 37024
rect 17827 36959 18143 36960
rect 26268 37024 26584 37025
rect 26268 36960 26274 37024
rect 26338 36960 26354 37024
rect 26418 36960 26434 37024
rect 26498 36960 26514 37024
rect 26578 36960 26584 37024
rect 26268 36959 26584 36960
rect 34709 37024 35025 37025
rect 34709 36960 34715 37024
rect 34779 36960 34795 37024
rect 34859 36960 34875 37024
rect 34939 36960 34955 37024
rect 35019 36960 35025 37024
rect 34709 36959 35025 36960
rect 5166 36480 5482 36481
rect 5166 36416 5172 36480
rect 5236 36416 5252 36480
rect 5316 36416 5332 36480
rect 5396 36416 5412 36480
rect 5476 36416 5482 36480
rect 5166 36415 5482 36416
rect 13607 36480 13923 36481
rect 13607 36416 13613 36480
rect 13677 36416 13693 36480
rect 13757 36416 13773 36480
rect 13837 36416 13853 36480
rect 13917 36416 13923 36480
rect 13607 36415 13923 36416
rect 22048 36480 22364 36481
rect 22048 36416 22054 36480
rect 22118 36416 22134 36480
rect 22198 36416 22214 36480
rect 22278 36416 22294 36480
rect 22358 36416 22364 36480
rect 22048 36415 22364 36416
rect 30489 36480 30805 36481
rect 30489 36416 30495 36480
rect 30559 36416 30575 36480
rect 30639 36416 30655 36480
rect 30719 36416 30735 36480
rect 30799 36416 30805 36480
rect 30489 36415 30805 36416
rect 9386 35936 9702 35937
rect 9386 35872 9392 35936
rect 9456 35872 9472 35936
rect 9536 35872 9552 35936
rect 9616 35872 9632 35936
rect 9696 35872 9702 35936
rect 9386 35871 9702 35872
rect 17827 35936 18143 35937
rect 17827 35872 17833 35936
rect 17897 35872 17913 35936
rect 17977 35872 17993 35936
rect 18057 35872 18073 35936
rect 18137 35872 18143 35936
rect 17827 35871 18143 35872
rect 26268 35936 26584 35937
rect 26268 35872 26274 35936
rect 26338 35872 26354 35936
rect 26418 35872 26434 35936
rect 26498 35872 26514 35936
rect 26578 35872 26584 35936
rect 26268 35871 26584 35872
rect 34709 35936 35025 35937
rect 34709 35872 34715 35936
rect 34779 35872 34795 35936
rect 34859 35872 34875 35936
rect 34939 35872 34955 35936
rect 35019 35872 35025 35936
rect 34709 35871 35025 35872
rect 5166 35392 5482 35393
rect 5166 35328 5172 35392
rect 5236 35328 5252 35392
rect 5316 35328 5332 35392
rect 5396 35328 5412 35392
rect 5476 35328 5482 35392
rect 5166 35327 5482 35328
rect 13607 35392 13923 35393
rect 13607 35328 13613 35392
rect 13677 35328 13693 35392
rect 13757 35328 13773 35392
rect 13837 35328 13853 35392
rect 13917 35328 13923 35392
rect 13607 35327 13923 35328
rect 22048 35392 22364 35393
rect 22048 35328 22054 35392
rect 22118 35328 22134 35392
rect 22198 35328 22214 35392
rect 22278 35328 22294 35392
rect 22358 35328 22364 35392
rect 22048 35327 22364 35328
rect 30489 35392 30805 35393
rect 30489 35328 30495 35392
rect 30559 35328 30575 35392
rect 30639 35328 30655 35392
rect 30719 35328 30735 35392
rect 30799 35328 30805 35392
rect 30489 35327 30805 35328
rect 9386 34848 9702 34849
rect 9386 34784 9392 34848
rect 9456 34784 9472 34848
rect 9536 34784 9552 34848
rect 9616 34784 9632 34848
rect 9696 34784 9702 34848
rect 9386 34783 9702 34784
rect 17827 34848 18143 34849
rect 17827 34784 17833 34848
rect 17897 34784 17913 34848
rect 17977 34784 17993 34848
rect 18057 34784 18073 34848
rect 18137 34784 18143 34848
rect 17827 34783 18143 34784
rect 26268 34848 26584 34849
rect 26268 34784 26274 34848
rect 26338 34784 26354 34848
rect 26418 34784 26434 34848
rect 26498 34784 26514 34848
rect 26578 34784 26584 34848
rect 26268 34783 26584 34784
rect 34709 34848 35025 34849
rect 34709 34784 34715 34848
rect 34779 34784 34795 34848
rect 34859 34784 34875 34848
rect 34939 34784 34955 34848
rect 35019 34784 35025 34848
rect 34709 34783 35025 34784
rect 5166 34304 5482 34305
rect 5166 34240 5172 34304
rect 5236 34240 5252 34304
rect 5316 34240 5332 34304
rect 5396 34240 5412 34304
rect 5476 34240 5482 34304
rect 5166 34239 5482 34240
rect 13607 34304 13923 34305
rect 13607 34240 13613 34304
rect 13677 34240 13693 34304
rect 13757 34240 13773 34304
rect 13837 34240 13853 34304
rect 13917 34240 13923 34304
rect 13607 34239 13923 34240
rect 22048 34304 22364 34305
rect 22048 34240 22054 34304
rect 22118 34240 22134 34304
rect 22198 34240 22214 34304
rect 22278 34240 22294 34304
rect 22358 34240 22364 34304
rect 22048 34239 22364 34240
rect 30489 34304 30805 34305
rect 30489 34240 30495 34304
rect 30559 34240 30575 34304
rect 30639 34240 30655 34304
rect 30719 34240 30735 34304
rect 30799 34240 30805 34304
rect 30489 34239 30805 34240
rect 9386 33760 9702 33761
rect 9386 33696 9392 33760
rect 9456 33696 9472 33760
rect 9536 33696 9552 33760
rect 9616 33696 9632 33760
rect 9696 33696 9702 33760
rect 9386 33695 9702 33696
rect 17827 33760 18143 33761
rect 17827 33696 17833 33760
rect 17897 33696 17913 33760
rect 17977 33696 17993 33760
rect 18057 33696 18073 33760
rect 18137 33696 18143 33760
rect 17827 33695 18143 33696
rect 26268 33760 26584 33761
rect 26268 33696 26274 33760
rect 26338 33696 26354 33760
rect 26418 33696 26434 33760
rect 26498 33696 26514 33760
rect 26578 33696 26584 33760
rect 26268 33695 26584 33696
rect 34709 33760 35025 33761
rect 34709 33696 34715 33760
rect 34779 33696 34795 33760
rect 34859 33696 34875 33760
rect 34939 33696 34955 33760
rect 35019 33696 35025 33760
rect 34709 33695 35025 33696
rect 5166 33216 5482 33217
rect 5166 33152 5172 33216
rect 5236 33152 5252 33216
rect 5316 33152 5332 33216
rect 5396 33152 5412 33216
rect 5476 33152 5482 33216
rect 5166 33151 5482 33152
rect 13607 33216 13923 33217
rect 13607 33152 13613 33216
rect 13677 33152 13693 33216
rect 13757 33152 13773 33216
rect 13837 33152 13853 33216
rect 13917 33152 13923 33216
rect 13607 33151 13923 33152
rect 22048 33216 22364 33217
rect 22048 33152 22054 33216
rect 22118 33152 22134 33216
rect 22198 33152 22214 33216
rect 22278 33152 22294 33216
rect 22358 33152 22364 33216
rect 22048 33151 22364 33152
rect 30489 33216 30805 33217
rect 30489 33152 30495 33216
rect 30559 33152 30575 33216
rect 30639 33152 30655 33216
rect 30719 33152 30735 33216
rect 30799 33152 30805 33216
rect 30489 33151 30805 33152
rect 9386 32672 9702 32673
rect 9386 32608 9392 32672
rect 9456 32608 9472 32672
rect 9536 32608 9552 32672
rect 9616 32608 9632 32672
rect 9696 32608 9702 32672
rect 9386 32607 9702 32608
rect 17827 32672 18143 32673
rect 17827 32608 17833 32672
rect 17897 32608 17913 32672
rect 17977 32608 17993 32672
rect 18057 32608 18073 32672
rect 18137 32608 18143 32672
rect 17827 32607 18143 32608
rect 26268 32672 26584 32673
rect 26268 32608 26274 32672
rect 26338 32608 26354 32672
rect 26418 32608 26434 32672
rect 26498 32608 26514 32672
rect 26578 32608 26584 32672
rect 26268 32607 26584 32608
rect 34709 32672 35025 32673
rect 34709 32608 34715 32672
rect 34779 32608 34795 32672
rect 34859 32608 34875 32672
rect 34939 32608 34955 32672
rect 35019 32608 35025 32672
rect 34709 32607 35025 32608
rect 5166 32128 5482 32129
rect 5166 32064 5172 32128
rect 5236 32064 5252 32128
rect 5316 32064 5332 32128
rect 5396 32064 5412 32128
rect 5476 32064 5482 32128
rect 5166 32063 5482 32064
rect 13607 32128 13923 32129
rect 13607 32064 13613 32128
rect 13677 32064 13693 32128
rect 13757 32064 13773 32128
rect 13837 32064 13853 32128
rect 13917 32064 13923 32128
rect 13607 32063 13923 32064
rect 22048 32128 22364 32129
rect 22048 32064 22054 32128
rect 22118 32064 22134 32128
rect 22198 32064 22214 32128
rect 22278 32064 22294 32128
rect 22358 32064 22364 32128
rect 22048 32063 22364 32064
rect 30489 32128 30805 32129
rect 30489 32064 30495 32128
rect 30559 32064 30575 32128
rect 30639 32064 30655 32128
rect 30719 32064 30735 32128
rect 30799 32064 30805 32128
rect 30489 32063 30805 32064
rect 34881 32058 34947 32061
rect 35200 32058 36000 32148
rect 34881 32056 36000 32058
rect 34881 32000 34886 32056
rect 34942 32000 36000 32056
rect 34881 31998 36000 32000
rect 34881 31995 34947 31998
rect 35200 31908 36000 31998
rect 9386 31584 9702 31585
rect 9386 31520 9392 31584
rect 9456 31520 9472 31584
rect 9536 31520 9552 31584
rect 9616 31520 9632 31584
rect 9696 31520 9702 31584
rect 9386 31519 9702 31520
rect 17827 31584 18143 31585
rect 17827 31520 17833 31584
rect 17897 31520 17913 31584
rect 17977 31520 17993 31584
rect 18057 31520 18073 31584
rect 18137 31520 18143 31584
rect 17827 31519 18143 31520
rect 26268 31584 26584 31585
rect 26268 31520 26274 31584
rect 26338 31520 26354 31584
rect 26418 31520 26434 31584
rect 26498 31520 26514 31584
rect 26578 31520 26584 31584
rect 26268 31519 26584 31520
rect 34709 31584 35025 31585
rect 34709 31520 34715 31584
rect 34779 31520 34795 31584
rect 34859 31520 34875 31584
rect 34939 31520 34955 31584
rect 35019 31520 35025 31584
rect 34709 31519 35025 31520
rect 5166 31040 5482 31041
rect 5166 30976 5172 31040
rect 5236 30976 5252 31040
rect 5316 30976 5332 31040
rect 5396 30976 5412 31040
rect 5476 30976 5482 31040
rect 5166 30975 5482 30976
rect 13607 31040 13923 31041
rect 13607 30976 13613 31040
rect 13677 30976 13693 31040
rect 13757 30976 13773 31040
rect 13837 30976 13853 31040
rect 13917 30976 13923 31040
rect 13607 30975 13923 30976
rect 22048 31040 22364 31041
rect 22048 30976 22054 31040
rect 22118 30976 22134 31040
rect 22198 30976 22214 31040
rect 22278 30976 22294 31040
rect 22358 30976 22364 31040
rect 22048 30975 22364 30976
rect 30489 31040 30805 31041
rect 30489 30976 30495 31040
rect 30559 30976 30575 31040
rect 30639 30976 30655 31040
rect 30719 30976 30735 31040
rect 30799 30976 30805 31040
rect 30489 30975 30805 30976
rect 18689 30698 18755 30701
rect 19241 30698 19307 30701
rect 18689 30696 19307 30698
rect 18689 30640 18694 30696
rect 18750 30640 19246 30696
rect 19302 30640 19307 30696
rect 18689 30638 19307 30640
rect 18689 30635 18755 30638
rect 19241 30635 19307 30638
rect 9386 30496 9702 30497
rect 9386 30432 9392 30496
rect 9456 30432 9472 30496
rect 9536 30432 9552 30496
rect 9616 30432 9632 30496
rect 9696 30432 9702 30496
rect 9386 30431 9702 30432
rect 17827 30496 18143 30497
rect 17827 30432 17833 30496
rect 17897 30432 17913 30496
rect 17977 30432 17993 30496
rect 18057 30432 18073 30496
rect 18137 30432 18143 30496
rect 17827 30431 18143 30432
rect 26268 30496 26584 30497
rect 26268 30432 26274 30496
rect 26338 30432 26354 30496
rect 26418 30432 26434 30496
rect 26498 30432 26514 30496
rect 26578 30432 26584 30496
rect 26268 30431 26584 30432
rect 34709 30496 35025 30497
rect 34709 30432 34715 30496
rect 34779 30432 34795 30496
rect 34859 30432 34875 30496
rect 34939 30432 34955 30496
rect 35019 30432 35025 30496
rect 34709 30431 35025 30432
rect 0 30018 800 30108
rect 933 30018 999 30021
rect 0 30016 999 30018
rect 0 29960 938 30016
rect 994 29960 999 30016
rect 0 29958 999 29960
rect 0 29868 800 29958
rect 933 29955 999 29958
rect 5166 29952 5482 29953
rect 5166 29888 5172 29952
rect 5236 29888 5252 29952
rect 5316 29888 5332 29952
rect 5396 29888 5412 29952
rect 5476 29888 5482 29952
rect 5166 29887 5482 29888
rect 13607 29952 13923 29953
rect 13607 29888 13613 29952
rect 13677 29888 13693 29952
rect 13757 29888 13773 29952
rect 13837 29888 13853 29952
rect 13917 29888 13923 29952
rect 13607 29887 13923 29888
rect 22048 29952 22364 29953
rect 22048 29888 22054 29952
rect 22118 29888 22134 29952
rect 22198 29888 22214 29952
rect 22278 29888 22294 29952
rect 22358 29888 22364 29952
rect 22048 29887 22364 29888
rect 30489 29952 30805 29953
rect 30489 29888 30495 29952
rect 30559 29888 30575 29952
rect 30639 29888 30655 29952
rect 30719 29888 30735 29952
rect 30799 29888 30805 29952
rect 30489 29887 30805 29888
rect 9386 29408 9702 29409
rect 9386 29344 9392 29408
rect 9456 29344 9472 29408
rect 9536 29344 9552 29408
rect 9616 29344 9632 29408
rect 9696 29344 9702 29408
rect 9386 29343 9702 29344
rect 17827 29408 18143 29409
rect 17827 29344 17833 29408
rect 17897 29344 17913 29408
rect 17977 29344 17993 29408
rect 18057 29344 18073 29408
rect 18137 29344 18143 29408
rect 17827 29343 18143 29344
rect 26268 29408 26584 29409
rect 26268 29344 26274 29408
rect 26338 29344 26354 29408
rect 26418 29344 26434 29408
rect 26498 29344 26514 29408
rect 26578 29344 26584 29408
rect 26268 29343 26584 29344
rect 34709 29408 35025 29409
rect 34709 29344 34715 29408
rect 34779 29344 34795 29408
rect 34859 29344 34875 29408
rect 34939 29344 34955 29408
rect 35019 29344 35025 29408
rect 34709 29343 35025 29344
rect 20345 29202 20411 29205
rect 20897 29202 20963 29205
rect 20345 29200 20963 29202
rect 20345 29144 20350 29200
rect 20406 29144 20902 29200
rect 20958 29144 20963 29200
rect 20345 29142 20963 29144
rect 20345 29139 20411 29142
rect 20897 29139 20963 29142
rect 5166 28864 5482 28865
rect 5166 28800 5172 28864
rect 5236 28800 5252 28864
rect 5316 28800 5332 28864
rect 5396 28800 5412 28864
rect 5476 28800 5482 28864
rect 5166 28799 5482 28800
rect 13607 28864 13923 28865
rect 13607 28800 13613 28864
rect 13677 28800 13693 28864
rect 13757 28800 13773 28864
rect 13837 28800 13853 28864
rect 13917 28800 13923 28864
rect 13607 28799 13923 28800
rect 22048 28864 22364 28865
rect 22048 28800 22054 28864
rect 22118 28800 22134 28864
rect 22198 28800 22214 28864
rect 22278 28800 22294 28864
rect 22358 28800 22364 28864
rect 22048 28799 22364 28800
rect 30489 28864 30805 28865
rect 30489 28800 30495 28864
rect 30559 28800 30575 28864
rect 30639 28800 30655 28864
rect 30719 28800 30735 28864
rect 30799 28800 30805 28864
rect 30489 28799 30805 28800
rect 9386 28320 9702 28321
rect 9386 28256 9392 28320
rect 9456 28256 9472 28320
rect 9536 28256 9552 28320
rect 9616 28256 9632 28320
rect 9696 28256 9702 28320
rect 9386 28255 9702 28256
rect 17827 28320 18143 28321
rect 17827 28256 17833 28320
rect 17897 28256 17913 28320
rect 17977 28256 17993 28320
rect 18057 28256 18073 28320
rect 18137 28256 18143 28320
rect 17827 28255 18143 28256
rect 26268 28320 26584 28321
rect 26268 28256 26274 28320
rect 26338 28256 26354 28320
rect 26418 28256 26434 28320
rect 26498 28256 26514 28320
rect 26578 28256 26584 28320
rect 26268 28255 26584 28256
rect 34709 28320 35025 28321
rect 34709 28256 34715 28320
rect 34779 28256 34795 28320
rect 34859 28256 34875 28320
rect 34939 28256 34955 28320
rect 35019 28256 35025 28320
rect 34709 28255 35025 28256
rect 5166 27776 5482 27777
rect 5166 27712 5172 27776
rect 5236 27712 5252 27776
rect 5316 27712 5332 27776
rect 5396 27712 5412 27776
rect 5476 27712 5482 27776
rect 5166 27711 5482 27712
rect 13607 27776 13923 27777
rect 13607 27712 13613 27776
rect 13677 27712 13693 27776
rect 13757 27712 13773 27776
rect 13837 27712 13853 27776
rect 13917 27712 13923 27776
rect 13607 27711 13923 27712
rect 22048 27776 22364 27777
rect 22048 27712 22054 27776
rect 22118 27712 22134 27776
rect 22198 27712 22214 27776
rect 22278 27712 22294 27776
rect 22358 27712 22364 27776
rect 22048 27711 22364 27712
rect 30489 27776 30805 27777
rect 30489 27712 30495 27776
rect 30559 27712 30575 27776
rect 30639 27712 30655 27776
rect 30719 27712 30735 27776
rect 30799 27712 30805 27776
rect 30489 27711 30805 27712
rect 20437 27434 20503 27437
rect 20805 27434 20871 27437
rect 20437 27432 20871 27434
rect 20437 27376 20442 27432
rect 20498 27376 20810 27432
rect 20866 27376 20871 27432
rect 20437 27374 20871 27376
rect 20437 27371 20503 27374
rect 20805 27371 20871 27374
rect 9386 27232 9702 27233
rect 9386 27168 9392 27232
rect 9456 27168 9472 27232
rect 9536 27168 9552 27232
rect 9616 27168 9632 27232
rect 9696 27168 9702 27232
rect 9386 27167 9702 27168
rect 17827 27232 18143 27233
rect 17827 27168 17833 27232
rect 17897 27168 17913 27232
rect 17977 27168 17993 27232
rect 18057 27168 18073 27232
rect 18137 27168 18143 27232
rect 17827 27167 18143 27168
rect 26268 27232 26584 27233
rect 26268 27168 26274 27232
rect 26338 27168 26354 27232
rect 26418 27168 26434 27232
rect 26498 27168 26514 27232
rect 26578 27168 26584 27232
rect 26268 27167 26584 27168
rect 34709 27232 35025 27233
rect 34709 27168 34715 27232
rect 34779 27168 34795 27232
rect 34859 27168 34875 27232
rect 34939 27168 34955 27232
rect 35019 27168 35025 27232
rect 34709 27167 35025 27168
rect 20805 27026 20871 27029
rect 21265 27026 21331 27029
rect 20805 27024 21331 27026
rect 20805 26968 20810 27024
rect 20866 26968 21270 27024
rect 21326 26968 21331 27024
rect 20805 26966 21331 26968
rect 20805 26963 20871 26966
rect 21265 26963 21331 26966
rect 20069 26890 20135 26893
rect 21357 26890 21423 26893
rect 20069 26888 21423 26890
rect 20069 26832 20074 26888
rect 20130 26832 21362 26888
rect 21418 26832 21423 26888
rect 20069 26830 21423 26832
rect 20069 26827 20135 26830
rect 21357 26827 21423 26830
rect 5166 26688 5482 26689
rect 5166 26624 5172 26688
rect 5236 26624 5252 26688
rect 5316 26624 5332 26688
rect 5396 26624 5412 26688
rect 5476 26624 5482 26688
rect 5166 26623 5482 26624
rect 13607 26688 13923 26689
rect 13607 26624 13613 26688
rect 13677 26624 13693 26688
rect 13757 26624 13773 26688
rect 13837 26624 13853 26688
rect 13917 26624 13923 26688
rect 13607 26623 13923 26624
rect 22048 26688 22364 26689
rect 22048 26624 22054 26688
rect 22118 26624 22134 26688
rect 22198 26624 22214 26688
rect 22278 26624 22294 26688
rect 22358 26624 22364 26688
rect 22048 26623 22364 26624
rect 30489 26688 30805 26689
rect 30489 26624 30495 26688
rect 30559 26624 30575 26688
rect 30639 26624 30655 26688
rect 30719 26624 30735 26688
rect 30799 26624 30805 26688
rect 30489 26623 30805 26624
rect 20897 26482 20963 26485
rect 21909 26482 21975 26485
rect 20897 26480 21975 26482
rect 20897 26424 20902 26480
rect 20958 26424 21914 26480
rect 21970 26424 21975 26480
rect 20897 26422 21975 26424
rect 20897 26419 20963 26422
rect 21909 26419 21975 26422
rect 20621 26346 20687 26349
rect 21357 26346 21423 26349
rect 25589 26346 25655 26349
rect 20621 26344 25655 26346
rect 20621 26288 20626 26344
rect 20682 26288 21362 26344
rect 21418 26288 25594 26344
rect 25650 26288 25655 26344
rect 20621 26286 25655 26288
rect 20621 26283 20687 26286
rect 21357 26283 21423 26286
rect 25589 26283 25655 26286
rect 9386 26144 9702 26145
rect 9386 26080 9392 26144
rect 9456 26080 9472 26144
rect 9536 26080 9552 26144
rect 9616 26080 9632 26144
rect 9696 26080 9702 26144
rect 9386 26079 9702 26080
rect 17827 26144 18143 26145
rect 17827 26080 17833 26144
rect 17897 26080 17913 26144
rect 17977 26080 17993 26144
rect 18057 26080 18073 26144
rect 18137 26080 18143 26144
rect 17827 26079 18143 26080
rect 26268 26144 26584 26145
rect 26268 26080 26274 26144
rect 26338 26080 26354 26144
rect 26418 26080 26434 26144
rect 26498 26080 26514 26144
rect 26578 26080 26584 26144
rect 26268 26079 26584 26080
rect 34709 26144 35025 26145
rect 34709 26080 34715 26144
rect 34779 26080 34795 26144
rect 34859 26080 34875 26144
rect 34939 26080 34955 26144
rect 35019 26080 35025 26144
rect 34709 26079 35025 26080
rect 5166 25600 5482 25601
rect 5166 25536 5172 25600
rect 5236 25536 5252 25600
rect 5316 25536 5332 25600
rect 5396 25536 5412 25600
rect 5476 25536 5482 25600
rect 5166 25535 5482 25536
rect 13607 25600 13923 25601
rect 13607 25536 13613 25600
rect 13677 25536 13693 25600
rect 13757 25536 13773 25600
rect 13837 25536 13853 25600
rect 13917 25536 13923 25600
rect 13607 25535 13923 25536
rect 22048 25600 22364 25601
rect 22048 25536 22054 25600
rect 22118 25536 22134 25600
rect 22198 25536 22214 25600
rect 22278 25536 22294 25600
rect 22358 25536 22364 25600
rect 22048 25535 22364 25536
rect 30489 25600 30805 25601
rect 30489 25536 30495 25600
rect 30559 25536 30575 25600
rect 30639 25536 30655 25600
rect 30719 25536 30735 25600
rect 30799 25536 30805 25600
rect 30489 25535 30805 25536
rect 29085 25258 29151 25261
rect 30097 25258 30163 25261
rect 29085 25256 30163 25258
rect 29085 25200 29090 25256
rect 29146 25200 30102 25256
rect 30158 25200 30163 25256
rect 29085 25198 30163 25200
rect 29085 25195 29151 25198
rect 30097 25195 30163 25198
rect 9386 25056 9702 25057
rect 9386 24992 9392 25056
rect 9456 24992 9472 25056
rect 9536 24992 9552 25056
rect 9616 24992 9632 25056
rect 9696 24992 9702 25056
rect 9386 24991 9702 24992
rect 17827 25056 18143 25057
rect 17827 24992 17833 25056
rect 17897 24992 17913 25056
rect 17977 24992 17993 25056
rect 18057 24992 18073 25056
rect 18137 24992 18143 25056
rect 17827 24991 18143 24992
rect 26268 25056 26584 25057
rect 26268 24992 26274 25056
rect 26338 24992 26354 25056
rect 26418 24992 26434 25056
rect 26498 24992 26514 25056
rect 26578 24992 26584 25056
rect 26268 24991 26584 24992
rect 34709 25056 35025 25057
rect 34709 24992 34715 25056
rect 34779 24992 34795 25056
rect 34859 24992 34875 25056
rect 34939 24992 34955 25056
rect 35019 24992 35025 25056
rect 34709 24991 35025 24992
rect 5166 24512 5482 24513
rect 5166 24448 5172 24512
rect 5236 24448 5252 24512
rect 5316 24448 5332 24512
rect 5396 24448 5412 24512
rect 5476 24448 5482 24512
rect 5166 24447 5482 24448
rect 13607 24512 13923 24513
rect 13607 24448 13613 24512
rect 13677 24448 13693 24512
rect 13757 24448 13773 24512
rect 13837 24448 13853 24512
rect 13917 24448 13923 24512
rect 13607 24447 13923 24448
rect 22048 24512 22364 24513
rect 22048 24448 22054 24512
rect 22118 24448 22134 24512
rect 22198 24448 22214 24512
rect 22278 24448 22294 24512
rect 22358 24448 22364 24512
rect 22048 24447 22364 24448
rect 30489 24512 30805 24513
rect 30489 24448 30495 24512
rect 30559 24448 30575 24512
rect 30639 24448 30655 24512
rect 30719 24448 30735 24512
rect 30799 24448 30805 24512
rect 30489 24447 30805 24448
rect 9386 23968 9702 23969
rect 9386 23904 9392 23968
rect 9456 23904 9472 23968
rect 9536 23904 9552 23968
rect 9616 23904 9632 23968
rect 9696 23904 9702 23968
rect 9386 23903 9702 23904
rect 17827 23968 18143 23969
rect 17827 23904 17833 23968
rect 17897 23904 17913 23968
rect 17977 23904 17993 23968
rect 18057 23904 18073 23968
rect 18137 23904 18143 23968
rect 17827 23903 18143 23904
rect 26268 23968 26584 23969
rect 26268 23904 26274 23968
rect 26338 23904 26354 23968
rect 26418 23904 26434 23968
rect 26498 23904 26514 23968
rect 26578 23904 26584 23968
rect 26268 23903 26584 23904
rect 34709 23968 35025 23969
rect 34709 23904 34715 23968
rect 34779 23904 34795 23968
rect 34859 23904 34875 23968
rect 34939 23904 34955 23968
rect 35019 23904 35025 23968
rect 34709 23903 35025 23904
rect 5166 23424 5482 23425
rect 5166 23360 5172 23424
rect 5236 23360 5252 23424
rect 5316 23360 5332 23424
rect 5396 23360 5412 23424
rect 5476 23360 5482 23424
rect 5166 23359 5482 23360
rect 13607 23424 13923 23425
rect 13607 23360 13613 23424
rect 13677 23360 13693 23424
rect 13757 23360 13773 23424
rect 13837 23360 13853 23424
rect 13917 23360 13923 23424
rect 13607 23359 13923 23360
rect 22048 23424 22364 23425
rect 22048 23360 22054 23424
rect 22118 23360 22134 23424
rect 22198 23360 22214 23424
rect 22278 23360 22294 23424
rect 22358 23360 22364 23424
rect 22048 23359 22364 23360
rect 30489 23424 30805 23425
rect 30489 23360 30495 23424
rect 30559 23360 30575 23424
rect 30639 23360 30655 23424
rect 30719 23360 30735 23424
rect 30799 23360 30805 23424
rect 30489 23359 30805 23360
rect 9386 22880 9702 22881
rect 9386 22816 9392 22880
rect 9456 22816 9472 22880
rect 9536 22816 9552 22880
rect 9616 22816 9632 22880
rect 9696 22816 9702 22880
rect 9386 22815 9702 22816
rect 17827 22880 18143 22881
rect 17827 22816 17833 22880
rect 17897 22816 17913 22880
rect 17977 22816 17993 22880
rect 18057 22816 18073 22880
rect 18137 22816 18143 22880
rect 17827 22815 18143 22816
rect 26268 22880 26584 22881
rect 26268 22816 26274 22880
rect 26338 22816 26354 22880
rect 26418 22816 26434 22880
rect 26498 22816 26514 22880
rect 26578 22816 26584 22880
rect 26268 22815 26584 22816
rect 34709 22880 35025 22881
rect 34709 22816 34715 22880
rect 34779 22816 34795 22880
rect 34859 22816 34875 22880
rect 34939 22816 34955 22880
rect 35019 22816 35025 22880
rect 34709 22815 35025 22816
rect 5166 22336 5482 22337
rect 5166 22272 5172 22336
rect 5236 22272 5252 22336
rect 5316 22272 5332 22336
rect 5396 22272 5412 22336
rect 5476 22272 5482 22336
rect 5166 22271 5482 22272
rect 13607 22336 13923 22337
rect 13607 22272 13613 22336
rect 13677 22272 13693 22336
rect 13757 22272 13773 22336
rect 13837 22272 13853 22336
rect 13917 22272 13923 22336
rect 13607 22271 13923 22272
rect 22048 22336 22364 22337
rect 22048 22272 22054 22336
rect 22118 22272 22134 22336
rect 22198 22272 22214 22336
rect 22278 22272 22294 22336
rect 22358 22272 22364 22336
rect 22048 22271 22364 22272
rect 30489 22336 30805 22337
rect 30489 22272 30495 22336
rect 30559 22272 30575 22336
rect 30639 22272 30655 22336
rect 30719 22272 30735 22336
rect 30799 22272 30805 22336
rect 30489 22271 30805 22272
rect 34881 21994 34947 21997
rect 34881 21992 35082 21994
rect 34881 21936 34886 21992
rect 34942 21960 35082 21992
rect 34942 21948 35266 21960
rect 34942 21936 36000 21948
rect 34881 21934 36000 21936
rect 34881 21931 34947 21934
rect 35022 21900 36000 21934
rect 9386 21792 9702 21793
rect 9386 21728 9392 21792
rect 9456 21728 9472 21792
rect 9536 21728 9552 21792
rect 9616 21728 9632 21792
rect 9696 21728 9702 21792
rect 9386 21727 9702 21728
rect 17827 21792 18143 21793
rect 17827 21728 17833 21792
rect 17897 21728 17913 21792
rect 17977 21728 17993 21792
rect 18057 21728 18073 21792
rect 18137 21728 18143 21792
rect 17827 21727 18143 21728
rect 26268 21792 26584 21793
rect 26268 21728 26274 21792
rect 26338 21728 26354 21792
rect 26418 21728 26434 21792
rect 26498 21728 26514 21792
rect 26578 21728 26584 21792
rect 26268 21727 26584 21728
rect 34709 21792 35025 21793
rect 34709 21728 34715 21792
rect 34779 21728 34795 21792
rect 34859 21728 34875 21792
rect 34939 21728 34955 21792
rect 35019 21728 35025 21792
rect 34709 21727 35025 21728
rect 35200 21708 36000 21900
rect 5166 21248 5482 21249
rect 5166 21184 5172 21248
rect 5236 21184 5252 21248
rect 5316 21184 5332 21248
rect 5396 21184 5412 21248
rect 5476 21184 5482 21248
rect 5166 21183 5482 21184
rect 13607 21248 13923 21249
rect 13607 21184 13613 21248
rect 13677 21184 13693 21248
rect 13757 21184 13773 21248
rect 13837 21184 13853 21248
rect 13917 21184 13923 21248
rect 13607 21183 13923 21184
rect 22048 21248 22364 21249
rect 22048 21184 22054 21248
rect 22118 21184 22134 21248
rect 22198 21184 22214 21248
rect 22278 21184 22294 21248
rect 22358 21184 22364 21248
rect 22048 21183 22364 21184
rect 30489 21248 30805 21249
rect 30489 21184 30495 21248
rect 30559 21184 30575 21248
rect 30639 21184 30655 21248
rect 30719 21184 30735 21248
rect 30799 21184 30805 21248
rect 30489 21183 30805 21184
rect 9386 20704 9702 20705
rect 9386 20640 9392 20704
rect 9456 20640 9472 20704
rect 9536 20640 9552 20704
rect 9616 20640 9632 20704
rect 9696 20640 9702 20704
rect 9386 20639 9702 20640
rect 17827 20704 18143 20705
rect 17827 20640 17833 20704
rect 17897 20640 17913 20704
rect 17977 20640 17993 20704
rect 18057 20640 18073 20704
rect 18137 20640 18143 20704
rect 17827 20639 18143 20640
rect 26268 20704 26584 20705
rect 26268 20640 26274 20704
rect 26338 20640 26354 20704
rect 26418 20640 26434 20704
rect 26498 20640 26514 20704
rect 26578 20640 26584 20704
rect 26268 20639 26584 20640
rect 34709 20704 35025 20705
rect 34709 20640 34715 20704
rect 34779 20640 34795 20704
rect 34859 20640 34875 20704
rect 34939 20640 34955 20704
rect 35019 20640 35025 20704
rect 34709 20639 35025 20640
rect 5166 20160 5482 20161
rect 5166 20096 5172 20160
rect 5236 20096 5252 20160
rect 5316 20096 5332 20160
rect 5396 20096 5412 20160
rect 5476 20096 5482 20160
rect 5166 20095 5482 20096
rect 13607 20160 13923 20161
rect 13607 20096 13613 20160
rect 13677 20096 13693 20160
rect 13757 20096 13773 20160
rect 13837 20096 13853 20160
rect 13917 20096 13923 20160
rect 13607 20095 13923 20096
rect 22048 20160 22364 20161
rect 22048 20096 22054 20160
rect 22118 20096 22134 20160
rect 22198 20096 22214 20160
rect 22278 20096 22294 20160
rect 22358 20096 22364 20160
rect 22048 20095 22364 20096
rect 30489 20160 30805 20161
rect 30489 20096 30495 20160
rect 30559 20096 30575 20160
rect 30639 20096 30655 20160
rect 30719 20096 30735 20160
rect 30799 20096 30805 20160
rect 30489 20095 30805 20096
rect 0 19818 800 19908
rect 933 19818 999 19821
rect 0 19816 999 19818
rect 0 19760 938 19816
rect 994 19760 999 19816
rect 0 19758 999 19760
rect 0 19668 800 19758
rect 933 19755 999 19758
rect 9386 19616 9702 19617
rect 9386 19552 9392 19616
rect 9456 19552 9472 19616
rect 9536 19552 9552 19616
rect 9616 19552 9632 19616
rect 9696 19552 9702 19616
rect 9386 19551 9702 19552
rect 17827 19616 18143 19617
rect 17827 19552 17833 19616
rect 17897 19552 17913 19616
rect 17977 19552 17993 19616
rect 18057 19552 18073 19616
rect 18137 19552 18143 19616
rect 17827 19551 18143 19552
rect 26268 19616 26584 19617
rect 26268 19552 26274 19616
rect 26338 19552 26354 19616
rect 26418 19552 26434 19616
rect 26498 19552 26514 19616
rect 26578 19552 26584 19616
rect 26268 19551 26584 19552
rect 34709 19616 35025 19617
rect 34709 19552 34715 19616
rect 34779 19552 34795 19616
rect 34859 19552 34875 19616
rect 34939 19552 34955 19616
rect 35019 19552 35025 19616
rect 34709 19551 35025 19552
rect 5166 19072 5482 19073
rect 5166 19008 5172 19072
rect 5236 19008 5252 19072
rect 5316 19008 5332 19072
rect 5396 19008 5412 19072
rect 5476 19008 5482 19072
rect 5166 19007 5482 19008
rect 13607 19072 13923 19073
rect 13607 19008 13613 19072
rect 13677 19008 13693 19072
rect 13757 19008 13773 19072
rect 13837 19008 13853 19072
rect 13917 19008 13923 19072
rect 13607 19007 13923 19008
rect 22048 19072 22364 19073
rect 22048 19008 22054 19072
rect 22118 19008 22134 19072
rect 22198 19008 22214 19072
rect 22278 19008 22294 19072
rect 22358 19008 22364 19072
rect 22048 19007 22364 19008
rect 30489 19072 30805 19073
rect 30489 19008 30495 19072
rect 30559 19008 30575 19072
rect 30639 19008 30655 19072
rect 30719 19008 30735 19072
rect 30799 19008 30805 19072
rect 30489 19007 30805 19008
rect 9386 18528 9702 18529
rect 9386 18464 9392 18528
rect 9456 18464 9472 18528
rect 9536 18464 9552 18528
rect 9616 18464 9632 18528
rect 9696 18464 9702 18528
rect 9386 18463 9702 18464
rect 17827 18528 18143 18529
rect 17827 18464 17833 18528
rect 17897 18464 17913 18528
rect 17977 18464 17993 18528
rect 18057 18464 18073 18528
rect 18137 18464 18143 18528
rect 17827 18463 18143 18464
rect 26268 18528 26584 18529
rect 26268 18464 26274 18528
rect 26338 18464 26354 18528
rect 26418 18464 26434 18528
rect 26498 18464 26514 18528
rect 26578 18464 26584 18528
rect 26268 18463 26584 18464
rect 34709 18528 35025 18529
rect 34709 18464 34715 18528
rect 34779 18464 34795 18528
rect 34859 18464 34875 18528
rect 34939 18464 34955 18528
rect 35019 18464 35025 18528
rect 34709 18463 35025 18464
rect 5166 17984 5482 17985
rect 5166 17920 5172 17984
rect 5236 17920 5252 17984
rect 5316 17920 5332 17984
rect 5396 17920 5412 17984
rect 5476 17920 5482 17984
rect 5166 17919 5482 17920
rect 13607 17984 13923 17985
rect 13607 17920 13613 17984
rect 13677 17920 13693 17984
rect 13757 17920 13773 17984
rect 13837 17920 13853 17984
rect 13917 17920 13923 17984
rect 13607 17919 13923 17920
rect 22048 17984 22364 17985
rect 22048 17920 22054 17984
rect 22118 17920 22134 17984
rect 22198 17920 22214 17984
rect 22278 17920 22294 17984
rect 22358 17920 22364 17984
rect 22048 17919 22364 17920
rect 30489 17984 30805 17985
rect 30489 17920 30495 17984
rect 30559 17920 30575 17984
rect 30639 17920 30655 17984
rect 30719 17920 30735 17984
rect 30799 17920 30805 17984
rect 30489 17919 30805 17920
rect 9386 17440 9702 17441
rect 9386 17376 9392 17440
rect 9456 17376 9472 17440
rect 9536 17376 9552 17440
rect 9616 17376 9632 17440
rect 9696 17376 9702 17440
rect 9386 17375 9702 17376
rect 17827 17440 18143 17441
rect 17827 17376 17833 17440
rect 17897 17376 17913 17440
rect 17977 17376 17993 17440
rect 18057 17376 18073 17440
rect 18137 17376 18143 17440
rect 17827 17375 18143 17376
rect 26268 17440 26584 17441
rect 26268 17376 26274 17440
rect 26338 17376 26354 17440
rect 26418 17376 26434 17440
rect 26498 17376 26514 17440
rect 26578 17376 26584 17440
rect 26268 17375 26584 17376
rect 34709 17440 35025 17441
rect 34709 17376 34715 17440
rect 34779 17376 34795 17440
rect 34859 17376 34875 17440
rect 34939 17376 34955 17440
rect 35019 17376 35025 17440
rect 34709 17375 35025 17376
rect 5166 16896 5482 16897
rect 5166 16832 5172 16896
rect 5236 16832 5252 16896
rect 5316 16832 5332 16896
rect 5396 16832 5412 16896
rect 5476 16832 5482 16896
rect 5166 16831 5482 16832
rect 13607 16896 13923 16897
rect 13607 16832 13613 16896
rect 13677 16832 13693 16896
rect 13757 16832 13773 16896
rect 13837 16832 13853 16896
rect 13917 16832 13923 16896
rect 13607 16831 13923 16832
rect 22048 16896 22364 16897
rect 22048 16832 22054 16896
rect 22118 16832 22134 16896
rect 22198 16832 22214 16896
rect 22278 16832 22294 16896
rect 22358 16832 22364 16896
rect 22048 16831 22364 16832
rect 30489 16896 30805 16897
rect 30489 16832 30495 16896
rect 30559 16832 30575 16896
rect 30639 16832 30655 16896
rect 30719 16832 30735 16896
rect 30799 16832 30805 16896
rect 30489 16831 30805 16832
rect 9386 16352 9702 16353
rect 9386 16288 9392 16352
rect 9456 16288 9472 16352
rect 9536 16288 9552 16352
rect 9616 16288 9632 16352
rect 9696 16288 9702 16352
rect 9386 16287 9702 16288
rect 17827 16352 18143 16353
rect 17827 16288 17833 16352
rect 17897 16288 17913 16352
rect 17977 16288 17993 16352
rect 18057 16288 18073 16352
rect 18137 16288 18143 16352
rect 17827 16287 18143 16288
rect 26268 16352 26584 16353
rect 26268 16288 26274 16352
rect 26338 16288 26354 16352
rect 26418 16288 26434 16352
rect 26498 16288 26514 16352
rect 26578 16288 26584 16352
rect 26268 16287 26584 16288
rect 34709 16352 35025 16353
rect 34709 16288 34715 16352
rect 34779 16288 34795 16352
rect 34859 16288 34875 16352
rect 34939 16288 34955 16352
rect 35019 16288 35025 16352
rect 34709 16287 35025 16288
rect 5166 15808 5482 15809
rect 5166 15744 5172 15808
rect 5236 15744 5252 15808
rect 5316 15744 5332 15808
rect 5396 15744 5412 15808
rect 5476 15744 5482 15808
rect 5166 15743 5482 15744
rect 13607 15808 13923 15809
rect 13607 15744 13613 15808
rect 13677 15744 13693 15808
rect 13757 15744 13773 15808
rect 13837 15744 13853 15808
rect 13917 15744 13923 15808
rect 13607 15743 13923 15744
rect 22048 15808 22364 15809
rect 22048 15744 22054 15808
rect 22118 15744 22134 15808
rect 22198 15744 22214 15808
rect 22278 15744 22294 15808
rect 22358 15744 22364 15808
rect 22048 15743 22364 15744
rect 30489 15808 30805 15809
rect 30489 15744 30495 15808
rect 30559 15744 30575 15808
rect 30639 15744 30655 15808
rect 30719 15744 30735 15808
rect 30799 15744 30805 15808
rect 30489 15743 30805 15744
rect 9386 15264 9702 15265
rect 9386 15200 9392 15264
rect 9456 15200 9472 15264
rect 9536 15200 9552 15264
rect 9616 15200 9632 15264
rect 9696 15200 9702 15264
rect 9386 15199 9702 15200
rect 17827 15264 18143 15265
rect 17827 15200 17833 15264
rect 17897 15200 17913 15264
rect 17977 15200 17993 15264
rect 18057 15200 18073 15264
rect 18137 15200 18143 15264
rect 17827 15199 18143 15200
rect 26268 15264 26584 15265
rect 26268 15200 26274 15264
rect 26338 15200 26354 15264
rect 26418 15200 26434 15264
rect 26498 15200 26514 15264
rect 26578 15200 26584 15264
rect 26268 15199 26584 15200
rect 34709 15264 35025 15265
rect 34709 15200 34715 15264
rect 34779 15200 34795 15264
rect 34859 15200 34875 15264
rect 34939 15200 34955 15264
rect 35019 15200 35025 15264
rect 34709 15199 35025 15200
rect 5166 14720 5482 14721
rect 5166 14656 5172 14720
rect 5236 14656 5252 14720
rect 5316 14656 5332 14720
rect 5396 14656 5412 14720
rect 5476 14656 5482 14720
rect 5166 14655 5482 14656
rect 13607 14720 13923 14721
rect 13607 14656 13613 14720
rect 13677 14656 13693 14720
rect 13757 14656 13773 14720
rect 13837 14656 13853 14720
rect 13917 14656 13923 14720
rect 13607 14655 13923 14656
rect 22048 14720 22364 14721
rect 22048 14656 22054 14720
rect 22118 14656 22134 14720
rect 22198 14656 22214 14720
rect 22278 14656 22294 14720
rect 22358 14656 22364 14720
rect 22048 14655 22364 14656
rect 30489 14720 30805 14721
rect 30489 14656 30495 14720
rect 30559 14656 30575 14720
rect 30639 14656 30655 14720
rect 30719 14656 30735 14720
rect 30799 14656 30805 14720
rect 30489 14655 30805 14656
rect 9386 14176 9702 14177
rect 9386 14112 9392 14176
rect 9456 14112 9472 14176
rect 9536 14112 9552 14176
rect 9616 14112 9632 14176
rect 9696 14112 9702 14176
rect 9386 14111 9702 14112
rect 17827 14176 18143 14177
rect 17827 14112 17833 14176
rect 17897 14112 17913 14176
rect 17977 14112 17993 14176
rect 18057 14112 18073 14176
rect 18137 14112 18143 14176
rect 17827 14111 18143 14112
rect 26268 14176 26584 14177
rect 26268 14112 26274 14176
rect 26338 14112 26354 14176
rect 26418 14112 26434 14176
rect 26498 14112 26514 14176
rect 26578 14112 26584 14176
rect 26268 14111 26584 14112
rect 34709 14176 35025 14177
rect 34709 14112 34715 14176
rect 34779 14112 34795 14176
rect 34859 14112 34875 14176
rect 34939 14112 34955 14176
rect 35019 14112 35025 14176
rect 34709 14111 35025 14112
rect 5166 13632 5482 13633
rect 5166 13568 5172 13632
rect 5236 13568 5252 13632
rect 5316 13568 5332 13632
rect 5396 13568 5412 13632
rect 5476 13568 5482 13632
rect 5166 13567 5482 13568
rect 13607 13632 13923 13633
rect 13607 13568 13613 13632
rect 13677 13568 13693 13632
rect 13757 13568 13773 13632
rect 13837 13568 13853 13632
rect 13917 13568 13923 13632
rect 13607 13567 13923 13568
rect 22048 13632 22364 13633
rect 22048 13568 22054 13632
rect 22118 13568 22134 13632
rect 22198 13568 22214 13632
rect 22278 13568 22294 13632
rect 22358 13568 22364 13632
rect 22048 13567 22364 13568
rect 30489 13632 30805 13633
rect 30489 13568 30495 13632
rect 30559 13568 30575 13632
rect 30639 13568 30655 13632
rect 30719 13568 30735 13632
rect 30799 13568 30805 13632
rect 30489 13567 30805 13568
rect 9386 13088 9702 13089
rect 9386 13024 9392 13088
rect 9456 13024 9472 13088
rect 9536 13024 9552 13088
rect 9616 13024 9632 13088
rect 9696 13024 9702 13088
rect 9386 13023 9702 13024
rect 17827 13088 18143 13089
rect 17827 13024 17833 13088
rect 17897 13024 17913 13088
rect 17977 13024 17993 13088
rect 18057 13024 18073 13088
rect 18137 13024 18143 13088
rect 17827 13023 18143 13024
rect 26268 13088 26584 13089
rect 26268 13024 26274 13088
rect 26338 13024 26354 13088
rect 26418 13024 26434 13088
rect 26498 13024 26514 13088
rect 26578 13024 26584 13088
rect 26268 13023 26584 13024
rect 34709 13088 35025 13089
rect 34709 13024 34715 13088
rect 34779 13024 34795 13088
rect 34859 13024 34875 13088
rect 34939 13024 34955 13088
rect 35019 13024 35025 13088
rect 34709 13023 35025 13024
rect 5166 12544 5482 12545
rect 5166 12480 5172 12544
rect 5236 12480 5252 12544
rect 5316 12480 5332 12544
rect 5396 12480 5412 12544
rect 5476 12480 5482 12544
rect 5166 12479 5482 12480
rect 13607 12544 13923 12545
rect 13607 12480 13613 12544
rect 13677 12480 13693 12544
rect 13757 12480 13773 12544
rect 13837 12480 13853 12544
rect 13917 12480 13923 12544
rect 13607 12479 13923 12480
rect 22048 12544 22364 12545
rect 22048 12480 22054 12544
rect 22118 12480 22134 12544
rect 22198 12480 22214 12544
rect 22278 12480 22294 12544
rect 22358 12480 22364 12544
rect 22048 12479 22364 12480
rect 30489 12544 30805 12545
rect 30489 12480 30495 12544
rect 30559 12480 30575 12544
rect 30639 12480 30655 12544
rect 30719 12480 30735 12544
rect 30799 12480 30805 12544
rect 30489 12479 30805 12480
rect 9386 12000 9702 12001
rect 9386 11936 9392 12000
rect 9456 11936 9472 12000
rect 9536 11936 9552 12000
rect 9616 11936 9632 12000
rect 9696 11936 9702 12000
rect 9386 11935 9702 11936
rect 17827 12000 18143 12001
rect 17827 11936 17833 12000
rect 17897 11936 17913 12000
rect 17977 11936 17993 12000
rect 18057 11936 18073 12000
rect 18137 11936 18143 12000
rect 17827 11935 18143 11936
rect 26268 12000 26584 12001
rect 26268 11936 26274 12000
rect 26338 11936 26354 12000
rect 26418 11936 26434 12000
rect 26498 11936 26514 12000
rect 26578 11936 26584 12000
rect 26268 11935 26584 11936
rect 34709 12000 35025 12001
rect 34709 11936 34715 12000
rect 34779 11936 34795 12000
rect 34859 11936 34875 12000
rect 34939 11936 34955 12000
rect 35019 11936 35025 12000
rect 34709 11935 35025 11936
rect 34513 11658 34579 11661
rect 35200 11658 36000 11748
rect 34513 11656 36000 11658
rect 34513 11600 34518 11656
rect 34574 11600 36000 11656
rect 34513 11598 36000 11600
rect 34513 11595 34579 11598
rect 35200 11508 36000 11598
rect 5166 11456 5482 11457
rect 5166 11392 5172 11456
rect 5236 11392 5252 11456
rect 5316 11392 5332 11456
rect 5396 11392 5412 11456
rect 5476 11392 5482 11456
rect 5166 11391 5482 11392
rect 13607 11456 13923 11457
rect 13607 11392 13613 11456
rect 13677 11392 13693 11456
rect 13757 11392 13773 11456
rect 13837 11392 13853 11456
rect 13917 11392 13923 11456
rect 13607 11391 13923 11392
rect 22048 11456 22364 11457
rect 22048 11392 22054 11456
rect 22118 11392 22134 11456
rect 22198 11392 22214 11456
rect 22278 11392 22294 11456
rect 22358 11392 22364 11456
rect 22048 11391 22364 11392
rect 30489 11456 30805 11457
rect 30489 11392 30495 11456
rect 30559 11392 30575 11456
rect 30639 11392 30655 11456
rect 30719 11392 30735 11456
rect 30799 11392 30805 11456
rect 30489 11391 30805 11392
rect 9386 10912 9702 10913
rect 9386 10848 9392 10912
rect 9456 10848 9472 10912
rect 9536 10848 9552 10912
rect 9616 10848 9632 10912
rect 9696 10848 9702 10912
rect 9386 10847 9702 10848
rect 17827 10912 18143 10913
rect 17827 10848 17833 10912
rect 17897 10848 17913 10912
rect 17977 10848 17993 10912
rect 18057 10848 18073 10912
rect 18137 10848 18143 10912
rect 17827 10847 18143 10848
rect 26268 10912 26584 10913
rect 26268 10848 26274 10912
rect 26338 10848 26354 10912
rect 26418 10848 26434 10912
rect 26498 10848 26514 10912
rect 26578 10848 26584 10912
rect 26268 10847 26584 10848
rect 34709 10912 35025 10913
rect 34709 10848 34715 10912
rect 34779 10848 34795 10912
rect 34859 10848 34875 10912
rect 34939 10848 34955 10912
rect 35019 10848 35025 10912
rect 34709 10847 35025 10848
rect 5166 10368 5482 10369
rect 5166 10304 5172 10368
rect 5236 10304 5252 10368
rect 5316 10304 5332 10368
rect 5396 10304 5412 10368
rect 5476 10304 5482 10368
rect 5166 10303 5482 10304
rect 13607 10368 13923 10369
rect 13607 10304 13613 10368
rect 13677 10304 13693 10368
rect 13757 10304 13773 10368
rect 13837 10304 13853 10368
rect 13917 10304 13923 10368
rect 13607 10303 13923 10304
rect 22048 10368 22364 10369
rect 22048 10304 22054 10368
rect 22118 10304 22134 10368
rect 22198 10304 22214 10368
rect 22278 10304 22294 10368
rect 22358 10304 22364 10368
rect 22048 10303 22364 10304
rect 30489 10368 30805 10369
rect 30489 10304 30495 10368
rect 30559 10304 30575 10368
rect 30639 10304 30655 10368
rect 30719 10304 30735 10368
rect 30799 10304 30805 10368
rect 30489 10303 30805 10304
rect 9386 9824 9702 9825
rect 9386 9760 9392 9824
rect 9456 9760 9472 9824
rect 9536 9760 9552 9824
rect 9616 9760 9632 9824
rect 9696 9760 9702 9824
rect 9386 9759 9702 9760
rect 17827 9824 18143 9825
rect 17827 9760 17833 9824
rect 17897 9760 17913 9824
rect 17977 9760 17993 9824
rect 18057 9760 18073 9824
rect 18137 9760 18143 9824
rect 17827 9759 18143 9760
rect 26268 9824 26584 9825
rect 26268 9760 26274 9824
rect 26338 9760 26354 9824
rect 26418 9760 26434 9824
rect 26498 9760 26514 9824
rect 26578 9760 26584 9824
rect 26268 9759 26584 9760
rect 34709 9824 35025 9825
rect 34709 9760 34715 9824
rect 34779 9760 34795 9824
rect 34859 9760 34875 9824
rect 34939 9760 34955 9824
rect 35019 9760 35025 9824
rect 34709 9759 35025 9760
rect 0 9618 800 9708
rect 1393 9618 1459 9621
rect 0 9616 1459 9618
rect 0 9560 1398 9616
rect 1454 9560 1459 9616
rect 0 9558 1459 9560
rect 0 9468 800 9558
rect 1393 9555 1459 9558
rect 5166 9280 5482 9281
rect 5166 9216 5172 9280
rect 5236 9216 5252 9280
rect 5316 9216 5332 9280
rect 5396 9216 5412 9280
rect 5476 9216 5482 9280
rect 5166 9215 5482 9216
rect 13607 9280 13923 9281
rect 13607 9216 13613 9280
rect 13677 9216 13693 9280
rect 13757 9216 13773 9280
rect 13837 9216 13853 9280
rect 13917 9216 13923 9280
rect 13607 9215 13923 9216
rect 22048 9280 22364 9281
rect 22048 9216 22054 9280
rect 22118 9216 22134 9280
rect 22198 9216 22214 9280
rect 22278 9216 22294 9280
rect 22358 9216 22364 9280
rect 22048 9215 22364 9216
rect 30489 9280 30805 9281
rect 30489 9216 30495 9280
rect 30559 9216 30575 9280
rect 30639 9216 30655 9280
rect 30719 9216 30735 9280
rect 30799 9216 30805 9280
rect 30489 9215 30805 9216
rect 9386 8736 9702 8737
rect 9386 8672 9392 8736
rect 9456 8672 9472 8736
rect 9536 8672 9552 8736
rect 9616 8672 9632 8736
rect 9696 8672 9702 8736
rect 9386 8671 9702 8672
rect 17827 8736 18143 8737
rect 17827 8672 17833 8736
rect 17897 8672 17913 8736
rect 17977 8672 17993 8736
rect 18057 8672 18073 8736
rect 18137 8672 18143 8736
rect 17827 8671 18143 8672
rect 26268 8736 26584 8737
rect 26268 8672 26274 8736
rect 26338 8672 26354 8736
rect 26418 8672 26434 8736
rect 26498 8672 26514 8736
rect 26578 8672 26584 8736
rect 26268 8671 26584 8672
rect 34709 8736 35025 8737
rect 34709 8672 34715 8736
rect 34779 8672 34795 8736
rect 34859 8672 34875 8736
rect 34939 8672 34955 8736
rect 35019 8672 35025 8736
rect 34709 8671 35025 8672
rect 5166 8192 5482 8193
rect 5166 8128 5172 8192
rect 5236 8128 5252 8192
rect 5316 8128 5332 8192
rect 5396 8128 5412 8192
rect 5476 8128 5482 8192
rect 5166 8127 5482 8128
rect 13607 8192 13923 8193
rect 13607 8128 13613 8192
rect 13677 8128 13693 8192
rect 13757 8128 13773 8192
rect 13837 8128 13853 8192
rect 13917 8128 13923 8192
rect 13607 8127 13923 8128
rect 22048 8192 22364 8193
rect 22048 8128 22054 8192
rect 22118 8128 22134 8192
rect 22198 8128 22214 8192
rect 22278 8128 22294 8192
rect 22358 8128 22364 8192
rect 22048 8127 22364 8128
rect 30489 8192 30805 8193
rect 30489 8128 30495 8192
rect 30559 8128 30575 8192
rect 30639 8128 30655 8192
rect 30719 8128 30735 8192
rect 30799 8128 30805 8192
rect 30489 8127 30805 8128
rect 9386 7648 9702 7649
rect 9386 7584 9392 7648
rect 9456 7584 9472 7648
rect 9536 7584 9552 7648
rect 9616 7584 9632 7648
rect 9696 7584 9702 7648
rect 9386 7583 9702 7584
rect 17827 7648 18143 7649
rect 17827 7584 17833 7648
rect 17897 7584 17913 7648
rect 17977 7584 17993 7648
rect 18057 7584 18073 7648
rect 18137 7584 18143 7648
rect 17827 7583 18143 7584
rect 26268 7648 26584 7649
rect 26268 7584 26274 7648
rect 26338 7584 26354 7648
rect 26418 7584 26434 7648
rect 26498 7584 26514 7648
rect 26578 7584 26584 7648
rect 26268 7583 26584 7584
rect 34709 7648 35025 7649
rect 34709 7584 34715 7648
rect 34779 7584 34795 7648
rect 34859 7584 34875 7648
rect 34939 7584 34955 7648
rect 35019 7584 35025 7648
rect 34709 7583 35025 7584
rect 5166 7104 5482 7105
rect 5166 7040 5172 7104
rect 5236 7040 5252 7104
rect 5316 7040 5332 7104
rect 5396 7040 5412 7104
rect 5476 7040 5482 7104
rect 5166 7039 5482 7040
rect 13607 7104 13923 7105
rect 13607 7040 13613 7104
rect 13677 7040 13693 7104
rect 13757 7040 13773 7104
rect 13837 7040 13853 7104
rect 13917 7040 13923 7104
rect 13607 7039 13923 7040
rect 22048 7104 22364 7105
rect 22048 7040 22054 7104
rect 22118 7040 22134 7104
rect 22198 7040 22214 7104
rect 22278 7040 22294 7104
rect 22358 7040 22364 7104
rect 22048 7039 22364 7040
rect 30489 7104 30805 7105
rect 30489 7040 30495 7104
rect 30559 7040 30575 7104
rect 30639 7040 30655 7104
rect 30719 7040 30735 7104
rect 30799 7040 30805 7104
rect 30489 7039 30805 7040
rect 9386 6560 9702 6561
rect 9386 6496 9392 6560
rect 9456 6496 9472 6560
rect 9536 6496 9552 6560
rect 9616 6496 9632 6560
rect 9696 6496 9702 6560
rect 9386 6495 9702 6496
rect 17827 6560 18143 6561
rect 17827 6496 17833 6560
rect 17897 6496 17913 6560
rect 17977 6496 17993 6560
rect 18057 6496 18073 6560
rect 18137 6496 18143 6560
rect 17827 6495 18143 6496
rect 26268 6560 26584 6561
rect 26268 6496 26274 6560
rect 26338 6496 26354 6560
rect 26418 6496 26434 6560
rect 26498 6496 26514 6560
rect 26578 6496 26584 6560
rect 26268 6495 26584 6496
rect 34709 6560 35025 6561
rect 34709 6496 34715 6560
rect 34779 6496 34795 6560
rect 34859 6496 34875 6560
rect 34939 6496 34955 6560
rect 35019 6496 35025 6560
rect 34709 6495 35025 6496
rect 5166 6016 5482 6017
rect 5166 5952 5172 6016
rect 5236 5952 5252 6016
rect 5316 5952 5332 6016
rect 5396 5952 5412 6016
rect 5476 5952 5482 6016
rect 5166 5951 5482 5952
rect 13607 6016 13923 6017
rect 13607 5952 13613 6016
rect 13677 5952 13693 6016
rect 13757 5952 13773 6016
rect 13837 5952 13853 6016
rect 13917 5952 13923 6016
rect 13607 5951 13923 5952
rect 22048 6016 22364 6017
rect 22048 5952 22054 6016
rect 22118 5952 22134 6016
rect 22198 5952 22214 6016
rect 22278 5952 22294 6016
rect 22358 5952 22364 6016
rect 22048 5951 22364 5952
rect 30489 6016 30805 6017
rect 30489 5952 30495 6016
rect 30559 5952 30575 6016
rect 30639 5952 30655 6016
rect 30719 5952 30735 6016
rect 30799 5952 30805 6016
rect 30489 5951 30805 5952
rect 9386 5472 9702 5473
rect 9386 5408 9392 5472
rect 9456 5408 9472 5472
rect 9536 5408 9552 5472
rect 9616 5408 9632 5472
rect 9696 5408 9702 5472
rect 9386 5407 9702 5408
rect 17827 5472 18143 5473
rect 17827 5408 17833 5472
rect 17897 5408 17913 5472
rect 17977 5408 17993 5472
rect 18057 5408 18073 5472
rect 18137 5408 18143 5472
rect 17827 5407 18143 5408
rect 26268 5472 26584 5473
rect 26268 5408 26274 5472
rect 26338 5408 26354 5472
rect 26418 5408 26434 5472
rect 26498 5408 26514 5472
rect 26578 5408 26584 5472
rect 26268 5407 26584 5408
rect 34709 5472 35025 5473
rect 34709 5408 34715 5472
rect 34779 5408 34795 5472
rect 34859 5408 34875 5472
rect 34939 5408 34955 5472
rect 35019 5408 35025 5472
rect 34709 5407 35025 5408
rect 5166 4928 5482 4929
rect 5166 4864 5172 4928
rect 5236 4864 5252 4928
rect 5316 4864 5332 4928
rect 5396 4864 5412 4928
rect 5476 4864 5482 4928
rect 5166 4863 5482 4864
rect 13607 4928 13923 4929
rect 13607 4864 13613 4928
rect 13677 4864 13693 4928
rect 13757 4864 13773 4928
rect 13837 4864 13853 4928
rect 13917 4864 13923 4928
rect 13607 4863 13923 4864
rect 22048 4928 22364 4929
rect 22048 4864 22054 4928
rect 22118 4864 22134 4928
rect 22198 4864 22214 4928
rect 22278 4864 22294 4928
rect 22358 4864 22364 4928
rect 22048 4863 22364 4864
rect 30489 4928 30805 4929
rect 30489 4864 30495 4928
rect 30559 4864 30575 4928
rect 30639 4864 30655 4928
rect 30719 4864 30735 4928
rect 30799 4864 30805 4928
rect 30489 4863 30805 4864
rect 9386 4384 9702 4385
rect 9386 4320 9392 4384
rect 9456 4320 9472 4384
rect 9536 4320 9552 4384
rect 9616 4320 9632 4384
rect 9696 4320 9702 4384
rect 9386 4319 9702 4320
rect 17827 4384 18143 4385
rect 17827 4320 17833 4384
rect 17897 4320 17913 4384
rect 17977 4320 17993 4384
rect 18057 4320 18073 4384
rect 18137 4320 18143 4384
rect 17827 4319 18143 4320
rect 26268 4384 26584 4385
rect 26268 4320 26274 4384
rect 26338 4320 26354 4384
rect 26418 4320 26434 4384
rect 26498 4320 26514 4384
rect 26578 4320 26584 4384
rect 26268 4319 26584 4320
rect 34709 4384 35025 4385
rect 34709 4320 34715 4384
rect 34779 4320 34795 4384
rect 34859 4320 34875 4384
rect 34939 4320 34955 4384
rect 35019 4320 35025 4384
rect 34709 4319 35025 4320
rect 5166 3840 5482 3841
rect 5166 3776 5172 3840
rect 5236 3776 5252 3840
rect 5316 3776 5332 3840
rect 5396 3776 5412 3840
rect 5476 3776 5482 3840
rect 5166 3775 5482 3776
rect 13607 3840 13923 3841
rect 13607 3776 13613 3840
rect 13677 3776 13693 3840
rect 13757 3776 13773 3840
rect 13837 3776 13853 3840
rect 13917 3776 13923 3840
rect 13607 3775 13923 3776
rect 22048 3840 22364 3841
rect 22048 3776 22054 3840
rect 22118 3776 22134 3840
rect 22198 3776 22214 3840
rect 22278 3776 22294 3840
rect 22358 3776 22364 3840
rect 22048 3775 22364 3776
rect 30489 3840 30805 3841
rect 30489 3776 30495 3840
rect 30559 3776 30575 3840
rect 30639 3776 30655 3840
rect 30719 3776 30735 3840
rect 30799 3776 30805 3840
rect 30489 3775 30805 3776
rect 9386 3296 9702 3297
rect 9386 3232 9392 3296
rect 9456 3232 9472 3296
rect 9536 3232 9552 3296
rect 9616 3232 9632 3296
rect 9696 3232 9702 3296
rect 9386 3231 9702 3232
rect 17827 3296 18143 3297
rect 17827 3232 17833 3296
rect 17897 3232 17913 3296
rect 17977 3232 17993 3296
rect 18057 3232 18073 3296
rect 18137 3232 18143 3296
rect 17827 3231 18143 3232
rect 26268 3296 26584 3297
rect 26268 3232 26274 3296
rect 26338 3232 26354 3296
rect 26418 3232 26434 3296
rect 26498 3232 26514 3296
rect 26578 3232 26584 3296
rect 26268 3231 26584 3232
rect 34709 3296 35025 3297
rect 34709 3232 34715 3296
rect 34779 3232 34795 3296
rect 34859 3232 34875 3296
rect 34939 3232 34955 3296
rect 35019 3232 35025 3296
rect 34709 3231 35025 3232
rect 5166 2752 5482 2753
rect 5166 2688 5172 2752
rect 5236 2688 5252 2752
rect 5316 2688 5332 2752
rect 5396 2688 5412 2752
rect 5476 2688 5482 2752
rect 5166 2687 5482 2688
rect 13607 2752 13923 2753
rect 13607 2688 13613 2752
rect 13677 2688 13693 2752
rect 13757 2688 13773 2752
rect 13837 2688 13853 2752
rect 13917 2688 13923 2752
rect 13607 2687 13923 2688
rect 22048 2752 22364 2753
rect 22048 2688 22054 2752
rect 22118 2688 22134 2752
rect 22198 2688 22214 2752
rect 22278 2688 22294 2752
rect 22358 2688 22364 2752
rect 22048 2687 22364 2688
rect 30489 2752 30805 2753
rect 30489 2688 30495 2752
rect 30559 2688 30575 2752
rect 30639 2688 30655 2752
rect 30719 2688 30735 2752
rect 30799 2688 30805 2752
rect 30489 2687 30805 2688
rect 9386 2208 9702 2209
rect 9386 2144 9392 2208
rect 9456 2144 9472 2208
rect 9536 2144 9552 2208
rect 9616 2144 9632 2208
rect 9696 2144 9702 2208
rect 9386 2143 9702 2144
rect 17827 2208 18143 2209
rect 17827 2144 17833 2208
rect 17897 2144 17913 2208
rect 17977 2144 17993 2208
rect 18057 2144 18073 2208
rect 18137 2144 18143 2208
rect 17827 2143 18143 2144
rect 26268 2208 26584 2209
rect 26268 2144 26274 2208
rect 26338 2144 26354 2208
rect 26418 2144 26434 2208
rect 26498 2144 26514 2208
rect 26578 2144 26584 2208
rect 26268 2143 26584 2144
rect 34709 2208 35025 2209
rect 34709 2144 34715 2208
rect 34779 2144 34795 2208
rect 34859 2144 34875 2208
rect 34939 2144 34955 2208
rect 35019 2144 35025 2208
rect 34709 2143 35025 2144
rect 35200 2141 36000 2228
rect 35157 2136 36000 2141
rect 35157 2080 35162 2136
rect 35218 2080 36000 2136
rect 35157 2075 36000 2080
rect 35200 1988 36000 2075
<< via3 >>
rect 5172 39740 5236 39744
rect 5172 39684 5176 39740
rect 5176 39684 5232 39740
rect 5232 39684 5236 39740
rect 5172 39680 5236 39684
rect 5252 39740 5316 39744
rect 5252 39684 5256 39740
rect 5256 39684 5312 39740
rect 5312 39684 5316 39740
rect 5252 39680 5316 39684
rect 5332 39740 5396 39744
rect 5332 39684 5336 39740
rect 5336 39684 5392 39740
rect 5392 39684 5396 39740
rect 5332 39680 5396 39684
rect 5412 39740 5476 39744
rect 5412 39684 5416 39740
rect 5416 39684 5472 39740
rect 5472 39684 5476 39740
rect 5412 39680 5476 39684
rect 13613 39740 13677 39744
rect 13613 39684 13617 39740
rect 13617 39684 13673 39740
rect 13673 39684 13677 39740
rect 13613 39680 13677 39684
rect 13693 39740 13757 39744
rect 13693 39684 13697 39740
rect 13697 39684 13753 39740
rect 13753 39684 13757 39740
rect 13693 39680 13757 39684
rect 13773 39740 13837 39744
rect 13773 39684 13777 39740
rect 13777 39684 13833 39740
rect 13833 39684 13837 39740
rect 13773 39680 13837 39684
rect 13853 39740 13917 39744
rect 13853 39684 13857 39740
rect 13857 39684 13913 39740
rect 13913 39684 13917 39740
rect 13853 39680 13917 39684
rect 22054 39740 22118 39744
rect 22054 39684 22058 39740
rect 22058 39684 22114 39740
rect 22114 39684 22118 39740
rect 22054 39680 22118 39684
rect 22134 39740 22198 39744
rect 22134 39684 22138 39740
rect 22138 39684 22194 39740
rect 22194 39684 22198 39740
rect 22134 39680 22198 39684
rect 22214 39740 22278 39744
rect 22214 39684 22218 39740
rect 22218 39684 22274 39740
rect 22274 39684 22278 39740
rect 22214 39680 22278 39684
rect 22294 39740 22358 39744
rect 22294 39684 22298 39740
rect 22298 39684 22354 39740
rect 22354 39684 22358 39740
rect 22294 39680 22358 39684
rect 30495 39740 30559 39744
rect 30495 39684 30499 39740
rect 30499 39684 30555 39740
rect 30555 39684 30559 39740
rect 30495 39680 30559 39684
rect 30575 39740 30639 39744
rect 30575 39684 30579 39740
rect 30579 39684 30635 39740
rect 30635 39684 30639 39740
rect 30575 39680 30639 39684
rect 30655 39740 30719 39744
rect 30655 39684 30659 39740
rect 30659 39684 30715 39740
rect 30715 39684 30719 39740
rect 30655 39680 30719 39684
rect 30735 39740 30799 39744
rect 30735 39684 30739 39740
rect 30739 39684 30795 39740
rect 30795 39684 30799 39740
rect 30735 39680 30799 39684
rect 9392 39196 9456 39200
rect 9392 39140 9396 39196
rect 9396 39140 9452 39196
rect 9452 39140 9456 39196
rect 9392 39136 9456 39140
rect 9472 39196 9536 39200
rect 9472 39140 9476 39196
rect 9476 39140 9532 39196
rect 9532 39140 9536 39196
rect 9472 39136 9536 39140
rect 9552 39196 9616 39200
rect 9552 39140 9556 39196
rect 9556 39140 9612 39196
rect 9612 39140 9616 39196
rect 9552 39136 9616 39140
rect 9632 39196 9696 39200
rect 9632 39140 9636 39196
rect 9636 39140 9692 39196
rect 9692 39140 9696 39196
rect 9632 39136 9696 39140
rect 17833 39196 17897 39200
rect 17833 39140 17837 39196
rect 17837 39140 17893 39196
rect 17893 39140 17897 39196
rect 17833 39136 17897 39140
rect 17913 39196 17977 39200
rect 17913 39140 17917 39196
rect 17917 39140 17973 39196
rect 17973 39140 17977 39196
rect 17913 39136 17977 39140
rect 17993 39196 18057 39200
rect 17993 39140 17997 39196
rect 17997 39140 18053 39196
rect 18053 39140 18057 39196
rect 17993 39136 18057 39140
rect 18073 39196 18137 39200
rect 18073 39140 18077 39196
rect 18077 39140 18133 39196
rect 18133 39140 18137 39196
rect 18073 39136 18137 39140
rect 26274 39196 26338 39200
rect 26274 39140 26278 39196
rect 26278 39140 26334 39196
rect 26334 39140 26338 39196
rect 26274 39136 26338 39140
rect 26354 39196 26418 39200
rect 26354 39140 26358 39196
rect 26358 39140 26414 39196
rect 26414 39140 26418 39196
rect 26354 39136 26418 39140
rect 26434 39196 26498 39200
rect 26434 39140 26438 39196
rect 26438 39140 26494 39196
rect 26494 39140 26498 39196
rect 26434 39136 26498 39140
rect 26514 39196 26578 39200
rect 26514 39140 26518 39196
rect 26518 39140 26574 39196
rect 26574 39140 26578 39196
rect 26514 39136 26578 39140
rect 34715 39196 34779 39200
rect 34715 39140 34719 39196
rect 34719 39140 34775 39196
rect 34775 39140 34779 39196
rect 34715 39136 34779 39140
rect 34795 39196 34859 39200
rect 34795 39140 34799 39196
rect 34799 39140 34855 39196
rect 34855 39140 34859 39196
rect 34795 39136 34859 39140
rect 34875 39196 34939 39200
rect 34875 39140 34879 39196
rect 34879 39140 34935 39196
rect 34935 39140 34939 39196
rect 34875 39136 34939 39140
rect 34955 39196 35019 39200
rect 34955 39140 34959 39196
rect 34959 39140 35015 39196
rect 35015 39140 35019 39196
rect 34955 39136 35019 39140
rect 5172 38652 5236 38656
rect 5172 38596 5176 38652
rect 5176 38596 5232 38652
rect 5232 38596 5236 38652
rect 5172 38592 5236 38596
rect 5252 38652 5316 38656
rect 5252 38596 5256 38652
rect 5256 38596 5312 38652
rect 5312 38596 5316 38652
rect 5252 38592 5316 38596
rect 5332 38652 5396 38656
rect 5332 38596 5336 38652
rect 5336 38596 5392 38652
rect 5392 38596 5396 38652
rect 5332 38592 5396 38596
rect 5412 38652 5476 38656
rect 5412 38596 5416 38652
rect 5416 38596 5472 38652
rect 5472 38596 5476 38652
rect 5412 38592 5476 38596
rect 13613 38652 13677 38656
rect 13613 38596 13617 38652
rect 13617 38596 13673 38652
rect 13673 38596 13677 38652
rect 13613 38592 13677 38596
rect 13693 38652 13757 38656
rect 13693 38596 13697 38652
rect 13697 38596 13753 38652
rect 13753 38596 13757 38652
rect 13693 38592 13757 38596
rect 13773 38652 13837 38656
rect 13773 38596 13777 38652
rect 13777 38596 13833 38652
rect 13833 38596 13837 38652
rect 13773 38592 13837 38596
rect 13853 38652 13917 38656
rect 13853 38596 13857 38652
rect 13857 38596 13913 38652
rect 13913 38596 13917 38652
rect 13853 38592 13917 38596
rect 22054 38652 22118 38656
rect 22054 38596 22058 38652
rect 22058 38596 22114 38652
rect 22114 38596 22118 38652
rect 22054 38592 22118 38596
rect 22134 38652 22198 38656
rect 22134 38596 22138 38652
rect 22138 38596 22194 38652
rect 22194 38596 22198 38652
rect 22134 38592 22198 38596
rect 22214 38652 22278 38656
rect 22214 38596 22218 38652
rect 22218 38596 22274 38652
rect 22274 38596 22278 38652
rect 22214 38592 22278 38596
rect 22294 38652 22358 38656
rect 22294 38596 22298 38652
rect 22298 38596 22354 38652
rect 22354 38596 22358 38652
rect 22294 38592 22358 38596
rect 30495 38652 30559 38656
rect 30495 38596 30499 38652
rect 30499 38596 30555 38652
rect 30555 38596 30559 38652
rect 30495 38592 30559 38596
rect 30575 38652 30639 38656
rect 30575 38596 30579 38652
rect 30579 38596 30635 38652
rect 30635 38596 30639 38652
rect 30575 38592 30639 38596
rect 30655 38652 30719 38656
rect 30655 38596 30659 38652
rect 30659 38596 30715 38652
rect 30715 38596 30719 38652
rect 30655 38592 30719 38596
rect 30735 38652 30799 38656
rect 30735 38596 30739 38652
rect 30739 38596 30795 38652
rect 30795 38596 30799 38652
rect 30735 38592 30799 38596
rect 9392 38108 9456 38112
rect 9392 38052 9396 38108
rect 9396 38052 9452 38108
rect 9452 38052 9456 38108
rect 9392 38048 9456 38052
rect 9472 38108 9536 38112
rect 9472 38052 9476 38108
rect 9476 38052 9532 38108
rect 9532 38052 9536 38108
rect 9472 38048 9536 38052
rect 9552 38108 9616 38112
rect 9552 38052 9556 38108
rect 9556 38052 9612 38108
rect 9612 38052 9616 38108
rect 9552 38048 9616 38052
rect 9632 38108 9696 38112
rect 9632 38052 9636 38108
rect 9636 38052 9692 38108
rect 9692 38052 9696 38108
rect 9632 38048 9696 38052
rect 17833 38108 17897 38112
rect 17833 38052 17837 38108
rect 17837 38052 17893 38108
rect 17893 38052 17897 38108
rect 17833 38048 17897 38052
rect 17913 38108 17977 38112
rect 17913 38052 17917 38108
rect 17917 38052 17973 38108
rect 17973 38052 17977 38108
rect 17913 38048 17977 38052
rect 17993 38108 18057 38112
rect 17993 38052 17997 38108
rect 17997 38052 18053 38108
rect 18053 38052 18057 38108
rect 17993 38048 18057 38052
rect 18073 38108 18137 38112
rect 18073 38052 18077 38108
rect 18077 38052 18133 38108
rect 18133 38052 18137 38108
rect 18073 38048 18137 38052
rect 26274 38108 26338 38112
rect 26274 38052 26278 38108
rect 26278 38052 26334 38108
rect 26334 38052 26338 38108
rect 26274 38048 26338 38052
rect 26354 38108 26418 38112
rect 26354 38052 26358 38108
rect 26358 38052 26414 38108
rect 26414 38052 26418 38108
rect 26354 38048 26418 38052
rect 26434 38108 26498 38112
rect 26434 38052 26438 38108
rect 26438 38052 26494 38108
rect 26494 38052 26498 38108
rect 26434 38048 26498 38052
rect 26514 38108 26578 38112
rect 26514 38052 26518 38108
rect 26518 38052 26574 38108
rect 26574 38052 26578 38108
rect 26514 38048 26578 38052
rect 34715 38108 34779 38112
rect 34715 38052 34719 38108
rect 34719 38052 34775 38108
rect 34775 38052 34779 38108
rect 34715 38048 34779 38052
rect 34795 38108 34859 38112
rect 34795 38052 34799 38108
rect 34799 38052 34855 38108
rect 34855 38052 34859 38108
rect 34795 38048 34859 38052
rect 34875 38108 34939 38112
rect 34875 38052 34879 38108
rect 34879 38052 34935 38108
rect 34935 38052 34939 38108
rect 34875 38048 34939 38052
rect 34955 38108 35019 38112
rect 34955 38052 34959 38108
rect 34959 38052 35015 38108
rect 35015 38052 35019 38108
rect 34955 38048 35019 38052
rect 5172 37564 5236 37568
rect 5172 37508 5176 37564
rect 5176 37508 5232 37564
rect 5232 37508 5236 37564
rect 5172 37504 5236 37508
rect 5252 37564 5316 37568
rect 5252 37508 5256 37564
rect 5256 37508 5312 37564
rect 5312 37508 5316 37564
rect 5252 37504 5316 37508
rect 5332 37564 5396 37568
rect 5332 37508 5336 37564
rect 5336 37508 5392 37564
rect 5392 37508 5396 37564
rect 5332 37504 5396 37508
rect 5412 37564 5476 37568
rect 5412 37508 5416 37564
rect 5416 37508 5472 37564
rect 5472 37508 5476 37564
rect 5412 37504 5476 37508
rect 13613 37564 13677 37568
rect 13613 37508 13617 37564
rect 13617 37508 13673 37564
rect 13673 37508 13677 37564
rect 13613 37504 13677 37508
rect 13693 37564 13757 37568
rect 13693 37508 13697 37564
rect 13697 37508 13753 37564
rect 13753 37508 13757 37564
rect 13693 37504 13757 37508
rect 13773 37564 13837 37568
rect 13773 37508 13777 37564
rect 13777 37508 13833 37564
rect 13833 37508 13837 37564
rect 13773 37504 13837 37508
rect 13853 37564 13917 37568
rect 13853 37508 13857 37564
rect 13857 37508 13913 37564
rect 13913 37508 13917 37564
rect 13853 37504 13917 37508
rect 22054 37564 22118 37568
rect 22054 37508 22058 37564
rect 22058 37508 22114 37564
rect 22114 37508 22118 37564
rect 22054 37504 22118 37508
rect 22134 37564 22198 37568
rect 22134 37508 22138 37564
rect 22138 37508 22194 37564
rect 22194 37508 22198 37564
rect 22134 37504 22198 37508
rect 22214 37564 22278 37568
rect 22214 37508 22218 37564
rect 22218 37508 22274 37564
rect 22274 37508 22278 37564
rect 22214 37504 22278 37508
rect 22294 37564 22358 37568
rect 22294 37508 22298 37564
rect 22298 37508 22354 37564
rect 22354 37508 22358 37564
rect 22294 37504 22358 37508
rect 30495 37564 30559 37568
rect 30495 37508 30499 37564
rect 30499 37508 30555 37564
rect 30555 37508 30559 37564
rect 30495 37504 30559 37508
rect 30575 37564 30639 37568
rect 30575 37508 30579 37564
rect 30579 37508 30635 37564
rect 30635 37508 30639 37564
rect 30575 37504 30639 37508
rect 30655 37564 30719 37568
rect 30655 37508 30659 37564
rect 30659 37508 30715 37564
rect 30715 37508 30719 37564
rect 30655 37504 30719 37508
rect 30735 37564 30799 37568
rect 30735 37508 30739 37564
rect 30739 37508 30795 37564
rect 30795 37508 30799 37564
rect 30735 37504 30799 37508
rect 9392 37020 9456 37024
rect 9392 36964 9396 37020
rect 9396 36964 9452 37020
rect 9452 36964 9456 37020
rect 9392 36960 9456 36964
rect 9472 37020 9536 37024
rect 9472 36964 9476 37020
rect 9476 36964 9532 37020
rect 9532 36964 9536 37020
rect 9472 36960 9536 36964
rect 9552 37020 9616 37024
rect 9552 36964 9556 37020
rect 9556 36964 9612 37020
rect 9612 36964 9616 37020
rect 9552 36960 9616 36964
rect 9632 37020 9696 37024
rect 9632 36964 9636 37020
rect 9636 36964 9692 37020
rect 9692 36964 9696 37020
rect 9632 36960 9696 36964
rect 17833 37020 17897 37024
rect 17833 36964 17837 37020
rect 17837 36964 17893 37020
rect 17893 36964 17897 37020
rect 17833 36960 17897 36964
rect 17913 37020 17977 37024
rect 17913 36964 17917 37020
rect 17917 36964 17973 37020
rect 17973 36964 17977 37020
rect 17913 36960 17977 36964
rect 17993 37020 18057 37024
rect 17993 36964 17997 37020
rect 17997 36964 18053 37020
rect 18053 36964 18057 37020
rect 17993 36960 18057 36964
rect 18073 37020 18137 37024
rect 18073 36964 18077 37020
rect 18077 36964 18133 37020
rect 18133 36964 18137 37020
rect 18073 36960 18137 36964
rect 26274 37020 26338 37024
rect 26274 36964 26278 37020
rect 26278 36964 26334 37020
rect 26334 36964 26338 37020
rect 26274 36960 26338 36964
rect 26354 37020 26418 37024
rect 26354 36964 26358 37020
rect 26358 36964 26414 37020
rect 26414 36964 26418 37020
rect 26354 36960 26418 36964
rect 26434 37020 26498 37024
rect 26434 36964 26438 37020
rect 26438 36964 26494 37020
rect 26494 36964 26498 37020
rect 26434 36960 26498 36964
rect 26514 37020 26578 37024
rect 26514 36964 26518 37020
rect 26518 36964 26574 37020
rect 26574 36964 26578 37020
rect 26514 36960 26578 36964
rect 34715 37020 34779 37024
rect 34715 36964 34719 37020
rect 34719 36964 34775 37020
rect 34775 36964 34779 37020
rect 34715 36960 34779 36964
rect 34795 37020 34859 37024
rect 34795 36964 34799 37020
rect 34799 36964 34855 37020
rect 34855 36964 34859 37020
rect 34795 36960 34859 36964
rect 34875 37020 34939 37024
rect 34875 36964 34879 37020
rect 34879 36964 34935 37020
rect 34935 36964 34939 37020
rect 34875 36960 34939 36964
rect 34955 37020 35019 37024
rect 34955 36964 34959 37020
rect 34959 36964 35015 37020
rect 35015 36964 35019 37020
rect 34955 36960 35019 36964
rect 5172 36476 5236 36480
rect 5172 36420 5176 36476
rect 5176 36420 5232 36476
rect 5232 36420 5236 36476
rect 5172 36416 5236 36420
rect 5252 36476 5316 36480
rect 5252 36420 5256 36476
rect 5256 36420 5312 36476
rect 5312 36420 5316 36476
rect 5252 36416 5316 36420
rect 5332 36476 5396 36480
rect 5332 36420 5336 36476
rect 5336 36420 5392 36476
rect 5392 36420 5396 36476
rect 5332 36416 5396 36420
rect 5412 36476 5476 36480
rect 5412 36420 5416 36476
rect 5416 36420 5472 36476
rect 5472 36420 5476 36476
rect 5412 36416 5476 36420
rect 13613 36476 13677 36480
rect 13613 36420 13617 36476
rect 13617 36420 13673 36476
rect 13673 36420 13677 36476
rect 13613 36416 13677 36420
rect 13693 36476 13757 36480
rect 13693 36420 13697 36476
rect 13697 36420 13753 36476
rect 13753 36420 13757 36476
rect 13693 36416 13757 36420
rect 13773 36476 13837 36480
rect 13773 36420 13777 36476
rect 13777 36420 13833 36476
rect 13833 36420 13837 36476
rect 13773 36416 13837 36420
rect 13853 36476 13917 36480
rect 13853 36420 13857 36476
rect 13857 36420 13913 36476
rect 13913 36420 13917 36476
rect 13853 36416 13917 36420
rect 22054 36476 22118 36480
rect 22054 36420 22058 36476
rect 22058 36420 22114 36476
rect 22114 36420 22118 36476
rect 22054 36416 22118 36420
rect 22134 36476 22198 36480
rect 22134 36420 22138 36476
rect 22138 36420 22194 36476
rect 22194 36420 22198 36476
rect 22134 36416 22198 36420
rect 22214 36476 22278 36480
rect 22214 36420 22218 36476
rect 22218 36420 22274 36476
rect 22274 36420 22278 36476
rect 22214 36416 22278 36420
rect 22294 36476 22358 36480
rect 22294 36420 22298 36476
rect 22298 36420 22354 36476
rect 22354 36420 22358 36476
rect 22294 36416 22358 36420
rect 30495 36476 30559 36480
rect 30495 36420 30499 36476
rect 30499 36420 30555 36476
rect 30555 36420 30559 36476
rect 30495 36416 30559 36420
rect 30575 36476 30639 36480
rect 30575 36420 30579 36476
rect 30579 36420 30635 36476
rect 30635 36420 30639 36476
rect 30575 36416 30639 36420
rect 30655 36476 30719 36480
rect 30655 36420 30659 36476
rect 30659 36420 30715 36476
rect 30715 36420 30719 36476
rect 30655 36416 30719 36420
rect 30735 36476 30799 36480
rect 30735 36420 30739 36476
rect 30739 36420 30795 36476
rect 30795 36420 30799 36476
rect 30735 36416 30799 36420
rect 9392 35932 9456 35936
rect 9392 35876 9396 35932
rect 9396 35876 9452 35932
rect 9452 35876 9456 35932
rect 9392 35872 9456 35876
rect 9472 35932 9536 35936
rect 9472 35876 9476 35932
rect 9476 35876 9532 35932
rect 9532 35876 9536 35932
rect 9472 35872 9536 35876
rect 9552 35932 9616 35936
rect 9552 35876 9556 35932
rect 9556 35876 9612 35932
rect 9612 35876 9616 35932
rect 9552 35872 9616 35876
rect 9632 35932 9696 35936
rect 9632 35876 9636 35932
rect 9636 35876 9692 35932
rect 9692 35876 9696 35932
rect 9632 35872 9696 35876
rect 17833 35932 17897 35936
rect 17833 35876 17837 35932
rect 17837 35876 17893 35932
rect 17893 35876 17897 35932
rect 17833 35872 17897 35876
rect 17913 35932 17977 35936
rect 17913 35876 17917 35932
rect 17917 35876 17973 35932
rect 17973 35876 17977 35932
rect 17913 35872 17977 35876
rect 17993 35932 18057 35936
rect 17993 35876 17997 35932
rect 17997 35876 18053 35932
rect 18053 35876 18057 35932
rect 17993 35872 18057 35876
rect 18073 35932 18137 35936
rect 18073 35876 18077 35932
rect 18077 35876 18133 35932
rect 18133 35876 18137 35932
rect 18073 35872 18137 35876
rect 26274 35932 26338 35936
rect 26274 35876 26278 35932
rect 26278 35876 26334 35932
rect 26334 35876 26338 35932
rect 26274 35872 26338 35876
rect 26354 35932 26418 35936
rect 26354 35876 26358 35932
rect 26358 35876 26414 35932
rect 26414 35876 26418 35932
rect 26354 35872 26418 35876
rect 26434 35932 26498 35936
rect 26434 35876 26438 35932
rect 26438 35876 26494 35932
rect 26494 35876 26498 35932
rect 26434 35872 26498 35876
rect 26514 35932 26578 35936
rect 26514 35876 26518 35932
rect 26518 35876 26574 35932
rect 26574 35876 26578 35932
rect 26514 35872 26578 35876
rect 34715 35932 34779 35936
rect 34715 35876 34719 35932
rect 34719 35876 34775 35932
rect 34775 35876 34779 35932
rect 34715 35872 34779 35876
rect 34795 35932 34859 35936
rect 34795 35876 34799 35932
rect 34799 35876 34855 35932
rect 34855 35876 34859 35932
rect 34795 35872 34859 35876
rect 34875 35932 34939 35936
rect 34875 35876 34879 35932
rect 34879 35876 34935 35932
rect 34935 35876 34939 35932
rect 34875 35872 34939 35876
rect 34955 35932 35019 35936
rect 34955 35876 34959 35932
rect 34959 35876 35015 35932
rect 35015 35876 35019 35932
rect 34955 35872 35019 35876
rect 5172 35388 5236 35392
rect 5172 35332 5176 35388
rect 5176 35332 5232 35388
rect 5232 35332 5236 35388
rect 5172 35328 5236 35332
rect 5252 35388 5316 35392
rect 5252 35332 5256 35388
rect 5256 35332 5312 35388
rect 5312 35332 5316 35388
rect 5252 35328 5316 35332
rect 5332 35388 5396 35392
rect 5332 35332 5336 35388
rect 5336 35332 5392 35388
rect 5392 35332 5396 35388
rect 5332 35328 5396 35332
rect 5412 35388 5476 35392
rect 5412 35332 5416 35388
rect 5416 35332 5472 35388
rect 5472 35332 5476 35388
rect 5412 35328 5476 35332
rect 13613 35388 13677 35392
rect 13613 35332 13617 35388
rect 13617 35332 13673 35388
rect 13673 35332 13677 35388
rect 13613 35328 13677 35332
rect 13693 35388 13757 35392
rect 13693 35332 13697 35388
rect 13697 35332 13753 35388
rect 13753 35332 13757 35388
rect 13693 35328 13757 35332
rect 13773 35388 13837 35392
rect 13773 35332 13777 35388
rect 13777 35332 13833 35388
rect 13833 35332 13837 35388
rect 13773 35328 13837 35332
rect 13853 35388 13917 35392
rect 13853 35332 13857 35388
rect 13857 35332 13913 35388
rect 13913 35332 13917 35388
rect 13853 35328 13917 35332
rect 22054 35388 22118 35392
rect 22054 35332 22058 35388
rect 22058 35332 22114 35388
rect 22114 35332 22118 35388
rect 22054 35328 22118 35332
rect 22134 35388 22198 35392
rect 22134 35332 22138 35388
rect 22138 35332 22194 35388
rect 22194 35332 22198 35388
rect 22134 35328 22198 35332
rect 22214 35388 22278 35392
rect 22214 35332 22218 35388
rect 22218 35332 22274 35388
rect 22274 35332 22278 35388
rect 22214 35328 22278 35332
rect 22294 35388 22358 35392
rect 22294 35332 22298 35388
rect 22298 35332 22354 35388
rect 22354 35332 22358 35388
rect 22294 35328 22358 35332
rect 30495 35388 30559 35392
rect 30495 35332 30499 35388
rect 30499 35332 30555 35388
rect 30555 35332 30559 35388
rect 30495 35328 30559 35332
rect 30575 35388 30639 35392
rect 30575 35332 30579 35388
rect 30579 35332 30635 35388
rect 30635 35332 30639 35388
rect 30575 35328 30639 35332
rect 30655 35388 30719 35392
rect 30655 35332 30659 35388
rect 30659 35332 30715 35388
rect 30715 35332 30719 35388
rect 30655 35328 30719 35332
rect 30735 35388 30799 35392
rect 30735 35332 30739 35388
rect 30739 35332 30795 35388
rect 30795 35332 30799 35388
rect 30735 35328 30799 35332
rect 9392 34844 9456 34848
rect 9392 34788 9396 34844
rect 9396 34788 9452 34844
rect 9452 34788 9456 34844
rect 9392 34784 9456 34788
rect 9472 34844 9536 34848
rect 9472 34788 9476 34844
rect 9476 34788 9532 34844
rect 9532 34788 9536 34844
rect 9472 34784 9536 34788
rect 9552 34844 9616 34848
rect 9552 34788 9556 34844
rect 9556 34788 9612 34844
rect 9612 34788 9616 34844
rect 9552 34784 9616 34788
rect 9632 34844 9696 34848
rect 9632 34788 9636 34844
rect 9636 34788 9692 34844
rect 9692 34788 9696 34844
rect 9632 34784 9696 34788
rect 17833 34844 17897 34848
rect 17833 34788 17837 34844
rect 17837 34788 17893 34844
rect 17893 34788 17897 34844
rect 17833 34784 17897 34788
rect 17913 34844 17977 34848
rect 17913 34788 17917 34844
rect 17917 34788 17973 34844
rect 17973 34788 17977 34844
rect 17913 34784 17977 34788
rect 17993 34844 18057 34848
rect 17993 34788 17997 34844
rect 17997 34788 18053 34844
rect 18053 34788 18057 34844
rect 17993 34784 18057 34788
rect 18073 34844 18137 34848
rect 18073 34788 18077 34844
rect 18077 34788 18133 34844
rect 18133 34788 18137 34844
rect 18073 34784 18137 34788
rect 26274 34844 26338 34848
rect 26274 34788 26278 34844
rect 26278 34788 26334 34844
rect 26334 34788 26338 34844
rect 26274 34784 26338 34788
rect 26354 34844 26418 34848
rect 26354 34788 26358 34844
rect 26358 34788 26414 34844
rect 26414 34788 26418 34844
rect 26354 34784 26418 34788
rect 26434 34844 26498 34848
rect 26434 34788 26438 34844
rect 26438 34788 26494 34844
rect 26494 34788 26498 34844
rect 26434 34784 26498 34788
rect 26514 34844 26578 34848
rect 26514 34788 26518 34844
rect 26518 34788 26574 34844
rect 26574 34788 26578 34844
rect 26514 34784 26578 34788
rect 34715 34844 34779 34848
rect 34715 34788 34719 34844
rect 34719 34788 34775 34844
rect 34775 34788 34779 34844
rect 34715 34784 34779 34788
rect 34795 34844 34859 34848
rect 34795 34788 34799 34844
rect 34799 34788 34855 34844
rect 34855 34788 34859 34844
rect 34795 34784 34859 34788
rect 34875 34844 34939 34848
rect 34875 34788 34879 34844
rect 34879 34788 34935 34844
rect 34935 34788 34939 34844
rect 34875 34784 34939 34788
rect 34955 34844 35019 34848
rect 34955 34788 34959 34844
rect 34959 34788 35015 34844
rect 35015 34788 35019 34844
rect 34955 34784 35019 34788
rect 5172 34300 5236 34304
rect 5172 34244 5176 34300
rect 5176 34244 5232 34300
rect 5232 34244 5236 34300
rect 5172 34240 5236 34244
rect 5252 34300 5316 34304
rect 5252 34244 5256 34300
rect 5256 34244 5312 34300
rect 5312 34244 5316 34300
rect 5252 34240 5316 34244
rect 5332 34300 5396 34304
rect 5332 34244 5336 34300
rect 5336 34244 5392 34300
rect 5392 34244 5396 34300
rect 5332 34240 5396 34244
rect 5412 34300 5476 34304
rect 5412 34244 5416 34300
rect 5416 34244 5472 34300
rect 5472 34244 5476 34300
rect 5412 34240 5476 34244
rect 13613 34300 13677 34304
rect 13613 34244 13617 34300
rect 13617 34244 13673 34300
rect 13673 34244 13677 34300
rect 13613 34240 13677 34244
rect 13693 34300 13757 34304
rect 13693 34244 13697 34300
rect 13697 34244 13753 34300
rect 13753 34244 13757 34300
rect 13693 34240 13757 34244
rect 13773 34300 13837 34304
rect 13773 34244 13777 34300
rect 13777 34244 13833 34300
rect 13833 34244 13837 34300
rect 13773 34240 13837 34244
rect 13853 34300 13917 34304
rect 13853 34244 13857 34300
rect 13857 34244 13913 34300
rect 13913 34244 13917 34300
rect 13853 34240 13917 34244
rect 22054 34300 22118 34304
rect 22054 34244 22058 34300
rect 22058 34244 22114 34300
rect 22114 34244 22118 34300
rect 22054 34240 22118 34244
rect 22134 34300 22198 34304
rect 22134 34244 22138 34300
rect 22138 34244 22194 34300
rect 22194 34244 22198 34300
rect 22134 34240 22198 34244
rect 22214 34300 22278 34304
rect 22214 34244 22218 34300
rect 22218 34244 22274 34300
rect 22274 34244 22278 34300
rect 22214 34240 22278 34244
rect 22294 34300 22358 34304
rect 22294 34244 22298 34300
rect 22298 34244 22354 34300
rect 22354 34244 22358 34300
rect 22294 34240 22358 34244
rect 30495 34300 30559 34304
rect 30495 34244 30499 34300
rect 30499 34244 30555 34300
rect 30555 34244 30559 34300
rect 30495 34240 30559 34244
rect 30575 34300 30639 34304
rect 30575 34244 30579 34300
rect 30579 34244 30635 34300
rect 30635 34244 30639 34300
rect 30575 34240 30639 34244
rect 30655 34300 30719 34304
rect 30655 34244 30659 34300
rect 30659 34244 30715 34300
rect 30715 34244 30719 34300
rect 30655 34240 30719 34244
rect 30735 34300 30799 34304
rect 30735 34244 30739 34300
rect 30739 34244 30795 34300
rect 30795 34244 30799 34300
rect 30735 34240 30799 34244
rect 9392 33756 9456 33760
rect 9392 33700 9396 33756
rect 9396 33700 9452 33756
rect 9452 33700 9456 33756
rect 9392 33696 9456 33700
rect 9472 33756 9536 33760
rect 9472 33700 9476 33756
rect 9476 33700 9532 33756
rect 9532 33700 9536 33756
rect 9472 33696 9536 33700
rect 9552 33756 9616 33760
rect 9552 33700 9556 33756
rect 9556 33700 9612 33756
rect 9612 33700 9616 33756
rect 9552 33696 9616 33700
rect 9632 33756 9696 33760
rect 9632 33700 9636 33756
rect 9636 33700 9692 33756
rect 9692 33700 9696 33756
rect 9632 33696 9696 33700
rect 17833 33756 17897 33760
rect 17833 33700 17837 33756
rect 17837 33700 17893 33756
rect 17893 33700 17897 33756
rect 17833 33696 17897 33700
rect 17913 33756 17977 33760
rect 17913 33700 17917 33756
rect 17917 33700 17973 33756
rect 17973 33700 17977 33756
rect 17913 33696 17977 33700
rect 17993 33756 18057 33760
rect 17993 33700 17997 33756
rect 17997 33700 18053 33756
rect 18053 33700 18057 33756
rect 17993 33696 18057 33700
rect 18073 33756 18137 33760
rect 18073 33700 18077 33756
rect 18077 33700 18133 33756
rect 18133 33700 18137 33756
rect 18073 33696 18137 33700
rect 26274 33756 26338 33760
rect 26274 33700 26278 33756
rect 26278 33700 26334 33756
rect 26334 33700 26338 33756
rect 26274 33696 26338 33700
rect 26354 33756 26418 33760
rect 26354 33700 26358 33756
rect 26358 33700 26414 33756
rect 26414 33700 26418 33756
rect 26354 33696 26418 33700
rect 26434 33756 26498 33760
rect 26434 33700 26438 33756
rect 26438 33700 26494 33756
rect 26494 33700 26498 33756
rect 26434 33696 26498 33700
rect 26514 33756 26578 33760
rect 26514 33700 26518 33756
rect 26518 33700 26574 33756
rect 26574 33700 26578 33756
rect 26514 33696 26578 33700
rect 34715 33756 34779 33760
rect 34715 33700 34719 33756
rect 34719 33700 34775 33756
rect 34775 33700 34779 33756
rect 34715 33696 34779 33700
rect 34795 33756 34859 33760
rect 34795 33700 34799 33756
rect 34799 33700 34855 33756
rect 34855 33700 34859 33756
rect 34795 33696 34859 33700
rect 34875 33756 34939 33760
rect 34875 33700 34879 33756
rect 34879 33700 34935 33756
rect 34935 33700 34939 33756
rect 34875 33696 34939 33700
rect 34955 33756 35019 33760
rect 34955 33700 34959 33756
rect 34959 33700 35015 33756
rect 35015 33700 35019 33756
rect 34955 33696 35019 33700
rect 5172 33212 5236 33216
rect 5172 33156 5176 33212
rect 5176 33156 5232 33212
rect 5232 33156 5236 33212
rect 5172 33152 5236 33156
rect 5252 33212 5316 33216
rect 5252 33156 5256 33212
rect 5256 33156 5312 33212
rect 5312 33156 5316 33212
rect 5252 33152 5316 33156
rect 5332 33212 5396 33216
rect 5332 33156 5336 33212
rect 5336 33156 5392 33212
rect 5392 33156 5396 33212
rect 5332 33152 5396 33156
rect 5412 33212 5476 33216
rect 5412 33156 5416 33212
rect 5416 33156 5472 33212
rect 5472 33156 5476 33212
rect 5412 33152 5476 33156
rect 13613 33212 13677 33216
rect 13613 33156 13617 33212
rect 13617 33156 13673 33212
rect 13673 33156 13677 33212
rect 13613 33152 13677 33156
rect 13693 33212 13757 33216
rect 13693 33156 13697 33212
rect 13697 33156 13753 33212
rect 13753 33156 13757 33212
rect 13693 33152 13757 33156
rect 13773 33212 13837 33216
rect 13773 33156 13777 33212
rect 13777 33156 13833 33212
rect 13833 33156 13837 33212
rect 13773 33152 13837 33156
rect 13853 33212 13917 33216
rect 13853 33156 13857 33212
rect 13857 33156 13913 33212
rect 13913 33156 13917 33212
rect 13853 33152 13917 33156
rect 22054 33212 22118 33216
rect 22054 33156 22058 33212
rect 22058 33156 22114 33212
rect 22114 33156 22118 33212
rect 22054 33152 22118 33156
rect 22134 33212 22198 33216
rect 22134 33156 22138 33212
rect 22138 33156 22194 33212
rect 22194 33156 22198 33212
rect 22134 33152 22198 33156
rect 22214 33212 22278 33216
rect 22214 33156 22218 33212
rect 22218 33156 22274 33212
rect 22274 33156 22278 33212
rect 22214 33152 22278 33156
rect 22294 33212 22358 33216
rect 22294 33156 22298 33212
rect 22298 33156 22354 33212
rect 22354 33156 22358 33212
rect 22294 33152 22358 33156
rect 30495 33212 30559 33216
rect 30495 33156 30499 33212
rect 30499 33156 30555 33212
rect 30555 33156 30559 33212
rect 30495 33152 30559 33156
rect 30575 33212 30639 33216
rect 30575 33156 30579 33212
rect 30579 33156 30635 33212
rect 30635 33156 30639 33212
rect 30575 33152 30639 33156
rect 30655 33212 30719 33216
rect 30655 33156 30659 33212
rect 30659 33156 30715 33212
rect 30715 33156 30719 33212
rect 30655 33152 30719 33156
rect 30735 33212 30799 33216
rect 30735 33156 30739 33212
rect 30739 33156 30795 33212
rect 30795 33156 30799 33212
rect 30735 33152 30799 33156
rect 9392 32668 9456 32672
rect 9392 32612 9396 32668
rect 9396 32612 9452 32668
rect 9452 32612 9456 32668
rect 9392 32608 9456 32612
rect 9472 32668 9536 32672
rect 9472 32612 9476 32668
rect 9476 32612 9532 32668
rect 9532 32612 9536 32668
rect 9472 32608 9536 32612
rect 9552 32668 9616 32672
rect 9552 32612 9556 32668
rect 9556 32612 9612 32668
rect 9612 32612 9616 32668
rect 9552 32608 9616 32612
rect 9632 32668 9696 32672
rect 9632 32612 9636 32668
rect 9636 32612 9692 32668
rect 9692 32612 9696 32668
rect 9632 32608 9696 32612
rect 17833 32668 17897 32672
rect 17833 32612 17837 32668
rect 17837 32612 17893 32668
rect 17893 32612 17897 32668
rect 17833 32608 17897 32612
rect 17913 32668 17977 32672
rect 17913 32612 17917 32668
rect 17917 32612 17973 32668
rect 17973 32612 17977 32668
rect 17913 32608 17977 32612
rect 17993 32668 18057 32672
rect 17993 32612 17997 32668
rect 17997 32612 18053 32668
rect 18053 32612 18057 32668
rect 17993 32608 18057 32612
rect 18073 32668 18137 32672
rect 18073 32612 18077 32668
rect 18077 32612 18133 32668
rect 18133 32612 18137 32668
rect 18073 32608 18137 32612
rect 26274 32668 26338 32672
rect 26274 32612 26278 32668
rect 26278 32612 26334 32668
rect 26334 32612 26338 32668
rect 26274 32608 26338 32612
rect 26354 32668 26418 32672
rect 26354 32612 26358 32668
rect 26358 32612 26414 32668
rect 26414 32612 26418 32668
rect 26354 32608 26418 32612
rect 26434 32668 26498 32672
rect 26434 32612 26438 32668
rect 26438 32612 26494 32668
rect 26494 32612 26498 32668
rect 26434 32608 26498 32612
rect 26514 32668 26578 32672
rect 26514 32612 26518 32668
rect 26518 32612 26574 32668
rect 26574 32612 26578 32668
rect 26514 32608 26578 32612
rect 34715 32668 34779 32672
rect 34715 32612 34719 32668
rect 34719 32612 34775 32668
rect 34775 32612 34779 32668
rect 34715 32608 34779 32612
rect 34795 32668 34859 32672
rect 34795 32612 34799 32668
rect 34799 32612 34855 32668
rect 34855 32612 34859 32668
rect 34795 32608 34859 32612
rect 34875 32668 34939 32672
rect 34875 32612 34879 32668
rect 34879 32612 34935 32668
rect 34935 32612 34939 32668
rect 34875 32608 34939 32612
rect 34955 32668 35019 32672
rect 34955 32612 34959 32668
rect 34959 32612 35015 32668
rect 35015 32612 35019 32668
rect 34955 32608 35019 32612
rect 5172 32124 5236 32128
rect 5172 32068 5176 32124
rect 5176 32068 5232 32124
rect 5232 32068 5236 32124
rect 5172 32064 5236 32068
rect 5252 32124 5316 32128
rect 5252 32068 5256 32124
rect 5256 32068 5312 32124
rect 5312 32068 5316 32124
rect 5252 32064 5316 32068
rect 5332 32124 5396 32128
rect 5332 32068 5336 32124
rect 5336 32068 5392 32124
rect 5392 32068 5396 32124
rect 5332 32064 5396 32068
rect 5412 32124 5476 32128
rect 5412 32068 5416 32124
rect 5416 32068 5472 32124
rect 5472 32068 5476 32124
rect 5412 32064 5476 32068
rect 13613 32124 13677 32128
rect 13613 32068 13617 32124
rect 13617 32068 13673 32124
rect 13673 32068 13677 32124
rect 13613 32064 13677 32068
rect 13693 32124 13757 32128
rect 13693 32068 13697 32124
rect 13697 32068 13753 32124
rect 13753 32068 13757 32124
rect 13693 32064 13757 32068
rect 13773 32124 13837 32128
rect 13773 32068 13777 32124
rect 13777 32068 13833 32124
rect 13833 32068 13837 32124
rect 13773 32064 13837 32068
rect 13853 32124 13917 32128
rect 13853 32068 13857 32124
rect 13857 32068 13913 32124
rect 13913 32068 13917 32124
rect 13853 32064 13917 32068
rect 22054 32124 22118 32128
rect 22054 32068 22058 32124
rect 22058 32068 22114 32124
rect 22114 32068 22118 32124
rect 22054 32064 22118 32068
rect 22134 32124 22198 32128
rect 22134 32068 22138 32124
rect 22138 32068 22194 32124
rect 22194 32068 22198 32124
rect 22134 32064 22198 32068
rect 22214 32124 22278 32128
rect 22214 32068 22218 32124
rect 22218 32068 22274 32124
rect 22274 32068 22278 32124
rect 22214 32064 22278 32068
rect 22294 32124 22358 32128
rect 22294 32068 22298 32124
rect 22298 32068 22354 32124
rect 22354 32068 22358 32124
rect 22294 32064 22358 32068
rect 30495 32124 30559 32128
rect 30495 32068 30499 32124
rect 30499 32068 30555 32124
rect 30555 32068 30559 32124
rect 30495 32064 30559 32068
rect 30575 32124 30639 32128
rect 30575 32068 30579 32124
rect 30579 32068 30635 32124
rect 30635 32068 30639 32124
rect 30575 32064 30639 32068
rect 30655 32124 30719 32128
rect 30655 32068 30659 32124
rect 30659 32068 30715 32124
rect 30715 32068 30719 32124
rect 30655 32064 30719 32068
rect 30735 32124 30799 32128
rect 30735 32068 30739 32124
rect 30739 32068 30795 32124
rect 30795 32068 30799 32124
rect 30735 32064 30799 32068
rect 9392 31580 9456 31584
rect 9392 31524 9396 31580
rect 9396 31524 9452 31580
rect 9452 31524 9456 31580
rect 9392 31520 9456 31524
rect 9472 31580 9536 31584
rect 9472 31524 9476 31580
rect 9476 31524 9532 31580
rect 9532 31524 9536 31580
rect 9472 31520 9536 31524
rect 9552 31580 9616 31584
rect 9552 31524 9556 31580
rect 9556 31524 9612 31580
rect 9612 31524 9616 31580
rect 9552 31520 9616 31524
rect 9632 31580 9696 31584
rect 9632 31524 9636 31580
rect 9636 31524 9692 31580
rect 9692 31524 9696 31580
rect 9632 31520 9696 31524
rect 17833 31580 17897 31584
rect 17833 31524 17837 31580
rect 17837 31524 17893 31580
rect 17893 31524 17897 31580
rect 17833 31520 17897 31524
rect 17913 31580 17977 31584
rect 17913 31524 17917 31580
rect 17917 31524 17973 31580
rect 17973 31524 17977 31580
rect 17913 31520 17977 31524
rect 17993 31580 18057 31584
rect 17993 31524 17997 31580
rect 17997 31524 18053 31580
rect 18053 31524 18057 31580
rect 17993 31520 18057 31524
rect 18073 31580 18137 31584
rect 18073 31524 18077 31580
rect 18077 31524 18133 31580
rect 18133 31524 18137 31580
rect 18073 31520 18137 31524
rect 26274 31580 26338 31584
rect 26274 31524 26278 31580
rect 26278 31524 26334 31580
rect 26334 31524 26338 31580
rect 26274 31520 26338 31524
rect 26354 31580 26418 31584
rect 26354 31524 26358 31580
rect 26358 31524 26414 31580
rect 26414 31524 26418 31580
rect 26354 31520 26418 31524
rect 26434 31580 26498 31584
rect 26434 31524 26438 31580
rect 26438 31524 26494 31580
rect 26494 31524 26498 31580
rect 26434 31520 26498 31524
rect 26514 31580 26578 31584
rect 26514 31524 26518 31580
rect 26518 31524 26574 31580
rect 26574 31524 26578 31580
rect 26514 31520 26578 31524
rect 34715 31580 34779 31584
rect 34715 31524 34719 31580
rect 34719 31524 34775 31580
rect 34775 31524 34779 31580
rect 34715 31520 34779 31524
rect 34795 31580 34859 31584
rect 34795 31524 34799 31580
rect 34799 31524 34855 31580
rect 34855 31524 34859 31580
rect 34795 31520 34859 31524
rect 34875 31580 34939 31584
rect 34875 31524 34879 31580
rect 34879 31524 34935 31580
rect 34935 31524 34939 31580
rect 34875 31520 34939 31524
rect 34955 31580 35019 31584
rect 34955 31524 34959 31580
rect 34959 31524 35015 31580
rect 35015 31524 35019 31580
rect 34955 31520 35019 31524
rect 5172 31036 5236 31040
rect 5172 30980 5176 31036
rect 5176 30980 5232 31036
rect 5232 30980 5236 31036
rect 5172 30976 5236 30980
rect 5252 31036 5316 31040
rect 5252 30980 5256 31036
rect 5256 30980 5312 31036
rect 5312 30980 5316 31036
rect 5252 30976 5316 30980
rect 5332 31036 5396 31040
rect 5332 30980 5336 31036
rect 5336 30980 5392 31036
rect 5392 30980 5396 31036
rect 5332 30976 5396 30980
rect 5412 31036 5476 31040
rect 5412 30980 5416 31036
rect 5416 30980 5472 31036
rect 5472 30980 5476 31036
rect 5412 30976 5476 30980
rect 13613 31036 13677 31040
rect 13613 30980 13617 31036
rect 13617 30980 13673 31036
rect 13673 30980 13677 31036
rect 13613 30976 13677 30980
rect 13693 31036 13757 31040
rect 13693 30980 13697 31036
rect 13697 30980 13753 31036
rect 13753 30980 13757 31036
rect 13693 30976 13757 30980
rect 13773 31036 13837 31040
rect 13773 30980 13777 31036
rect 13777 30980 13833 31036
rect 13833 30980 13837 31036
rect 13773 30976 13837 30980
rect 13853 31036 13917 31040
rect 13853 30980 13857 31036
rect 13857 30980 13913 31036
rect 13913 30980 13917 31036
rect 13853 30976 13917 30980
rect 22054 31036 22118 31040
rect 22054 30980 22058 31036
rect 22058 30980 22114 31036
rect 22114 30980 22118 31036
rect 22054 30976 22118 30980
rect 22134 31036 22198 31040
rect 22134 30980 22138 31036
rect 22138 30980 22194 31036
rect 22194 30980 22198 31036
rect 22134 30976 22198 30980
rect 22214 31036 22278 31040
rect 22214 30980 22218 31036
rect 22218 30980 22274 31036
rect 22274 30980 22278 31036
rect 22214 30976 22278 30980
rect 22294 31036 22358 31040
rect 22294 30980 22298 31036
rect 22298 30980 22354 31036
rect 22354 30980 22358 31036
rect 22294 30976 22358 30980
rect 30495 31036 30559 31040
rect 30495 30980 30499 31036
rect 30499 30980 30555 31036
rect 30555 30980 30559 31036
rect 30495 30976 30559 30980
rect 30575 31036 30639 31040
rect 30575 30980 30579 31036
rect 30579 30980 30635 31036
rect 30635 30980 30639 31036
rect 30575 30976 30639 30980
rect 30655 31036 30719 31040
rect 30655 30980 30659 31036
rect 30659 30980 30715 31036
rect 30715 30980 30719 31036
rect 30655 30976 30719 30980
rect 30735 31036 30799 31040
rect 30735 30980 30739 31036
rect 30739 30980 30795 31036
rect 30795 30980 30799 31036
rect 30735 30976 30799 30980
rect 9392 30492 9456 30496
rect 9392 30436 9396 30492
rect 9396 30436 9452 30492
rect 9452 30436 9456 30492
rect 9392 30432 9456 30436
rect 9472 30492 9536 30496
rect 9472 30436 9476 30492
rect 9476 30436 9532 30492
rect 9532 30436 9536 30492
rect 9472 30432 9536 30436
rect 9552 30492 9616 30496
rect 9552 30436 9556 30492
rect 9556 30436 9612 30492
rect 9612 30436 9616 30492
rect 9552 30432 9616 30436
rect 9632 30492 9696 30496
rect 9632 30436 9636 30492
rect 9636 30436 9692 30492
rect 9692 30436 9696 30492
rect 9632 30432 9696 30436
rect 17833 30492 17897 30496
rect 17833 30436 17837 30492
rect 17837 30436 17893 30492
rect 17893 30436 17897 30492
rect 17833 30432 17897 30436
rect 17913 30492 17977 30496
rect 17913 30436 17917 30492
rect 17917 30436 17973 30492
rect 17973 30436 17977 30492
rect 17913 30432 17977 30436
rect 17993 30492 18057 30496
rect 17993 30436 17997 30492
rect 17997 30436 18053 30492
rect 18053 30436 18057 30492
rect 17993 30432 18057 30436
rect 18073 30492 18137 30496
rect 18073 30436 18077 30492
rect 18077 30436 18133 30492
rect 18133 30436 18137 30492
rect 18073 30432 18137 30436
rect 26274 30492 26338 30496
rect 26274 30436 26278 30492
rect 26278 30436 26334 30492
rect 26334 30436 26338 30492
rect 26274 30432 26338 30436
rect 26354 30492 26418 30496
rect 26354 30436 26358 30492
rect 26358 30436 26414 30492
rect 26414 30436 26418 30492
rect 26354 30432 26418 30436
rect 26434 30492 26498 30496
rect 26434 30436 26438 30492
rect 26438 30436 26494 30492
rect 26494 30436 26498 30492
rect 26434 30432 26498 30436
rect 26514 30492 26578 30496
rect 26514 30436 26518 30492
rect 26518 30436 26574 30492
rect 26574 30436 26578 30492
rect 26514 30432 26578 30436
rect 34715 30492 34779 30496
rect 34715 30436 34719 30492
rect 34719 30436 34775 30492
rect 34775 30436 34779 30492
rect 34715 30432 34779 30436
rect 34795 30492 34859 30496
rect 34795 30436 34799 30492
rect 34799 30436 34855 30492
rect 34855 30436 34859 30492
rect 34795 30432 34859 30436
rect 34875 30492 34939 30496
rect 34875 30436 34879 30492
rect 34879 30436 34935 30492
rect 34935 30436 34939 30492
rect 34875 30432 34939 30436
rect 34955 30492 35019 30496
rect 34955 30436 34959 30492
rect 34959 30436 35015 30492
rect 35015 30436 35019 30492
rect 34955 30432 35019 30436
rect 5172 29948 5236 29952
rect 5172 29892 5176 29948
rect 5176 29892 5232 29948
rect 5232 29892 5236 29948
rect 5172 29888 5236 29892
rect 5252 29948 5316 29952
rect 5252 29892 5256 29948
rect 5256 29892 5312 29948
rect 5312 29892 5316 29948
rect 5252 29888 5316 29892
rect 5332 29948 5396 29952
rect 5332 29892 5336 29948
rect 5336 29892 5392 29948
rect 5392 29892 5396 29948
rect 5332 29888 5396 29892
rect 5412 29948 5476 29952
rect 5412 29892 5416 29948
rect 5416 29892 5472 29948
rect 5472 29892 5476 29948
rect 5412 29888 5476 29892
rect 13613 29948 13677 29952
rect 13613 29892 13617 29948
rect 13617 29892 13673 29948
rect 13673 29892 13677 29948
rect 13613 29888 13677 29892
rect 13693 29948 13757 29952
rect 13693 29892 13697 29948
rect 13697 29892 13753 29948
rect 13753 29892 13757 29948
rect 13693 29888 13757 29892
rect 13773 29948 13837 29952
rect 13773 29892 13777 29948
rect 13777 29892 13833 29948
rect 13833 29892 13837 29948
rect 13773 29888 13837 29892
rect 13853 29948 13917 29952
rect 13853 29892 13857 29948
rect 13857 29892 13913 29948
rect 13913 29892 13917 29948
rect 13853 29888 13917 29892
rect 22054 29948 22118 29952
rect 22054 29892 22058 29948
rect 22058 29892 22114 29948
rect 22114 29892 22118 29948
rect 22054 29888 22118 29892
rect 22134 29948 22198 29952
rect 22134 29892 22138 29948
rect 22138 29892 22194 29948
rect 22194 29892 22198 29948
rect 22134 29888 22198 29892
rect 22214 29948 22278 29952
rect 22214 29892 22218 29948
rect 22218 29892 22274 29948
rect 22274 29892 22278 29948
rect 22214 29888 22278 29892
rect 22294 29948 22358 29952
rect 22294 29892 22298 29948
rect 22298 29892 22354 29948
rect 22354 29892 22358 29948
rect 22294 29888 22358 29892
rect 30495 29948 30559 29952
rect 30495 29892 30499 29948
rect 30499 29892 30555 29948
rect 30555 29892 30559 29948
rect 30495 29888 30559 29892
rect 30575 29948 30639 29952
rect 30575 29892 30579 29948
rect 30579 29892 30635 29948
rect 30635 29892 30639 29948
rect 30575 29888 30639 29892
rect 30655 29948 30719 29952
rect 30655 29892 30659 29948
rect 30659 29892 30715 29948
rect 30715 29892 30719 29948
rect 30655 29888 30719 29892
rect 30735 29948 30799 29952
rect 30735 29892 30739 29948
rect 30739 29892 30795 29948
rect 30795 29892 30799 29948
rect 30735 29888 30799 29892
rect 9392 29404 9456 29408
rect 9392 29348 9396 29404
rect 9396 29348 9452 29404
rect 9452 29348 9456 29404
rect 9392 29344 9456 29348
rect 9472 29404 9536 29408
rect 9472 29348 9476 29404
rect 9476 29348 9532 29404
rect 9532 29348 9536 29404
rect 9472 29344 9536 29348
rect 9552 29404 9616 29408
rect 9552 29348 9556 29404
rect 9556 29348 9612 29404
rect 9612 29348 9616 29404
rect 9552 29344 9616 29348
rect 9632 29404 9696 29408
rect 9632 29348 9636 29404
rect 9636 29348 9692 29404
rect 9692 29348 9696 29404
rect 9632 29344 9696 29348
rect 17833 29404 17897 29408
rect 17833 29348 17837 29404
rect 17837 29348 17893 29404
rect 17893 29348 17897 29404
rect 17833 29344 17897 29348
rect 17913 29404 17977 29408
rect 17913 29348 17917 29404
rect 17917 29348 17973 29404
rect 17973 29348 17977 29404
rect 17913 29344 17977 29348
rect 17993 29404 18057 29408
rect 17993 29348 17997 29404
rect 17997 29348 18053 29404
rect 18053 29348 18057 29404
rect 17993 29344 18057 29348
rect 18073 29404 18137 29408
rect 18073 29348 18077 29404
rect 18077 29348 18133 29404
rect 18133 29348 18137 29404
rect 18073 29344 18137 29348
rect 26274 29404 26338 29408
rect 26274 29348 26278 29404
rect 26278 29348 26334 29404
rect 26334 29348 26338 29404
rect 26274 29344 26338 29348
rect 26354 29404 26418 29408
rect 26354 29348 26358 29404
rect 26358 29348 26414 29404
rect 26414 29348 26418 29404
rect 26354 29344 26418 29348
rect 26434 29404 26498 29408
rect 26434 29348 26438 29404
rect 26438 29348 26494 29404
rect 26494 29348 26498 29404
rect 26434 29344 26498 29348
rect 26514 29404 26578 29408
rect 26514 29348 26518 29404
rect 26518 29348 26574 29404
rect 26574 29348 26578 29404
rect 26514 29344 26578 29348
rect 34715 29404 34779 29408
rect 34715 29348 34719 29404
rect 34719 29348 34775 29404
rect 34775 29348 34779 29404
rect 34715 29344 34779 29348
rect 34795 29404 34859 29408
rect 34795 29348 34799 29404
rect 34799 29348 34855 29404
rect 34855 29348 34859 29404
rect 34795 29344 34859 29348
rect 34875 29404 34939 29408
rect 34875 29348 34879 29404
rect 34879 29348 34935 29404
rect 34935 29348 34939 29404
rect 34875 29344 34939 29348
rect 34955 29404 35019 29408
rect 34955 29348 34959 29404
rect 34959 29348 35015 29404
rect 35015 29348 35019 29404
rect 34955 29344 35019 29348
rect 5172 28860 5236 28864
rect 5172 28804 5176 28860
rect 5176 28804 5232 28860
rect 5232 28804 5236 28860
rect 5172 28800 5236 28804
rect 5252 28860 5316 28864
rect 5252 28804 5256 28860
rect 5256 28804 5312 28860
rect 5312 28804 5316 28860
rect 5252 28800 5316 28804
rect 5332 28860 5396 28864
rect 5332 28804 5336 28860
rect 5336 28804 5392 28860
rect 5392 28804 5396 28860
rect 5332 28800 5396 28804
rect 5412 28860 5476 28864
rect 5412 28804 5416 28860
rect 5416 28804 5472 28860
rect 5472 28804 5476 28860
rect 5412 28800 5476 28804
rect 13613 28860 13677 28864
rect 13613 28804 13617 28860
rect 13617 28804 13673 28860
rect 13673 28804 13677 28860
rect 13613 28800 13677 28804
rect 13693 28860 13757 28864
rect 13693 28804 13697 28860
rect 13697 28804 13753 28860
rect 13753 28804 13757 28860
rect 13693 28800 13757 28804
rect 13773 28860 13837 28864
rect 13773 28804 13777 28860
rect 13777 28804 13833 28860
rect 13833 28804 13837 28860
rect 13773 28800 13837 28804
rect 13853 28860 13917 28864
rect 13853 28804 13857 28860
rect 13857 28804 13913 28860
rect 13913 28804 13917 28860
rect 13853 28800 13917 28804
rect 22054 28860 22118 28864
rect 22054 28804 22058 28860
rect 22058 28804 22114 28860
rect 22114 28804 22118 28860
rect 22054 28800 22118 28804
rect 22134 28860 22198 28864
rect 22134 28804 22138 28860
rect 22138 28804 22194 28860
rect 22194 28804 22198 28860
rect 22134 28800 22198 28804
rect 22214 28860 22278 28864
rect 22214 28804 22218 28860
rect 22218 28804 22274 28860
rect 22274 28804 22278 28860
rect 22214 28800 22278 28804
rect 22294 28860 22358 28864
rect 22294 28804 22298 28860
rect 22298 28804 22354 28860
rect 22354 28804 22358 28860
rect 22294 28800 22358 28804
rect 30495 28860 30559 28864
rect 30495 28804 30499 28860
rect 30499 28804 30555 28860
rect 30555 28804 30559 28860
rect 30495 28800 30559 28804
rect 30575 28860 30639 28864
rect 30575 28804 30579 28860
rect 30579 28804 30635 28860
rect 30635 28804 30639 28860
rect 30575 28800 30639 28804
rect 30655 28860 30719 28864
rect 30655 28804 30659 28860
rect 30659 28804 30715 28860
rect 30715 28804 30719 28860
rect 30655 28800 30719 28804
rect 30735 28860 30799 28864
rect 30735 28804 30739 28860
rect 30739 28804 30795 28860
rect 30795 28804 30799 28860
rect 30735 28800 30799 28804
rect 9392 28316 9456 28320
rect 9392 28260 9396 28316
rect 9396 28260 9452 28316
rect 9452 28260 9456 28316
rect 9392 28256 9456 28260
rect 9472 28316 9536 28320
rect 9472 28260 9476 28316
rect 9476 28260 9532 28316
rect 9532 28260 9536 28316
rect 9472 28256 9536 28260
rect 9552 28316 9616 28320
rect 9552 28260 9556 28316
rect 9556 28260 9612 28316
rect 9612 28260 9616 28316
rect 9552 28256 9616 28260
rect 9632 28316 9696 28320
rect 9632 28260 9636 28316
rect 9636 28260 9692 28316
rect 9692 28260 9696 28316
rect 9632 28256 9696 28260
rect 17833 28316 17897 28320
rect 17833 28260 17837 28316
rect 17837 28260 17893 28316
rect 17893 28260 17897 28316
rect 17833 28256 17897 28260
rect 17913 28316 17977 28320
rect 17913 28260 17917 28316
rect 17917 28260 17973 28316
rect 17973 28260 17977 28316
rect 17913 28256 17977 28260
rect 17993 28316 18057 28320
rect 17993 28260 17997 28316
rect 17997 28260 18053 28316
rect 18053 28260 18057 28316
rect 17993 28256 18057 28260
rect 18073 28316 18137 28320
rect 18073 28260 18077 28316
rect 18077 28260 18133 28316
rect 18133 28260 18137 28316
rect 18073 28256 18137 28260
rect 26274 28316 26338 28320
rect 26274 28260 26278 28316
rect 26278 28260 26334 28316
rect 26334 28260 26338 28316
rect 26274 28256 26338 28260
rect 26354 28316 26418 28320
rect 26354 28260 26358 28316
rect 26358 28260 26414 28316
rect 26414 28260 26418 28316
rect 26354 28256 26418 28260
rect 26434 28316 26498 28320
rect 26434 28260 26438 28316
rect 26438 28260 26494 28316
rect 26494 28260 26498 28316
rect 26434 28256 26498 28260
rect 26514 28316 26578 28320
rect 26514 28260 26518 28316
rect 26518 28260 26574 28316
rect 26574 28260 26578 28316
rect 26514 28256 26578 28260
rect 34715 28316 34779 28320
rect 34715 28260 34719 28316
rect 34719 28260 34775 28316
rect 34775 28260 34779 28316
rect 34715 28256 34779 28260
rect 34795 28316 34859 28320
rect 34795 28260 34799 28316
rect 34799 28260 34855 28316
rect 34855 28260 34859 28316
rect 34795 28256 34859 28260
rect 34875 28316 34939 28320
rect 34875 28260 34879 28316
rect 34879 28260 34935 28316
rect 34935 28260 34939 28316
rect 34875 28256 34939 28260
rect 34955 28316 35019 28320
rect 34955 28260 34959 28316
rect 34959 28260 35015 28316
rect 35015 28260 35019 28316
rect 34955 28256 35019 28260
rect 5172 27772 5236 27776
rect 5172 27716 5176 27772
rect 5176 27716 5232 27772
rect 5232 27716 5236 27772
rect 5172 27712 5236 27716
rect 5252 27772 5316 27776
rect 5252 27716 5256 27772
rect 5256 27716 5312 27772
rect 5312 27716 5316 27772
rect 5252 27712 5316 27716
rect 5332 27772 5396 27776
rect 5332 27716 5336 27772
rect 5336 27716 5392 27772
rect 5392 27716 5396 27772
rect 5332 27712 5396 27716
rect 5412 27772 5476 27776
rect 5412 27716 5416 27772
rect 5416 27716 5472 27772
rect 5472 27716 5476 27772
rect 5412 27712 5476 27716
rect 13613 27772 13677 27776
rect 13613 27716 13617 27772
rect 13617 27716 13673 27772
rect 13673 27716 13677 27772
rect 13613 27712 13677 27716
rect 13693 27772 13757 27776
rect 13693 27716 13697 27772
rect 13697 27716 13753 27772
rect 13753 27716 13757 27772
rect 13693 27712 13757 27716
rect 13773 27772 13837 27776
rect 13773 27716 13777 27772
rect 13777 27716 13833 27772
rect 13833 27716 13837 27772
rect 13773 27712 13837 27716
rect 13853 27772 13917 27776
rect 13853 27716 13857 27772
rect 13857 27716 13913 27772
rect 13913 27716 13917 27772
rect 13853 27712 13917 27716
rect 22054 27772 22118 27776
rect 22054 27716 22058 27772
rect 22058 27716 22114 27772
rect 22114 27716 22118 27772
rect 22054 27712 22118 27716
rect 22134 27772 22198 27776
rect 22134 27716 22138 27772
rect 22138 27716 22194 27772
rect 22194 27716 22198 27772
rect 22134 27712 22198 27716
rect 22214 27772 22278 27776
rect 22214 27716 22218 27772
rect 22218 27716 22274 27772
rect 22274 27716 22278 27772
rect 22214 27712 22278 27716
rect 22294 27772 22358 27776
rect 22294 27716 22298 27772
rect 22298 27716 22354 27772
rect 22354 27716 22358 27772
rect 22294 27712 22358 27716
rect 30495 27772 30559 27776
rect 30495 27716 30499 27772
rect 30499 27716 30555 27772
rect 30555 27716 30559 27772
rect 30495 27712 30559 27716
rect 30575 27772 30639 27776
rect 30575 27716 30579 27772
rect 30579 27716 30635 27772
rect 30635 27716 30639 27772
rect 30575 27712 30639 27716
rect 30655 27772 30719 27776
rect 30655 27716 30659 27772
rect 30659 27716 30715 27772
rect 30715 27716 30719 27772
rect 30655 27712 30719 27716
rect 30735 27772 30799 27776
rect 30735 27716 30739 27772
rect 30739 27716 30795 27772
rect 30795 27716 30799 27772
rect 30735 27712 30799 27716
rect 9392 27228 9456 27232
rect 9392 27172 9396 27228
rect 9396 27172 9452 27228
rect 9452 27172 9456 27228
rect 9392 27168 9456 27172
rect 9472 27228 9536 27232
rect 9472 27172 9476 27228
rect 9476 27172 9532 27228
rect 9532 27172 9536 27228
rect 9472 27168 9536 27172
rect 9552 27228 9616 27232
rect 9552 27172 9556 27228
rect 9556 27172 9612 27228
rect 9612 27172 9616 27228
rect 9552 27168 9616 27172
rect 9632 27228 9696 27232
rect 9632 27172 9636 27228
rect 9636 27172 9692 27228
rect 9692 27172 9696 27228
rect 9632 27168 9696 27172
rect 17833 27228 17897 27232
rect 17833 27172 17837 27228
rect 17837 27172 17893 27228
rect 17893 27172 17897 27228
rect 17833 27168 17897 27172
rect 17913 27228 17977 27232
rect 17913 27172 17917 27228
rect 17917 27172 17973 27228
rect 17973 27172 17977 27228
rect 17913 27168 17977 27172
rect 17993 27228 18057 27232
rect 17993 27172 17997 27228
rect 17997 27172 18053 27228
rect 18053 27172 18057 27228
rect 17993 27168 18057 27172
rect 18073 27228 18137 27232
rect 18073 27172 18077 27228
rect 18077 27172 18133 27228
rect 18133 27172 18137 27228
rect 18073 27168 18137 27172
rect 26274 27228 26338 27232
rect 26274 27172 26278 27228
rect 26278 27172 26334 27228
rect 26334 27172 26338 27228
rect 26274 27168 26338 27172
rect 26354 27228 26418 27232
rect 26354 27172 26358 27228
rect 26358 27172 26414 27228
rect 26414 27172 26418 27228
rect 26354 27168 26418 27172
rect 26434 27228 26498 27232
rect 26434 27172 26438 27228
rect 26438 27172 26494 27228
rect 26494 27172 26498 27228
rect 26434 27168 26498 27172
rect 26514 27228 26578 27232
rect 26514 27172 26518 27228
rect 26518 27172 26574 27228
rect 26574 27172 26578 27228
rect 26514 27168 26578 27172
rect 34715 27228 34779 27232
rect 34715 27172 34719 27228
rect 34719 27172 34775 27228
rect 34775 27172 34779 27228
rect 34715 27168 34779 27172
rect 34795 27228 34859 27232
rect 34795 27172 34799 27228
rect 34799 27172 34855 27228
rect 34855 27172 34859 27228
rect 34795 27168 34859 27172
rect 34875 27228 34939 27232
rect 34875 27172 34879 27228
rect 34879 27172 34935 27228
rect 34935 27172 34939 27228
rect 34875 27168 34939 27172
rect 34955 27228 35019 27232
rect 34955 27172 34959 27228
rect 34959 27172 35015 27228
rect 35015 27172 35019 27228
rect 34955 27168 35019 27172
rect 5172 26684 5236 26688
rect 5172 26628 5176 26684
rect 5176 26628 5232 26684
rect 5232 26628 5236 26684
rect 5172 26624 5236 26628
rect 5252 26684 5316 26688
rect 5252 26628 5256 26684
rect 5256 26628 5312 26684
rect 5312 26628 5316 26684
rect 5252 26624 5316 26628
rect 5332 26684 5396 26688
rect 5332 26628 5336 26684
rect 5336 26628 5392 26684
rect 5392 26628 5396 26684
rect 5332 26624 5396 26628
rect 5412 26684 5476 26688
rect 5412 26628 5416 26684
rect 5416 26628 5472 26684
rect 5472 26628 5476 26684
rect 5412 26624 5476 26628
rect 13613 26684 13677 26688
rect 13613 26628 13617 26684
rect 13617 26628 13673 26684
rect 13673 26628 13677 26684
rect 13613 26624 13677 26628
rect 13693 26684 13757 26688
rect 13693 26628 13697 26684
rect 13697 26628 13753 26684
rect 13753 26628 13757 26684
rect 13693 26624 13757 26628
rect 13773 26684 13837 26688
rect 13773 26628 13777 26684
rect 13777 26628 13833 26684
rect 13833 26628 13837 26684
rect 13773 26624 13837 26628
rect 13853 26684 13917 26688
rect 13853 26628 13857 26684
rect 13857 26628 13913 26684
rect 13913 26628 13917 26684
rect 13853 26624 13917 26628
rect 22054 26684 22118 26688
rect 22054 26628 22058 26684
rect 22058 26628 22114 26684
rect 22114 26628 22118 26684
rect 22054 26624 22118 26628
rect 22134 26684 22198 26688
rect 22134 26628 22138 26684
rect 22138 26628 22194 26684
rect 22194 26628 22198 26684
rect 22134 26624 22198 26628
rect 22214 26684 22278 26688
rect 22214 26628 22218 26684
rect 22218 26628 22274 26684
rect 22274 26628 22278 26684
rect 22214 26624 22278 26628
rect 22294 26684 22358 26688
rect 22294 26628 22298 26684
rect 22298 26628 22354 26684
rect 22354 26628 22358 26684
rect 22294 26624 22358 26628
rect 30495 26684 30559 26688
rect 30495 26628 30499 26684
rect 30499 26628 30555 26684
rect 30555 26628 30559 26684
rect 30495 26624 30559 26628
rect 30575 26684 30639 26688
rect 30575 26628 30579 26684
rect 30579 26628 30635 26684
rect 30635 26628 30639 26684
rect 30575 26624 30639 26628
rect 30655 26684 30719 26688
rect 30655 26628 30659 26684
rect 30659 26628 30715 26684
rect 30715 26628 30719 26684
rect 30655 26624 30719 26628
rect 30735 26684 30799 26688
rect 30735 26628 30739 26684
rect 30739 26628 30795 26684
rect 30795 26628 30799 26684
rect 30735 26624 30799 26628
rect 9392 26140 9456 26144
rect 9392 26084 9396 26140
rect 9396 26084 9452 26140
rect 9452 26084 9456 26140
rect 9392 26080 9456 26084
rect 9472 26140 9536 26144
rect 9472 26084 9476 26140
rect 9476 26084 9532 26140
rect 9532 26084 9536 26140
rect 9472 26080 9536 26084
rect 9552 26140 9616 26144
rect 9552 26084 9556 26140
rect 9556 26084 9612 26140
rect 9612 26084 9616 26140
rect 9552 26080 9616 26084
rect 9632 26140 9696 26144
rect 9632 26084 9636 26140
rect 9636 26084 9692 26140
rect 9692 26084 9696 26140
rect 9632 26080 9696 26084
rect 17833 26140 17897 26144
rect 17833 26084 17837 26140
rect 17837 26084 17893 26140
rect 17893 26084 17897 26140
rect 17833 26080 17897 26084
rect 17913 26140 17977 26144
rect 17913 26084 17917 26140
rect 17917 26084 17973 26140
rect 17973 26084 17977 26140
rect 17913 26080 17977 26084
rect 17993 26140 18057 26144
rect 17993 26084 17997 26140
rect 17997 26084 18053 26140
rect 18053 26084 18057 26140
rect 17993 26080 18057 26084
rect 18073 26140 18137 26144
rect 18073 26084 18077 26140
rect 18077 26084 18133 26140
rect 18133 26084 18137 26140
rect 18073 26080 18137 26084
rect 26274 26140 26338 26144
rect 26274 26084 26278 26140
rect 26278 26084 26334 26140
rect 26334 26084 26338 26140
rect 26274 26080 26338 26084
rect 26354 26140 26418 26144
rect 26354 26084 26358 26140
rect 26358 26084 26414 26140
rect 26414 26084 26418 26140
rect 26354 26080 26418 26084
rect 26434 26140 26498 26144
rect 26434 26084 26438 26140
rect 26438 26084 26494 26140
rect 26494 26084 26498 26140
rect 26434 26080 26498 26084
rect 26514 26140 26578 26144
rect 26514 26084 26518 26140
rect 26518 26084 26574 26140
rect 26574 26084 26578 26140
rect 26514 26080 26578 26084
rect 34715 26140 34779 26144
rect 34715 26084 34719 26140
rect 34719 26084 34775 26140
rect 34775 26084 34779 26140
rect 34715 26080 34779 26084
rect 34795 26140 34859 26144
rect 34795 26084 34799 26140
rect 34799 26084 34855 26140
rect 34855 26084 34859 26140
rect 34795 26080 34859 26084
rect 34875 26140 34939 26144
rect 34875 26084 34879 26140
rect 34879 26084 34935 26140
rect 34935 26084 34939 26140
rect 34875 26080 34939 26084
rect 34955 26140 35019 26144
rect 34955 26084 34959 26140
rect 34959 26084 35015 26140
rect 35015 26084 35019 26140
rect 34955 26080 35019 26084
rect 5172 25596 5236 25600
rect 5172 25540 5176 25596
rect 5176 25540 5232 25596
rect 5232 25540 5236 25596
rect 5172 25536 5236 25540
rect 5252 25596 5316 25600
rect 5252 25540 5256 25596
rect 5256 25540 5312 25596
rect 5312 25540 5316 25596
rect 5252 25536 5316 25540
rect 5332 25596 5396 25600
rect 5332 25540 5336 25596
rect 5336 25540 5392 25596
rect 5392 25540 5396 25596
rect 5332 25536 5396 25540
rect 5412 25596 5476 25600
rect 5412 25540 5416 25596
rect 5416 25540 5472 25596
rect 5472 25540 5476 25596
rect 5412 25536 5476 25540
rect 13613 25596 13677 25600
rect 13613 25540 13617 25596
rect 13617 25540 13673 25596
rect 13673 25540 13677 25596
rect 13613 25536 13677 25540
rect 13693 25596 13757 25600
rect 13693 25540 13697 25596
rect 13697 25540 13753 25596
rect 13753 25540 13757 25596
rect 13693 25536 13757 25540
rect 13773 25596 13837 25600
rect 13773 25540 13777 25596
rect 13777 25540 13833 25596
rect 13833 25540 13837 25596
rect 13773 25536 13837 25540
rect 13853 25596 13917 25600
rect 13853 25540 13857 25596
rect 13857 25540 13913 25596
rect 13913 25540 13917 25596
rect 13853 25536 13917 25540
rect 22054 25596 22118 25600
rect 22054 25540 22058 25596
rect 22058 25540 22114 25596
rect 22114 25540 22118 25596
rect 22054 25536 22118 25540
rect 22134 25596 22198 25600
rect 22134 25540 22138 25596
rect 22138 25540 22194 25596
rect 22194 25540 22198 25596
rect 22134 25536 22198 25540
rect 22214 25596 22278 25600
rect 22214 25540 22218 25596
rect 22218 25540 22274 25596
rect 22274 25540 22278 25596
rect 22214 25536 22278 25540
rect 22294 25596 22358 25600
rect 22294 25540 22298 25596
rect 22298 25540 22354 25596
rect 22354 25540 22358 25596
rect 22294 25536 22358 25540
rect 30495 25596 30559 25600
rect 30495 25540 30499 25596
rect 30499 25540 30555 25596
rect 30555 25540 30559 25596
rect 30495 25536 30559 25540
rect 30575 25596 30639 25600
rect 30575 25540 30579 25596
rect 30579 25540 30635 25596
rect 30635 25540 30639 25596
rect 30575 25536 30639 25540
rect 30655 25596 30719 25600
rect 30655 25540 30659 25596
rect 30659 25540 30715 25596
rect 30715 25540 30719 25596
rect 30655 25536 30719 25540
rect 30735 25596 30799 25600
rect 30735 25540 30739 25596
rect 30739 25540 30795 25596
rect 30795 25540 30799 25596
rect 30735 25536 30799 25540
rect 9392 25052 9456 25056
rect 9392 24996 9396 25052
rect 9396 24996 9452 25052
rect 9452 24996 9456 25052
rect 9392 24992 9456 24996
rect 9472 25052 9536 25056
rect 9472 24996 9476 25052
rect 9476 24996 9532 25052
rect 9532 24996 9536 25052
rect 9472 24992 9536 24996
rect 9552 25052 9616 25056
rect 9552 24996 9556 25052
rect 9556 24996 9612 25052
rect 9612 24996 9616 25052
rect 9552 24992 9616 24996
rect 9632 25052 9696 25056
rect 9632 24996 9636 25052
rect 9636 24996 9692 25052
rect 9692 24996 9696 25052
rect 9632 24992 9696 24996
rect 17833 25052 17897 25056
rect 17833 24996 17837 25052
rect 17837 24996 17893 25052
rect 17893 24996 17897 25052
rect 17833 24992 17897 24996
rect 17913 25052 17977 25056
rect 17913 24996 17917 25052
rect 17917 24996 17973 25052
rect 17973 24996 17977 25052
rect 17913 24992 17977 24996
rect 17993 25052 18057 25056
rect 17993 24996 17997 25052
rect 17997 24996 18053 25052
rect 18053 24996 18057 25052
rect 17993 24992 18057 24996
rect 18073 25052 18137 25056
rect 18073 24996 18077 25052
rect 18077 24996 18133 25052
rect 18133 24996 18137 25052
rect 18073 24992 18137 24996
rect 26274 25052 26338 25056
rect 26274 24996 26278 25052
rect 26278 24996 26334 25052
rect 26334 24996 26338 25052
rect 26274 24992 26338 24996
rect 26354 25052 26418 25056
rect 26354 24996 26358 25052
rect 26358 24996 26414 25052
rect 26414 24996 26418 25052
rect 26354 24992 26418 24996
rect 26434 25052 26498 25056
rect 26434 24996 26438 25052
rect 26438 24996 26494 25052
rect 26494 24996 26498 25052
rect 26434 24992 26498 24996
rect 26514 25052 26578 25056
rect 26514 24996 26518 25052
rect 26518 24996 26574 25052
rect 26574 24996 26578 25052
rect 26514 24992 26578 24996
rect 34715 25052 34779 25056
rect 34715 24996 34719 25052
rect 34719 24996 34775 25052
rect 34775 24996 34779 25052
rect 34715 24992 34779 24996
rect 34795 25052 34859 25056
rect 34795 24996 34799 25052
rect 34799 24996 34855 25052
rect 34855 24996 34859 25052
rect 34795 24992 34859 24996
rect 34875 25052 34939 25056
rect 34875 24996 34879 25052
rect 34879 24996 34935 25052
rect 34935 24996 34939 25052
rect 34875 24992 34939 24996
rect 34955 25052 35019 25056
rect 34955 24996 34959 25052
rect 34959 24996 35015 25052
rect 35015 24996 35019 25052
rect 34955 24992 35019 24996
rect 5172 24508 5236 24512
rect 5172 24452 5176 24508
rect 5176 24452 5232 24508
rect 5232 24452 5236 24508
rect 5172 24448 5236 24452
rect 5252 24508 5316 24512
rect 5252 24452 5256 24508
rect 5256 24452 5312 24508
rect 5312 24452 5316 24508
rect 5252 24448 5316 24452
rect 5332 24508 5396 24512
rect 5332 24452 5336 24508
rect 5336 24452 5392 24508
rect 5392 24452 5396 24508
rect 5332 24448 5396 24452
rect 5412 24508 5476 24512
rect 5412 24452 5416 24508
rect 5416 24452 5472 24508
rect 5472 24452 5476 24508
rect 5412 24448 5476 24452
rect 13613 24508 13677 24512
rect 13613 24452 13617 24508
rect 13617 24452 13673 24508
rect 13673 24452 13677 24508
rect 13613 24448 13677 24452
rect 13693 24508 13757 24512
rect 13693 24452 13697 24508
rect 13697 24452 13753 24508
rect 13753 24452 13757 24508
rect 13693 24448 13757 24452
rect 13773 24508 13837 24512
rect 13773 24452 13777 24508
rect 13777 24452 13833 24508
rect 13833 24452 13837 24508
rect 13773 24448 13837 24452
rect 13853 24508 13917 24512
rect 13853 24452 13857 24508
rect 13857 24452 13913 24508
rect 13913 24452 13917 24508
rect 13853 24448 13917 24452
rect 22054 24508 22118 24512
rect 22054 24452 22058 24508
rect 22058 24452 22114 24508
rect 22114 24452 22118 24508
rect 22054 24448 22118 24452
rect 22134 24508 22198 24512
rect 22134 24452 22138 24508
rect 22138 24452 22194 24508
rect 22194 24452 22198 24508
rect 22134 24448 22198 24452
rect 22214 24508 22278 24512
rect 22214 24452 22218 24508
rect 22218 24452 22274 24508
rect 22274 24452 22278 24508
rect 22214 24448 22278 24452
rect 22294 24508 22358 24512
rect 22294 24452 22298 24508
rect 22298 24452 22354 24508
rect 22354 24452 22358 24508
rect 22294 24448 22358 24452
rect 30495 24508 30559 24512
rect 30495 24452 30499 24508
rect 30499 24452 30555 24508
rect 30555 24452 30559 24508
rect 30495 24448 30559 24452
rect 30575 24508 30639 24512
rect 30575 24452 30579 24508
rect 30579 24452 30635 24508
rect 30635 24452 30639 24508
rect 30575 24448 30639 24452
rect 30655 24508 30719 24512
rect 30655 24452 30659 24508
rect 30659 24452 30715 24508
rect 30715 24452 30719 24508
rect 30655 24448 30719 24452
rect 30735 24508 30799 24512
rect 30735 24452 30739 24508
rect 30739 24452 30795 24508
rect 30795 24452 30799 24508
rect 30735 24448 30799 24452
rect 9392 23964 9456 23968
rect 9392 23908 9396 23964
rect 9396 23908 9452 23964
rect 9452 23908 9456 23964
rect 9392 23904 9456 23908
rect 9472 23964 9536 23968
rect 9472 23908 9476 23964
rect 9476 23908 9532 23964
rect 9532 23908 9536 23964
rect 9472 23904 9536 23908
rect 9552 23964 9616 23968
rect 9552 23908 9556 23964
rect 9556 23908 9612 23964
rect 9612 23908 9616 23964
rect 9552 23904 9616 23908
rect 9632 23964 9696 23968
rect 9632 23908 9636 23964
rect 9636 23908 9692 23964
rect 9692 23908 9696 23964
rect 9632 23904 9696 23908
rect 17833 23964 17897 23968
rect 17833 23908 17837 23964
rect 17837 23908 17893 23964
rect 17893 23908 17897 23964
rect 17833 23904 17897 23908
rect 17913 23964 17977 23968
rect 17913 23908 17917 23964
rect 17917 23908 17973 23964
rect 17973 23908 17977 23964
rect 17913 23904 17977 23908
rect 17993 23964 18057 23968
rect 17993 23908 17997 23964
rect 17997 23908 18053 23964
rect 18053 23908 18057 23964
rect 17993 23904 18057 23908
rect 18073 23964 18137 23968
rect 18073 23908 18077 23964
rect 18077 23908 18133 23964
rect 18133 23908 18137 23964
rect 18073 23904 18137 23908
rect 26274 23964 26338 23968
rect 26274 23908 26278 23964
rect 26278 23908 26334 23964
rect 26334 23908 26338 23964
rect 26274 23904 26338 23908
rect 26354 23964 26418 23968
rect 26354 23908 26358 23964
rect 26358 23908 26414 23964
rect 26414 23908 26418 23964
rect 26354 23904 26418 23908
rect 26434 23964 26498 23968
rect 26434 23908 26438 23964
rect 26438 23908 26494 23964
rect 26494 23908 26498 23964
rect 26434 23904 26498 23908
rect 26514 23964 26578 23968
rect 26514 23908 26518 23964
rect 26518 23908 26574 23964
rect 26574 23908 26578 23964
rect 26514 23904 26578 23908
rect 34715 23964 34779 23968
rect 34715 23908 34719 23964
rect 34719 23908 34775 23964
rect 34775 23908 34779 23964
rect 34715 23904 34779 23908
rect 34795 23964 34859 23968
rect 34795 23908 34799 23964
rect 34799 23908 34855 23964
rect 34855 23908 34859 23964
rect 34795 23904 34859 23908
rect 34875 23964 34939 23968
rect 34875 23908 34879 23964
rect 34879 23908 34935 23964
rect 34935 23908 34939 23964
rect 34875 23904 34939 23908
rect 34955 23964 35019 23968
rect 34955 23908 34959 23964
rect 34959 23908 35015 23964
rect 35015 23908 35019 23964
rect 34955 23904 35019 23908
rect 5172 23420 5236 23424
rect 5172 23364 5176 23420
rect 5176 23364 5232 23420
rect 5232 23364 5236 23420
rect 5172 23360 5236 23364
rect 5252 23420 5316 23424
rect 5252 23364 5256 23420
rect 5256 23364 5312 23420
rect 5312 23364 5316 23420
rect 5252 23360 5316 23364
rect 5332 23420 5396 23424
rect 5332 23364 5336 23420
rect 5336 23364 5392 23420
rect 5392 23364 5396 23420
rect 5332 23360 5396 23364
rect 5412 23420 5476 23424
rect 5412 23364 5416 23420
rect 5416 23364 5472 23420
rect 5472 23364 5476 23420
rect 5412 23360 5476 23364
rect 13613 23420 13677 23424
rect 13613 23364 13617 23420
rect 13617 23364 13673 23420
rect 13673 23364 13677 23420
rect 13613 23360 13677 23364
rect 13693 23420 13757 23424
rect 13693 23364 13697 23420
rect 13697 23364 13753 23420
rect 13753 23364 13757 23420
rect 13693 23360 13757 23364
rect 13773 23420 13837 23424
rect 13773 23364 13777 23420
rect 13777 23364 13833 23420
rect 13833 23364 13837 23420
rect 13773 23360 13837 23364
rect 13853 23420 13917 23424
rect 13853 23364 13857 23420
rect 13857 23364 13913 23420
rect 13913 23364 13917 23420
rect 13853 23360 13917 23364
rect 22054 23420 22118 23424
rect 22054 23364 22058 23420
rect 22058 23364 22114 23420
rect 22114 23364 22118 23420
rect 22054 23360 22118 23364
rect 22134 23420 22198 23424
rect 22134 23364 22138 23420
rect 22138 23364 22194 23420
rect 22194 23364 22198 23420
rect 22134 23360 22198 23364
rect 22214 23420 22278 23424
rect 22214 23364 22218 23420
rect 22218 23364 22274 23420
rect 22274 23364 22278 23420
rect 22214 23360 22278 23364
rect 22294 23420 22358 23424
rect 22294 23364 22298 23420
rect 22298 23364 22354 23420
rect 22354 23364 22358 23420
rect 22294 23360 22358 23364
rect 30495 23420 30559 23424
rect 30495 23364 30499 23420
rect 30499 23364 30555 23420
rect 30555 23364 30559 23420
rect 30495 23360 30559 23364
rect 30575 23420 30639 23424
rect 30575 23364 30579 23420
rect 30579 23364 30635 23420
rect 30635 23364 30639 23420
rect 30575 23360 30639 23364
rect 30655 23420 30719 23424
rect 30655 23364 30659 23420
rect 30659 23364 30715 23420
rect 30715 23364 30719 23420
rect 30655 23360 30719 23364
rect 30735 23420 30799 23424
rect 30735 23364 30739 23420
rect 30739 23364 30795 23420
rect 30795 23364 30799 23420
rect 30735 23360 30799 23364
rect 9392 22876 9456 22880
rect 9392 22820 9396 22876
rect 9396 22820 9452 22876
rect 9452 22820 9456 22876
rect 9392 22816 9456 22820
rect 9472 22876 9536 22880
rect 9472 22820 9476 22876
rect 9476 22820 9532 22876
rect 9532 22820 9536 22876
rect 9472 22816 9536 22820
rect 9552 22876 9616 22880
rect 9552 22820 9556 22876
rect 9556 22820 9612 22876
rect 9612 22820 9616 22876
rect 9552 22816 9616 22820
rect 9632 22876 9696 22880
rect 9632 22820 9636 22876
rect 9636 22820 9692 22876
rect 9692 22820 9696 22876
rect 9632 22816 9696 22820
rect 17833 22876 17897 22880
rect 17833 22820 17837 22876
rect 17837 22820 17893 22876
rect 17893 22820 17897 22876
rect 17833 22816 17897 22820
rect 17913 22876 17977 22880
rect 17913 22820 17917 22876
rect 17917 22820 17973 22876
rect 17973 22820 17977 22876
rect 17913 22816 17977 22820
rect 17993 22876 18057 22880
rect 17993 22820 17997 22876
rect 17997 22820 18053 22876
rect 18053 22820 18057 22876
rect 17993 22816 18057 22820
rect 18073 22876 18137 22880
rect 18073 22820 18077 22876
rect 18077 22820 18133 22876
rect 18133 22820 18137 22876
rect 18073 22816 18137 22820
rect 26274 22876 26338 22880
rect 26274 22820 26278 22876
rect 26278 22820 26334 22876
rect 26334 22820 26338 22876
rect 26274 22816 26338 22820
rect 26354 22876 26418 22880
rect 26354 22820 26358 22876
rect 26358 22820 26414 22876
rect 26414 22820 26418 22876
rect 26354 22816 26418 22820
rect 26434 22876 26498 22880
rect 26434 22820 26438 22876
rect 26438 22820 26494 22876
rect 26494 22820 26498 22876
rect 26434 22816 26498 22820
rect 26514 22876 26578 22880
rect 26514 22820 26518 22876
rect 26518 22820 26574 22876
rect 26574 22820 26578 22876
rect 26514 22816 26578 22820
rect 34715 22876 34779 22880
rect 34715 22820 34719 22876
rect 34719 22820 34775 22876
rect 34775 22820 34779 22876
rect 34715 22816 34779 22820
rect 34795 22876 34859 22880
rect 34795 22820 34799 22876
rect 34799 22820 34855 22876
rect 34855 22820 34859 22876
rect 34795 22816 34859 22820
rect 34875 22876 34939 22880
rect 34875 22820 34879 22876
rect 34879 22820 34935 22876
rect 34935 22820 34939 22876
rect 34875 22816 34939 22820
rect 34955 22876 35019 22880
rect 34955 22820 34959 22876
rect 34959 22820 35015 22876
rect 35015 22820 35019 22876
rect 34955 22816 35019 22820
rect 5172 22332 5236 22336
rect 5172 22276 5176 22332
rect 5176 22276 5232 22332
rect 5232 22276 5236 22332
rect 5172 22272 5236 22276
rect 5252 22332 5316 22336
rect 5252 22276 5256 22332
rect 5256 22276 5312 22332
rect 5312 22276 5316 22332
rect 5252 22272 5316 22276
rect 5332 22332 5396 22336
rect 5332 22276 5336 22332
rect 5336 22276 5392 22332
rect 5392 22276 5396 22332
rect 5332 22272 5396 22276
rect 5412 22332 5476 22336
rect 5412 22276 5416 22332
rect 5416 22276 5472 22332
rect 5472 22276 5476 22332
rect 5412 22272 5476 22276
rect 13613 22332 13677 22336
rect 13613 22276 13617 22332
rect 13617 22276 13673 22332
rect 13673 22276 13677 22332
rect 13613 22272 13677 22276
rect 13693 22332 13757 22336
rect 13693 22276 13697 22332
rect 13697 22276 13753 22332
rect 13753 22276 13757 22332
rect 13693 22272 13757 22276
rect 13773 22332 13837 22336
rect 13773 22276 13777 22332
rect 13777 22276 13833 22332
rect 13833 22276 13837 22332
rect 13773 22272 13837 22276
rect 13853 22332 13917 22336
rect 13853 22276 13857 22332
rect 13857 22276 13913 22332
rect 13913 22276 13917 22332
rect 13853 22272 13917 22276
rect 22054 22332 22118 22336
rect 22054 22276 22058 22332
rect 22058 22276 22114 22332
rect 22114 22276 22118 22332
rect 22054 22272 22118 22276
rect 22134 22332 22198 22336
rect 22134 22276 22138 22332
rect 22138 22276 22194 22332
rect 22194 22276 22198 22332
rect 22134 22272 22198 22276
rect 22214 22332 22278 22336
rect 22214 22276 22218 22332
rect 22218 22276 22274 22332
rect 22274 22276 22278 22332
rect 22214 22272 22278 22276
rect 22294 22332 22358 22336
rect 22294 22276 22298 22332
rect 22298 22276 22354 22332
rect 22354 22276 22358 22332
rect 22294 22272 22358 22276
rect 30495 22332 30559 22336
rect 30495 22276 30499 22332
rect 30499 22276 30555 22332
rect 30555 22276 30559 22332
rect 30495 22272 30559 22276
rect 30575 22332 30639 22336
rect 30575 22276 30579 22332
rect 30579 22276 30635 22332
rect 30635 22276 30639 22332
rect 30575 22272 30639 22276
rect 30655 22332 30719 22336
rect 30655 22276 30659 22332
rect 30659 22276 30715 22332
rect 30715 22276 30719 22332
rect 30655 22272 30719 22276
rect 30735 22332 30799 22336
rect 30735 22276 30739 22332
rect 30739 22276 30795 22332
rect 30795 22276 30799 22332
rect 30735 22272 30799 22276
rect 9392 21788 9456 21792
rect 9392 21732 9396 21788
rect 9396 21732 9452 21788
rect 9452 21732 9456 21788
rect 9392 21728 9456 21732
rect 9472 21788 9536 21792
rect 9472 21732 9476 21788
rect 9476 21732 9532 21788
rect 9532 21732 9536 21788
rect 9472 21728 9536 21732
rect 9552 21788 9616 21792
rect 9552 21732 9556 21788
rect 9556 21732 9612 21788
rect 9612 21732 9616 21788
rect 9552 21728 9616 21732
rect 9632 21788 9696 21792
rect 9632 21732 9636 21788
rect 9636 21732 9692 21788
rect 9692 21732 9696 21788
rect 9632 21728 9696 21732
rect 17833 21788 17897 21792
rect 17833 21732 17837 21788
rect 17837 21732 17893 21788
rect 17893 21732 17897 21788
rect 17833 21728 17897 21732
rect 17913 21788 17977 21792
rect 17913 21732 17917 21788
rect 17917 21732 17973 21788
rect 17973 21732 17977 21788
rect 17913 21728 17977 21732
rect 17993 21788 18057 21792
rect 17993 21732 17997 21788
rect 17997 21732 18053 21788
rect 18053 21732 18057 21788
rect 17993 21728 18057 21732
rect 18073 21788 18137 21792
rect 18073 21732 18077 21788
rect 18077 21732 18133 21788
rect 18133 21732 18137 21788
rect 18073 21728 18137 21732
rect 26274 21788 26338 21792
rect 26274 21732 26278 21788
rect 26278 21732 26334 21788
rect 26334 21732 26338 21788
rect 26274 21728 26338 21732
rect 26354 21788 26418 21792
rect 26354 21732 26358 21788
rect 26358 21732 26414 21788
rect 26414 21732 26418 21788
rect 26354 21728 26418 21732
rect 26434 21788 26498 21792
rect 26434 21732 26438 21788
rect 26438 21732 26494 21788
rect 26494 21732 26498 21788
rect 26434 21728 26498 21732
rect 26514 21788 26578 21792
rect 26514 21732 26518 21788
rect 26518 21732 26574 21788
rect 26574 21732 26578 21788
rect 26514 21728 26578 21732
rect 34715 21788 34779 21792
rect 34715 21732 34719 21788
rect 34719 21732 34775 21788
rect 34775 21732 34779 21788
rect 34715 21728 34779 21732
rect 34795 21788 34859 21792
rect 34795 21732 34799 21788
rect 34799 21732 34855 21788
rect 34855 21732 34859 21788
rect 34795 21728 34859 21732
rect 34875 21788 34939 21792
rect 34875 21732 34879 21788
rect 34879 21732 34935 21788
rect 34935 21732 34939 21788
rect 34875 21728 34939 21732
rect 34955 21788 35019 21792
rect 34955 21732 34959 21788
rect 34959 21732 35015 21788
rect 35015 21732 35019 21788
rect 34955 21728 35019 21732
rect 5172 21244 5236 21248
rect 5172 21188 5176 21244
rect 5176 21188 5232 21244
rect 5232 21188 5236 21244
rect 5172 21184 5236 21188
rect 5252 21244 5316 21248
rect 5252 21188 5256 21244
rect 5256 21188 5312 21244
rect 5312 21188 5316 21244
rect 5252 21184 5316 21188
rect 5332 21244 5396 21248
rect 5332 21188 5336 21244
rect 5336 21188 5392 21244
rect 5392 21188 5396 21244
rect 5332 21184 5396 21188
rect 5412 21244 5476 21248
rect 5412 21188 5416 21244
rect 5416 21188 5472 21244
rect 5472 21188 5476 21244
rect 5412 21184 5476 21188
rect 13613 21244 13677 21248
rect 13613 21188 13617 21244
rect 13617 21188 13673 21244
rect 13673 21188 13677 21244
rect 13613 21184 13677 21188
rect 13693 21244 13757 21248
rect 13693 21188 13697 21244
rect 13697 21188 13753 21244
rect 13753 21188 13757 21244
rect 13693 21184 13757 21188
rect 13773 21244 13837 21248
rect 13773 21188 13777 21244
rect 13777 21188 13833 21244
rect 13833 21188 13837 21244
rect 13773 21184 13837 21188
rect 13853 21244 13917 21248
rect 13853 21188 13857 21244
rect 13857 21188 13913 21244
rect 13913 21188 13917 21244
rect 13853 21184 13917 21188
rect 22054 21244 22118 21248
rect 22054 21188 22058 21244
rect 22058 21188 22114 21244
rect 22114 21188 22118 21244
rect 22054 21184 22118 21188
rect 22134 21244 22198 21248
rect 22134 21188 22138 21244
rect 22138 21188 22194 21244
rect 22194 21188 22198 21244
rect 22134 21184 22198 21188
rect 22214 21244 22278 21248
rect 22214 21188 22218 21244
rect 22218 21188 22274 21244
rect 22274 21188 22278 21244
rect 22214 21184 22278 21188
rect 22294 21244 22358 21248
rect 22294 21188 22298 21244
rect 22298 21188 22354 21244
rect 22354 21188 22358 21244
rect 22294 21184 22358 21188
rect 30495 21244 30559 21248
rect 30495 21188 30499 21244
rect 30499 21188 30555 21244
rect 30555 21188 30559 21244
rect 30495 21184 30559 21188
rect 30575 21244 30639 21248
rect 30575 21188 30579 21244
rect 30579 21188 30635 21244
rect 30635 21188 30639 21244
rect 30575 21184 30639 21188
rect 30655 21244 30719 21248
rect 30655 21188 30659 21244
rect 30659 21188 30715 21244
rect 30715 21188 30719 21244
rect 30655 21184 30719 21188
rect 30735 21244 30799 21248
rect 30735 21188 30739 21244
rect 30739 21188 30795 21244
rect 30795 21188 30799 21244
rect 30735 21184 30799 21188
rect 9392 20700 9456 20704
rect 9392 20644 9396 20700
rect 9396 20644 9452 20700
rect 9452 20644 9456 20700
rect 9392 20640 9456 20644
rect 9472 20700 9536 20704
rect 9472 20644 9476 20700
rect 9476 20644 9532 20700
rect 9532 20644 9536 20700
rect 9472 20640 9536 20644
rect 9552 20700 9616 20704
rect 9552 20644 9556 20700
rect 9556 20644 9612 20700
rect 9612 20644 9616 20700
rect 9552 20640 9616 20644
rect 9632 20700 9696 20704
rect 9632 20644 9636 20700
rect 9636 20644 9692 20700
rect 9692 20644 9696 20700
rect 9632 20640 9696 20644
rect 17833 20700 17897 20704
rect 17833 20644 17837 20700
rect 17837 20644 17893 20700
rect 17893 20644 17897 20700
rect 17833 20640 17897 20644
rect 17913 20700 17977 20704
rect 17913 20644 17917 20700
rect 17917 20644 17973 20700
rect 17973 20644 17977 20700
rect 17913 20640 17977 20644
rect 17993 20700 18057 20704
rect 17993 20644 17997 20700
rect 17997 20644 18053 20700
rect 18053 20644 18057 20700
rect 17993 20640 18057 20644
rect 18073 20700 18137 20704
rect 18073 20644 18077 20700
rect 18077 20644 18133 20700
rect 18133 20644 18137 20700
rect 18073 20640 18137 20644
rect 26274 20700 26338 20704
rect 26274 20644 26278 20700
rect 26278 20644 26334 20700
rect 26334 20644 26338 20700
rect 26274 20640 26338 20644
rect 26354 20700 26418 20704
rect 26354 20644 26358 20700
rect 26358 20644 26414 20700
rect 26414 20644 26418 20700
rect 26354 20640 26418 20644
rect 26434 20700 26498 20704
rect 26434 20644 26438 20700
rect 26438 20644 26494 20700
rect 26494 20644 26498 20700
rect 26434 20640 26498 20644
rect 26514 20700 26578 20704
rect 26514 20644 26518 20700
rect 26518 20644 26574 20700
rect 26574 20644 26578 20700
rect 26514 20640 26578 20644
rect 34715 20700 34779 20704
rect 34715 20644 34719 20700
rect 34719 20644 34775 20700
rect 34775 20644 34779 20700
rect 34715 20640 34779 20644
rect 34795 20700 34859 20704
rect 34795 20644 34799 20700
rect 34799 20644 34855 20700
rect 34855 20644 34859 20700
rect 34795 20640 34859 20644
rect 34875 20700 34939 20704
rect 34875 20644 34879 20700
rect 34879 20644 34935 20700
rect 34935 20644 34939 20700
rect 34875 20640 34939 20644
rect 34955 20700 35019 20704
rect 34955 20644 34959 20700
rect 34959 20644 35015 20700
rect 35015 20644 35019 20700
rect 34955 20640 35019 20644
rect 5172 20156 5236 20160
rect 5172 20100 5176 20156
rect 5176 20100 5232 20156
rect 5232 20100 5236 20156
rect 5172 20096 5236 20100
rect 5252 20156 5316 20160
rect 5252 20100 5256 20156
rect 5256 20100 5312 20156
rect 5312 20100 5316 20156
rect 5252 20096 5316 20100
rect 5332 20156 5396 20160
rect 5332 20100 5336 20156
rect 5336 20100 5392 20156
rect 5392 20100 5396 20156
rect 5332 20096 5396 20100
rect 5412 20156 5476 20160
rect 5412 20100 5416 20156
rect 5416 20100 5472 20156
rect 5472 20100 5476 20156
rect 5412 20096 5476 20100
rect 13613 20156 13677 20160
rect 13613 20100 13617 20156
rect 13617 20100 13673 20156
rect 13673 20100 13677 20156
rect 13613 20096 13677 20100
rect 13693 20156 13757 20160
rect 13693 20100 13697 20156
rect 13697 20100 13753 20156
rect 13753 20100 13757 20156
rect 13693 20096 13757 20100
rect 13773 20156 13837 20160
rect 13773 20100 13777 20156
rect 13777 20100 13833 20156
rect 13833 20100 13837 20156
rect 13773 20096 13837 20100
rect 13853 20156 13917 20160
rect 13853 20100 13857 20156
rect 13857 20100 13913 20156
rect 13913 20100 13917 20156
rect 13853 20096 13917 20100
rect 22054 20156 22118 20160
rect 22054 20100 22058 20156
rect 22058 20100 22114 20156
rect 22114 20100 22118 20156
rect 22054 20096 22118 20100
rect 22134 20156 22198 20160
rect 22134 20100 22138 20156
rect 22138 20100 22194 20156
rect 22194 20100 22198 20156
rect 22134 20096 22198 20100
rect 22214 20156 22278 20160
rect 22214 20100 22218 20156
rect 22218 20100 22274 20156
rect 22274 20100 22278 20156
rect 22214 20096 22278 20100
rect 22294 20156 22358 20160
rect 22294 20100 22298 20156
rect 22298 20100 22354 20156
rect 22354 20100 22358 20156
rect 22294 20096 22358 20100
rect 30495 20156 30559 20160
rect 30495 20100 30499 20156
rect 30499 20100 30555 20156
rect 30555 20100 30559 20156
rect 30495 20096 30559 20100
rect 30575 20156 30639 20160
rect 30575 20100 30579 20156
rect 30579 20100 30635 20156
rect 30635 20100 30639 20156
rect 30575 20096 30639 20100
rect 30655 20156 30719 20160
rect 30655 20100 30659 20156
rect 30659 20100 30715 20156
rect 30715 20100 30719 20156
rect 30655 20096 30719 20100
rect 30735 20156 30799 20160
rect 30735 20100 30739 20156
rect 30739 20100 30795 20156
rect 30795 20100 30799 20156
rect 30735 20096 30799 20100
rect 9392 19612 9456 19616
rect 9392 19556 9396 19612
rect 9396 19556 9452 19612
rect 9452 19556 9456 19612
rect 9392 19552 9456 19556
rect 9472 19612 9536 19616
rect 9472 19556 9476 19612
rect 9476 19556 9532 19612
rect 9532 19556 9536 19612
rect 9472 19552 9536 19556
rect 9552 19612 9616 19616
rect 9552 19556 9556 19612
rect 9556 19556 9612 19612
rect 9612 19556 9616 19612
rect 9552 19552 9616 19556
rect 9632 19612 9696 19616
rect 9632 19556 9636 19612
rect 9636 19556 9692 19612
rect 9692 19556 9696 19612
rect 9632 19552 9696 19556
rect 17833 19612 17897 19616
rect 17833 19556 17837 19612
rect 17837 19556 17893 19612
rect 17893 19556 17897 19612
rect 17833 19552 17897 19556
rect 17913 19612 17977 19616
rect 17913 19556 17917 19612
rect 17917 19556 17973 19612
rect 17973 19556 17977 19612
rect 17913 19552 17977 19556
rect 17993 19612 18057 19616
rect 17993 19556 17997 19612
rect 17997 19556 18053 19612
rect 18053 19556 18057 19612
rect 17993 19552 18057 19556
rect 18073 19612 18137 19616
rect 18073 19556 18077 19612
rect 18077 19556 18133 19612
rect 18133 19556 18137 19612
rect 18073 19552 18137 19556
rect 26274 19612 26338 19616
rect 26274 19556 26278 19612
rect 26278 19556 26334 19612
rect 26334 19556 26338 19612
rect 26274 19552 26338 19556
rect 26354 19612 26418 19616
rect 26354 19556 26358 19612
rect 26358 19556 26414 19612
rect 26414 19556 26418 19612
rect 26354 19552 26418 19556
rect 26434 19612 26498 19616
rect 26434 19556 26438 19612
rect 26438 19556 26494 19612
rect 26494 19556 26498 19612
rect 26434 19552 26498 19556
rect 26514 19612 26578 19616
rect 26514 19556 26518 19612
rect 26518 19556 26574 19612
rect 26574 19556 26578 19612
rect 26514 19552 26578 19556
rect 34715 19612 34779 19616
rect 34715 19556 34719 19612
rect 34719 19556 34775 19612
rect 34775 19556 34779 19612
rect 34715 19552 34779 19556
rect 34795 19612 34859 19616
rect 34795 19556 34799 19612
rect 34799 19556 34855 19612
rect 34855 19556 34859 19612
rect 34795 19552 34859 19556
rect 34875 19612 34939 19616
rect 34875 19556 34879 19612
rect 34879 19556 34935 19612
rect 34935 19556 34939 19612
rect 34875 19552 34939 19556
rect 34955 19612 35019 19616
rect 34955 19556 34959 19612
rect 34959 19556 35015 19612
rect 35015 19556 35019 19612
rect 34955 19552 35019 19556
rect 5172 19068 5236 19072
rect 5172 19012 5176 19068
rect 5176 19012 5232 19068
rect 5232 19012 5236 19068
rect 5172 19008 5236 19012
rect 5252 19068 5316 19072
rect 5252 19012 5256 19068
rect 5256 19012 5312 19068
rect 5312 19012 5316 19068
rect 5252 19008 5316 19012
rect 5332 19068 5396 19072
rect 5332 19012 5336 19068
rect 5336 19012 5392 19068
rect 5392 19012 5396 19068
rect 5332 19008 5396 19012
rect 5412 19068 5476 19072
rect 5412 19012 5416 19068
rect 5416 19012 5472 19068
rect 5472 19012 5476 19068
rect 5412 19008 5476 19012
rect 13613 19068 13677 19072
rect 13613 19012 13617 19068
rect 13617 19012 13673 19068
rect 13673 19012 13677 19068
rect 13613 19008 13677 19012
rect 13693 19068 13757 19072
rect 13693 19012 13697 19068
rect 13697 19012 13753 19068
rect 13753 19012 13757 19068
rect 13693 19008 13757 19012
rect 13773 19068 13837 19072
rect 13773 19012 13777 19068
rect 13777 19012 13833 19068
rect 13833 19012 13837 19068
rect 13773 19008 13837 19012
rect 13853 19068 13917 19072
rect 13853 19012 13857 19068
rect 13857 19012 13913 19068
rect 13913 19012 13917 19068
rect 13853 19008 13917 19012
rect 22054 19068 22118 19072
rect 22054 19012 22058 19068
rect 22058 19012 22114 19068
rect 22114 19012 22118 19068
rect 22054 19008 22118 19012
rect 22134 19068 22198 19072
rect 22134 19012 22138 19068
rect 22138 19012 22194 19068
rect 22194 19012 22198 19068
rect 22134 19008 22198 19012
rect 22214 19068 22278 19072
rect 22214 19012 22218 19068
rect 22218 19012 22274 19068
rect 22274 19012 22278 19068
rect 22214 19008 22278 19012
rect 22294 19068 22358 19072
rect 22294 19012 22298 19068
rect 22298 19012 22354 19068
rect 22354 19012 22358 19068
rect 22294 19008 22358 19012
rect 30495 19068 30559 19072
rect 30495 19012 30499 19068
rect 30499 19012 30555 19068
rect 30555 19012 30559 19068
rect 30495 19008 30559 19012
rect 30575 19068 30639 19072
rect 30575 19012 30579 19068
rect 30579 19012 30635 19068
rect 30635 19012 30639 19068
rect 30575 19008 30639 19012
rect 30655 19068 30719 19072
rect 30655 19012 30659 19068
rect 30659 19012 30715 19068
rect 30715 19012 30719 19068
rect 30655 19008 30719 19012
rect 30735 19068 30799 19072
rect 30735 19012 30739 19068
rect 30739 19012 30795 19068
rect 30795 19012 30799 19068
rect 30735 19008 30799 19012
rect 9392 18524 9456 18528
rect 9392 18468 9396 18524
rect 9396 18468 9452 18524
rect 9452 18468 9456 18524
rect 9392 18464 9456 18468
rect 9472 18524 9536 18528
rect 9472 18468 9476 18524
rect 9476 18468 9532 18524
rect 9532 18468 9536 18524
rect 9472 18464 9536 18468
rect 9552 18524 9616 18528
rect 9552 18468 9556 18524
rect 9556 18468 9612 18524
rect 9612 18468 9616 18524
rect 9552 18464 9616 18468
rect 9632 18524 9696 18528
rect 9632 18468 9636 18524
rect 9636 18468 9692 18524
rect 9692 18468 9696 18524
rect 9632 18464 9696 18468
rect 17833 18524 17897 18528
rect 17833 18468 17837 18524
rect 17837 18468 17893 18524
rect 17893 18468 17897 18524
rect 17833 18464 17897 18468
rect 17913 18524 17977 18528
rect 17913 18468 17917 18524
rect 17917 18468 17973 18524
rect 17973 18468 17977 18524
rect 17913 18464 17977 18468
rect 17993 18524 18057 18528
rect 17993 18468 17997 18524
rect 17997 18468 18053 18524
rect 18053 18468 18057 18524
rect 17993 18464 18057 18468
rect 18073 18524 18137 18528
rect 18073 18468 18077 18524
rect 18077 18468 18133 18524
rect 18133 18468 18137 18524
rect 18073 18464 18137 18468
rect 26274 18524 26338 18528
rect 26274 18468 26278 18524
rect 26278 18468 26334 18524
rect 26334 18468 26338 18524
rect 26274 18464 26338 18468
rect 26354 18524 26418 18528
rect 26354 18468 26358 18524
rect 26358 18468 26414 18524
rect 26414 18468 26418 18524
rect 26354 18464 26418 18468
rect 26434 18524 26498 18528
rect 26434 18468 26438 18524
rect 26438 18468 26494 18524
rect 26494 18468 26498 18524
rect 26434 18464 26498 18468
rect 26514 18524 26578 18528
rect 26514 18468 26518 18524
rect 26518 18468 26574 18524
rect 26574 18468 26578 18524
rect 26514 18464 26578 18468
rect 34715 18524 34779 18528
rect 34715 18468 34719 18524
rect 34719 18468 34775 18524
rect 34775 18468 34779 18524
rect 34715 18464 34779 18468
rect 34795 18524 34859 18528
rect 34795 18468 34799 18524
rect 34799 18468 34855 18524
rect 34855 18468 34859 18524
rect 34795 18464 34859 18468
rect 34875 18524 34939 18528
rect 34875 18468 34879 18524
rect 34879 18468 34935 18524
rect 34935 18468 34939 18524
rect 34875 18464 34939 18468
rect 34955 18524 35019 18528
rect 34955 18468 34959 18524
rect 34959 18468 35015 18524
rect 35015 18468 35019 18524
rect 34955 18464 35019 18468
rect 5172 17980 5236 17984
rect 5172 17924 5176 17980
rect 5176 17924 5232 17980
rect 5232 17924 5236 17980
rect 5172 17920 5236 17924
rect 5252 17980 5316 17984
rect 5252 17924 5256 17980
rect 5256 17924 5312 17980
rect 5312 17924 5316 17980
rect 5252 17920 5316 17924
rect 5332 17980 5396 17984
rect 5332 17924 5336 17980
rect 5336 17924 5392 17980
rect 5392 17924 5396 17980
rect 5332 17920 5396 17924
rect 5412 17980 5476 17984
rect 5412 17924 5416 17980
rect 5416 17924 5472 17980
rect 5472 17924 5476 17980
rect 5412 17920 5476 17924
rect 13613 17980 13677 17984
rect 13613 17924 13617 17980
rect 13617 17924 13673 17980
rect 13673 17924 13677 17980
rect 13613 17920 13677 17924
rect 13693 17980 13757 17984
rect 13693 17924 13697 17980
rect 13697 17924 13753 17980
rect 13753 17924 13757 17980
rect 13693 17920 13757 17924
rect 13773 17980 13837 17984
rect 13773 17924 13777 17980
rect 13777 17924 13833 17980
rect 13833 17924 13837 17980
rect 13773 17920 13837 17924
rect 13853 17980 13917 17984
rect 13853 17924 13857 17980
rect 13857 17924 13913 17980
rect 13913 17924 13917 17980
rect 13853 17920 13917 17924
rect 22054 17980 22118 17984
rect 22054 17924 22058 17980
rect 22058 17924 22114 17980
rect 22114 17924 22118 17980
rect 22054 17920 22118 17924
rect 22134 17980 22198 17984
rect 22134 17924 22138 17980
rect 22138 17924 22194 17980
rect 22194 17924 22198 17980
rect 22134 17920 22198 17924
rect 22214 17980 22278 17984
rect 22214 17924 22218 17980
rect 22218 17924 22274 17980
rect 22274 17924 22278 17980
rect 22214 17920 22278 17924
rect 22294 17980 22358 17984
rect 22294 17924 22298 17980
rect 22298 17924 22354 17980
rect 22354 17924 22358 17980
rect 22294 17920 22358 17924
rect 30495 17980 30559 17984
rect 30495 17924 30499 17980
rect 30499 17924 30555 17980
rect 30555 17924 30559 17980
rect 30495 17920 30559 17924
rect 30575 17980 30639 17984
rect 30575 17924 30579 17980
rect 30579 17924 30635 17980
rect 30635 17924 30639 17980
rect 30575 17920 30639 17924
rect 30655 17980 30719 17984
rect 30655 17924 30659 17980
rect 30659 17924 30715 17980
rect 30715 17924 30719 17980
rect 30655 17920 30719 17924
rect 30735 17980 30799 17984
rect 30735 17924 30739 17980
rect 30739 17924 30795 17980
rect 30795 17924 30799 17980
rect 30735 17920 30799 17924
rect 9392 17436 9456 17440
rect 9392 17380 9396 17436
rect 9396 17380 9452 17436
rect 9452 17380 9456 17436
rect 9392 17376 9456 17380
rect 9472 17436 9536 17440
rect 9472 17380 9476 17436
rect 9476 17380 9532 17436
rect 9532 17380 9536 17436
rect 9472 17376 9536 17380
rect 9552 17436 9616 17440
rect 9552 17380 9556 17436
rect 9556 17380 9612 17436
rect 9612 17380 9616 17436
rect 9552 17376 9616 17380
rect 9632 17436 9696 17440
rect 9632 17380 9636 17436
rect 9636 17380 9692 17436
rect 9692 17380 9696 17436
rect 9632 17376 9696 17380
rect 17833 17436 17897 17440
rect 17833 17380 17837 17436
rect 17837 17380 17893 17436
rect 17893 17380 17897 17436
rect 17833 17376 17897 17380
rect 17913 17436 17977 17440
rect 17913 17380 17917 17436
rect 17917 17380 17973 17436
rect 17973 17380 17977 17436
rect 17913 17376 17977 17380
rect 17993 17436 18057 17440
rect 17993 17380 17997 17436
rect 17997 17380 18053 17436
rect 18053 17380 18057 17436
rect 17993 17376 18057 17380
rect 18073 17436 18137 17440
rect 18073 17380 18077 17436
rect 18077 17380 18133 17436
rect 18133 17380 18137 17436
rect 18073 17376 18137 17380
rect 26274 17436 26338 17440
rect 26274 17380 26278 17436
rect 26278 17380 26334 17436
rect 26334 17380 26338 17436
rect 26274 17376 26338 17380
rect 26354 17436 26418 17440
rect 26354 17380 26358 17436
rect 26358 17380 26414 17436
rect 26414 17380 26418 17436
rect 26354 17376 26418 17380
rect 26434 17436 26498 17440
rect 26434 17380 26438 17436
rect 26438 17380 26494 17436
rect 26494 17380 26498 17436
rect 26434 17376 26498 17380
rect 26514 17436 26578 17440
rect 26514 17380 26518 17436
rect 26518 17380 26574 17436
rect 26574 17380 26578 17436
rect 26514 17376 26578 17380
rect 34715 17436 34779 17440
rect 34715 17380 34719 17436
rect 34719 17380 34775 17436
rect 34775 17380 34779 17436
rect 34715 17376 34779 17380
rect 34795 17436 34859 17440
rect 34795 17380 34799 17436
rect 34799 17380 34855 17436
rect 34855 17380 34859 17436
rect 34795 17376 34859 17380
rect 34875 17436 34939 17440
rect 34875 17380 34879 17436
rect 34879 17380 34935 17436
rect 34935 17380 34939 17436
rect 34875 17376 34939 17380
rect 34955 17436 35019 17440
rect 34955 17380 34959 17436
rect 34959 17380 35015 17436
rect 35015 17380 35019 17436
rect 34955 17376 35019 17380
rect 5172 16892 5236 16896
rect 5172 16836 5176 16892
rect 5176 16836 5232 16892
rect 5232 16836 5236 16892
rect 5172 16832 5236 16836
rect 5252 16892 5316 16896
rect 5252 16836 5256 16892
rect 5256 16836 5312 16892
rect 5312 16836 5316 16892
rect 5252 16832 5316 16836
rect 5332 16892 5396 16896
rect 5332 16836 5336 16892
rect 5336 16836 5392 16892
rect 5392 16836 5396 16892
rect 5332 16832 5396 16836
rect 5412 16892 5476 16896
rect 5412 16836 5416 16892
rect 5416 16836 5472 16892
rect 5472 16836 5476 16892
rect 5412 16832 5476 16836
rect 13613 16892 13677 16896
rect 13613 16836 13617 16892
rect 13617 16836 13673 16892
rect 13673 16836 13677 16892
rect 13613 16832 13677 16836
rect 13693 16892 13757 16896
rect 13693 16836 13697 16892
rect 13697 16836 13753 16892
rect 13753 16836 13757 16892
rect 13693 16832 13757 16836
rect 13773 16892 13837 16896
rect 13773 16836 13777 16892
rect 13777 16836 13833 16892
rect 13833 16836 13837 16892
rect 13773 16832 13837 16836
rect 13853 16892 13917 16896
rect 13853 16836 13857 16892
rect 13857 16836 13913 16892
rect 13913 16836 13917 16892
rect 13853 16832 13917 16836
rect 22054 16892 22118 16896
rect 22054 16836 22058 16892
rect 22058 16836 22114 16892
rect 22114 16836 22118 16892
rect 22054 16832 22118 16836
rect 22134 16892 22198 16896
rect 22134 16836 22138 16892
rect 22138 16836 22194 16892
rect 22194 16836 22198 16892
rect 22134 16832 22198 16836
rect 22214 16892 22278 16896
rect 22214 16836 22218 16892
rect 22218 16836 22274 16892
rect 22274 16836 22278 16892
rect 22214 16832 22278 16836
rect 22294 16892 22358 16896
rect 22294 16836 22298 16892
rect 22298 16836 22354 16892
rect 22354 16836 22358 16892
rect 22294 16832 22358 16836
rect 30495 16892 30559 16896
rect 30495 16836 30499 16892
rect 30499 16836 30555 16892
rect 30555 16836 30559 16892
rect 30495 16832 30559 16836
rect 30575 16892 30639 16896
rect 30575 16836 30579 16892
rect 30579 16836 30635 16892
rect 30635 16836 30639 16892
rect 30575 16832 30639 16836
rect 30655 16892 30719 16896
rect 30655 16836 30659 16892
rect 30659 16836 30715 16892
rect 30715 16836 30719 16892
rect 30655 16832 30719 16836
rect 30735 16892 30799 16896
rect 30735 16836 30739 16892
rect 30739 16836 30795 16892
rect 30795 16836 30799 16892
rect 30735 16832 30799 16836
rect 9392 16348 9456 16352
rect 9392 16292 9396 16348
rect 9396 16292 9452 16348
rect 9452 16292 9456 16348
rect 9392 16288 9456 16292
rect 9472 16348 9536 16352
rect 9472 16292 9476 16348
rect 9476 16292 9532 16348
rect 9532 16292 9536 16348
rect 9472 16288 9536 16292
rect 9552 16348 9616 16352
rect 9552 16292 9556 16348
rect 9556 16292 9612 16348
rect 9612 16292 9616 16348
rect 9552 16288 9616 16292
rect 9632 16348 9696 16352
rect 9632 16292 9636 16348
rect 9636 16292 9692 16348
rect 9692 16292 9696 16348
rect 9632 16288 9696 16292
rect 17833 16348 17897 16352
rect 17833 16292 17837 16348
rect 17837 16292 17893 16348
rect 17893 16292 17897 16348
rect 17833 16288 17897 16292
rect 17913 16348 17977 16352
rect 17913 16292 17917 16348
rect 17917 16292 17973 16348
rect 17973 16292 17977 16348
rect 17913 16288 17977 16292
rect 17993 16348 18057 16352
rect 17993 16292 17997 16348
rect 17997 16292 18053 16348
rect 18053 16292 18057 16348
rect 17993 16288 18057 16292
rect 18073 16348 18137 16352
rect 18073 16292 18077 16348
rect 18077 16292 18133 16348
rect 18133 16292 18137 16348
rect 18073 16288 18137 16292
rect 26274 16348 26338 16352
rect 26274 16292 26278 16348
rect 26278 16292 26334 16348
rect 26334 16292 26338 16348
rect 26274 16288 26338 16292
rect 26354 16348 26418 16352
rect 26354 16292 26358 16348
rect 26358 16292 26414 16348
rect 26414 16292 26418 16348
rect 26354 16288 26418 16292
rect 26434 16348 26498 16352
rect 26434 16292 26438 16348
rect 26438 16292 26494 16348
rect 26494 16292 26498 16348
rect 26434 16288 26498 16292
rect 26514 16348 26578 16352
rect 26514 16292 26518 16348
rect 26518 16292 26574 16348
rect 26574 16292 26578 16348
rect 26514 16288 26578 16292
rect 34715 16348 34779 16352
rect 34715 16292 34719 16348
rect 34719 16292 34775 16348
rect 34775 16292 34779 16348
rect 34715 16288 34779 16292
rect 34795 16348 34859 16352
rect 34795 16292 34799 16348
rect 34799 16292 34855 16348
rect 34855 16292 34859 16348
rect 34795 16288 34859 16292
rect 34875 16348 34939 16352
rect 34875 16292 34879 16348
rect 34879 16292 34935 16348
rect 34935 16292 34939 16348
rect 34875 16288 34939 16292
rect 34955 16348 35019 16352
rect 34955 16292 34959 16348
rect 34959 16292 35015 16348
rect 35015 16292 35019 16348
rect 34955 16288 35019 16292
rect 5172 15804 5236 15808
rect 5172 15748 5176 15804
rect 5176 15748 5232 15804
rect 5232 15748 5236 15804
rect 5172 15744 5236 15748
rect 5252 15804 5316 15808
rect 5252 15748 5256 15804
rect 5256 15748 5312 15804
rect 5312 15748 5316 15804
rect 5252 15744 5316 15748
rect 5332 15804 5396 15808
rect 5332 15748 5336 15804
rect 5336 15748 5392 15804
rect 5392 15748 5396 15804
rect 5332 15744 5396 15748
rect 5412 15804 5476 15808
rect 5412 15748 5416 15804
rect 5416 15748 5472 15804
rect 5472 15748 5476 15804
rect 5412 15744 5476 15748
rect 13613 15804 13677 15808
rect 13613 15748 13617 15804
rect 13617 15748 13673 15804
rect 13673 15748 13677 15804
rect 13613 15744 13677 15748
rect 13693 15804 13757 15808
rect 13693 15748 13697 15804
rect 13697 15748 13753 15804
rect 13753 15748 13757 15804
rect 13693 15744 13757 15748
rect 13773 15804 13837 15808
rect 13773 15748 13777 15804
rect 13777 15748 13833 15804
rect 13833 15748 13837 15804
rect 13773 15744 13837 15748
rect 13853 15804 13917 15808
rect 13853 15748 13857 15804
rect 13857 15748 13913 15804
rect 13913 15748 13917 15804
rect 13853 15744 13917 15748
rect 22054 15804 22118 15808
rect 22054 15748 22058 15804
rect 22058 15748 22114 15804
rect 22114 15748 22118 15804
rect 22054 15744 22118 15748
rect 22134 15804 22198 15808
rect 22134 15748 22138 15804
rect 22138 15748 22194 15804
rect 22194 15748 22198 15804
rect 22134 15744 22198 15748
rect 22214 15804 22278 15808
rect 22214 15748 22218 15804
rect 22218 15748 22274 15804
rect 22274 15748 22278 15804
rect 22214 15744 22278 15748
rect 22294 15804 22358 15808
rect 22294 15748 22298 15804
rect 22298 15748 22354 15804
rect 22354 15748 22358 15804
rect 22294 15744 22358 15748
rect 30495 15804 30559 15808
rect 30495 15748 30499 15804
rect 30499 15748 30555 15804
rect 30555 15748 30559 15804
rect 30495 15744 30559 15748
rect 30575 15804 30639 15808
rect 30575 15748 30579 15804
rect 30579 15748 30635 15804
rect 30635 15748 30639 15804
rect 30575 15744 30639 15748
rect 30655 15804 30719 15808
rect 30655 15748 30659 15804
rect 30659 15748 30715 15804
rect 30715 15748 30719 15804
rect 30655 15744 30719 15748
rect 30735 15804 30799 15808
rect 30735 15748 30739 15804
rect 30739 15748 30795 15804
rect 30795 15748 30799 15804
rect 30735 15744 30799 15748
rect 9392 15260 9456 15264
rect 9392 15204 9396 15260
rect 9396 15204 9452 15260
rect 9452 15204 9456 15260
rect 9392 15200 9456 15204
rect 9472 15260 9536 15264
rect 9472 15204 9476 15260
rect 9476 15204 9532 15260
rect 9532 15204 9536 15260
rect 9472 15200 9536 15204
rect 9552 15260 9616 15264
rect 9552 15204 9556 15260
rect 9556 15204 9612 15260
rect 9612 15204 9616 15260
rect 9552 15200 9616 15204
rect 9632 15260 9696 15264
rect 9632 15204 9636 15260
rect 9636 15204 9692 15260
rect 9692 15204 9696 15260
rect 9632 15200 9696 15204
rect 17833 15260 17897 15264
rect 17833 15204 17837 15260
rect 17837 15204 17893 15260
rect 17893 15204 17897 15260
rect 17833 15200 17897 15204
rect 17913 15260 17977 15264
rect 17913 15204 17917 15260
rect 17917 15204 17973 15260
rect 17973 15204 17977 15260
rect 17913 15200 17977 15204
rect 17993 15260 18057 15264
rect 17993 15204 17997 15260
rect 17997 15204 18053 15260
rect 18053 15204 18057 15260
rect 17993 15200 18057 15204
rect 18073 15260 18137 15264
rect 18073 15204 18077 15260
rect 18077 15204 18133 15260
rect 18133 15204 18137 15260
rect 18073 15200 18137 15204
rect 26274 15260 26338 15264
rect 26274 15204 26278 15260
rect 26278 15204 26334 15260
rect 26334 15204 26338 15260
rect 26274 15200 26338 15204
rect 26354 15260 26418 15264
rect 26354 15204 26358 15260
rect 26358 15204 26414 15260
rect 26414 15204 26418 15260
rect 26354 15200 26418 15204
rect 26434 15260 26498 15264
rect 26434 15204 26438 15260
rect 26438 15204 26494 15260
rect 26494 15204 26498 15260
rect 26434 15200 26498 15204
rect 26514 15260 26578 15264
rect 26514 15204 26518 15260
rect 26518 15204 26574 15260
rect 26574 15204 26578 15260
rect 26514 15200 26578 15204
rect 34715 15260 34779 15264
rect 34715 15204 34719 15260
rect 34719 15204 34775 15260
rect 34775 15204 34779 15260
rect 34715 15200 34779 15204
rect 34795 15260 34859 15264
rect 34795 15204 34799 15260
rect 34799 15204 34855 15260
rect 34855 15204 34859 15260
rect 34795 15200 34859 15204
rect 34875 15260 34939 15264
rect 34875 15204 34879 15260
rect 34879 15204 34935 15260
rect 34935 15204 34939 15260
rect 34875 15200 34939 15204
rect 34955 15260 35019 15264
rect 34955 15204 34959 15260
rect 34959 15204 35015 15260
rect 35015 15204 35019 15260
rect 34955 15200 35019 15204
rect 5172 14716 5236 14720
rect 5172 14660 5176 14716
rect 5176 14660 5232 14716
rect 5232 14660 5236 14716
rect 5172 14656 5236 14660
rect 5252 14716 5316 14720
rect 5252 14660 5256 14716
rect 5256 14660 5312 14716
rect 5312 14660 5316 14716
rect 5252 14656 5316 14660
rect 5332 14716 5396 14720
rect 5332 14660 5336 14716
rect 5336 14660 5392 14716
rect 5392 14660 5396 14716
rect 5332 14656 5396 14660
rect 5412 14716 5476 14720
rect 5412 14660 5416 14716
rect 5416 14660 5472 14716
rect 5472 14660 5476 14716
rect 5412 14656 5476 14660
rect 13613 14716 13677 14720
rect 13613 14660 13617 14716
rect 13617 14660 13673 14716
rect 13673 14660 13677 14716
rect 13613 14656 13677 14660
rect 13693 14716 13757 14720
rect 13693 14660 13697 14716
rect 13697 14660 13753 14716
rect 13753 14660 13757 14716
rect 13693 14656 13757 14660
rect 13773 14716 13837 14720
rect 13773 14660 13777 14716
rect 13777 14660 13833 14716
rect 13833 14660 13837 14716
rect 13773 14656 13837 14660
rect 13853 14716 13917 14720
rect 13853 14660 13857 14716
rect 13857 14660 13913 14716
rect 13913 14660 13917 14716
rect 13853 14656 13917 14660
rect 22054 14716 22118 14720
rect 22054 14660 22058 14716
rect 22058 14660 22114 14716
rect 22114 14660 22118 14716
rect 22054 14656 22118 14660
rect 22134 14716 22198 14720
rect 22134 14660 22138 14716
rect 22138 14660 22194 14716
rect 22194 14660 22198 14716
rect 22134 14656 22198 14660
rect 22214 14716 22278 14720
rect 22214 14660 22218 14716
rect 22218 14660 22274 14716
rect 22274 14660 22278 14716
rect 22214 14656 22278 14660
rect 22294 14716 22358 14720
rect 22294 14660 22298 14716
rect 22298 14660 22354 14716
rect 22354 14660 22358 14716
rect 22294 14656 22358 14660
rect 30495 14716 30559 14720
rect 30495 14660 30499 14716
rect 30499 14660 30555 14716
rect 30555 14660 30559 14716
rect 30495 14656 30559 14660
rect 30575 14716 30639 14720
rect 30575 14660 30579 14716
rect 30579 14660 30635 14716
rect 30635 14660 30639 14716
rect 30575 14656 30639 14660
rect 30655 14716 30719 14720
rect 30655 14660 30659 14716
rect 30659 14660 30715 14716
rect 30715 14660 30719 14716
rect 30655 14656 30719 14660
rect 30735 14716 30799 14720
rect 30735 14660 30739 14716
rect 30739 14660 30795 14716
rect 30795 14660 30799 14716
rect 30735 14656 30799 14660
rect 9392 14172 9456 14176
rect 9392 14116 9396 14172
rect 9396 14116 9452 14172
rect 9452 14116 9456 14172
rect 9392 14112 9456 14116
rect 9472 14172 9536 14176
rect 9472 14116 9476 14172
rect 9476 14116 9532 14172
rect 9532 14116 9536 14172
rect 9472 14112 9536 14116
rect 9552 14172 9616 14176
rect 9552 14116 9556 14172
rect 9556 14116 9612 14172
rect 9612 14116 9616 14172
rect 9552 14112 9616 14116
rect 9632 14172 9696 14176
rect 9632 14116 9636 14172
rect 9636 14116 9692 14172
rect 9692 14116 9696 14172
rect 9632 14112 9696 14116
rect 17833 14172 17897 14176
rect 17833 14116 17837 14172
rect 17837 14116 17893 14172
rect 17893 14116 17897 14172
rect 17833 14112 17897 14116
rect 17913 14172 17977 14176
rect 17913 14116 17917 14172
rect 17917 14116 17973 14172
rect 17973 14116 17977 14172
rect 17913 14112 17977 14116
rect 17993 14172 18057 14176
rect 17993 14116 17997 14172
rect 17997 14116 18053 14172
rect 18053 14116 18057 14172
rect 17993 14112 18057 14116
rect 18073 14172 18137 14176
rect 18073 14116 18077 14172
rect 18077 14116 18133 14172
rect 18133 14116 18137 14172
rect 18073 14112 18137 14116
rect 26274 14172 26338 14176
rect 26274 14116 26278 14172
rect 26278 14116 26334 14172
rect 26334 14116 26338 14172
rect 26274 14112 26338 14116
rect 26354 14172 26418 14176
rect 26354 14116 26358 14172
rect 26358 14116 26414 14172
rect 26414 14116 26418 14172
rect 26354 14112 26418 14116
rect 26434 14172 26498 14176
rect 26434 14116 26438 14172
rect 26438 14116 26494 14172
rect 26494 14116 26498 14172
rect 26434 14112 26498 14116
rect 26514 14172 26578 14176
rect 26514 14116 26518 14172
rect 26518 14116 26574 14172
rect 26574 14116 26578 14172
rect 26514 14112 26578 14116
rect 34715 14172 34779 14176
rect 34715 14116 34719 14172
rect 34719 14116 34775 14172
rect 34775 14116 34779 14172
rect 34715 14112 34779 14116
rect 34795 14172 34859 14176
rect 34795 14116 34799 14172
rect 34799 14116 34855 14172
rect 34855 14116 34859 14172
rect 34795 14112 34859 14116
rect 34875 14172 34939 14176
rect 34875 14116 34879 14172
rect 34879 14116 34935 14172
rect 34935 14116 34939 14172
rect 34875 14112 34939 14116
rect 34955 14172 35019 14176
rect 34955 14116 34959 14172
rect 34959 14116 35015 14172
rect 35015 14116 35019 14172
rect 34955 14112 35019 14116
rect 5172 13628 5236 13632
rect 5172 13572 5176 13628
rect 5176 13572 5232 13628
rect 5232 13572 5236 13628
rect 5172 13568 5236 13572
rect 5252 13628 5316 13632
rect 5252 13572 5256 13628
rect 5256 13572 5312 13628
rect 5312 13572 5316 13628
rect 5252 13568 5316 13572
rect 5332 13628 5396 13632
rect 5332 13572 5336 13628
rect 5336 13572 5392 13628
rect 5392 13572 5396 13628
rect 5332 13568 5396 13572
rect 5412 13628 5476 13632
rect 5412 13572 5416 13628
rect 5416 13572 5472 13628
rect 5472 13572 5476 13628
rect 5412 13568 5476 13572
rect 13613 13628 13677 13632
rect 13613 13572 13617 13628
rect 13617 13572 13673 13628
rect 13673 13572 13677 13628
rect 13613 13568 13677 13572
rect 13693 13628 13757 13632
rect 13693 13572 13697 13628
rect 13697 13572 13753 13628
rect 13753 13572 13757 13628
rect 13693 13568 13757 13572
rect 13773 13628 13837 13632
rect 13773 13572 13777 13628
rect 13777 13572 13833 13628
rect 13833 13572 13837 13628
rect 13773 13568 13837 13572
rect 13853 13628 13917 13632
rect 13853 13572 13857 13628
rect 13857 13572 13913 13628
rect 13913 13572 13917 13628
rect 13853 13568 13917 13572
rect 22054 13628 22118 13632
rect 22054 13572 22058 13628
rect 22058 13572 22114 13628
rect 22114 13572 22118 13628
rect 22054 13568 22118 13572
rect 22134 13628 22198 13632
rect 22134 13572 22138 13628
rect 22138 13572 22194 13628
rect 22194 13572 22198 13628
rect 22134 13568 22198 13572
rect 22214 13628 22278 13632
rect 22214 13572 22218 13628
rect 22218 13572 22274 13628
rect 22274 13572 22278 13628
rect 22214 13568 22278 13572
rect 22294 13628 22358 13632
rect 22294 13572 22298 13628
rect 22298 13572 22354 13628
rect 22354 13572 22358 13628
rect 22294 13568 22358 13572
rect 30495 13628 30559 13632
rect 30495 13572 30499 13628
rect 30499 13572 30555 13628
rect 30555 13572 30559 13628
rect 30495 13568 30559 13572
rect 30575 13628 30639 13632
rect 30575 13572 30579 13628
rect 30579 13572 30635 13628
rect 30635 13572 30639 13628
rect 30575 13568 30639 13572
rect 30655 13628 30719 13632
rect 30655 13572 30659 13628
rect 30659 13572 30715 13628
rect 30715 13572 30719 13628
rect 30655 13568 30719 13572
rect 30735 13628 30799 13632
rect 30735 13572 30739 13628
rect 30739 13572 30795 13628
rect 30795 13572 30799 13628
rect 30735 13568 30799 13572
rect 9392 13084 9456 13088
rect 9392 13028 9396 13084
rect 9396 13028 9452 13084
rect 9452 13028 9456 13084
rect 9392 13024 9456 13028
rect 9472 13084 9536 13088
rect 9472 13028 9476 13084
rect 9476 13028 9532 13084
rect 9532 13028 9536 13084
rect 9472 13024 9536 13028
rect 9552 13084 9616 13088
rect 9552 13028 9556 13084
rect 9556 13028 9612 13084
rect 9612 13028 9616 13084
rect 9552 13024 9616 13028
rect 9632 13084 9696 13088
rect 9632 13028 9636 13084
rect 9636 13028 9692 13084
rect 9692 13028 9696 13084
rect 9632 13024 9696 13028
rect 17833 13084 17897 13088
rect 17833 13028 17837 13084
rect 17837 13028 17893 13084
rect 17893 13028 17897 13084
rect 17833 13024 17897 13028
rect 17913 13084 17977 13088
rect 17913 13028 17917 13084
rect 17917 13028 17973 13084
rect 17973 13028 17977 13084
rect 17913 13024 17977 13028
rect 17993 13084 18057 13088
rect 17993 13028 17997 13084
rect 17997 13028 18053 13084
rect 18053 13028 18057 13084
rect 17993 13024 18057 13028
rect 18073 13084 18137 13088
rect 18073 13028 18077 13084
rect 18077 13028 18133 13084
rect 18133 13028 18137 13084
rect 18073 13024 18137 13028
rect 26274 13084 26338 13088
rect 26274 13028 26278 13084
rect 26278 13028 26334 13084
rect 26334 13028 26338 13084
rect 26274 13024 26338 13028
rect 26354 13084 26418 13088
rect 26354 13028 26358 13084
rect 26358 13028 26414 13084
rect 26414 13028 26418 13084
rect 26354 13024 26418 13028
rect 26434 13084 26498 13088
rect 26434 13028 26438 13084
rect 26438 13028 26494 13084
rect 26494 13028 26498 13084
rect 26434 13024 26498 13028
rect 26514 13084 26578 13088
rect 26514 13028 26518 13084
rect 26518 13028 26574 13084
rect 26574 13028 26578 13084
rect 26514 13024 26578 13028
rect 34715 13084 34779 13088
rect 34715 13028 34719 13084
rect 34719 13028 34775 13084
rect 34775 13028 34779 13084
rect 34715 13024 34779 13028
rect 34795 13084 34859 13088
rect 34795 13028 34799 13084
rect 34799 13028 34855 13084
rect 34855 13028 34859 13084
rect 34795 13024 34859 13028
rect 34875 13084 34939 13088
rect 34875 13028 34879 13084
rect 34879 13028 34935 13084
rect 34935 13028 34939 13084
rect 34875 13024 34939 13028
rect 34955 13084 35019 13088
rect 34955 13028 34959 13084
rect 34959 13028 35015 13084
rect 35015 13028 35019 13084
rect 34955 13024 35019 13028
rect 5172 12540 5236 12544
rect 5172 12484 5176 12540
rect 5176 12484 5232 12540
rect 5232 12484 5236 12540
rect 5172 12480 5236 12484
rect 5252 12540 5316 12544
rect 5252 12484 5256 12540
rect 5256 12484 5312 12540
rect 5312 12484 5316 12540
rect 5252 12480 5316 12484
rect 5332 12540 5396 12544
rect 5332 12484 5336 12540
rect 5336 12484 5392 12540
rect 5392 12484 5396 12540
rect 5332 12480 5396 12484
rect 5412 12540 5476 12544
rect 5412 12484 5416 12540
rect 5416 12484 5472 12540
rect 5472 12484 5476 12540
rect 5412 12480 5476 12484
rect 13613 12540 13677 12544
rect 13613 12484 13617 12540
rect 13617 12484 13673 12540
rect 13673 12484 13677 12540
rect 13613 12480 13677 12484
rect 13693 12540 13757 12544
rect 13693 12484 13697 12540
rect 13697 12484 13753 12540
rect 13753 12484 13757 12540
rect 13693 12480 13757 12484
rect 13773 12540 13837 12544
rect 13773 12484 13777 12540
rect 13777 12484 13833 12540
rect 13833 12484 13837 12540
rect 13773 12480 13837 12484
rect 13853 12540 13917 12544
rect 13853 12484 13857 12540
rect 13857 12484 13913 12540
rect 13913 12484 13917 12540
rect 13853 12480 13917 12484
rect 22054 12540 22118 12544
rect 22054 12484 22058 12540
rect 22058 12484 22114 12540
rect 22114 12484 22118 12540
rect 22054 12480 22118 12484
rect 22134 12540 22198 12544
rect 22134 12484 22138 12540
rect 22138 12484 22194 12540
rect 22194 12484 22198 12540
rect 22134 12480 22198 12484
rect 22214 12540 22278 12544
rect 22214 12484 22218 12540
rect 22218 12484 22274 12540
rect 22274 12484 22278 12540
rect 22214 12480 22278 12484
rect 22294 12540 22358 12544
rect 22294 12484 22298 12540
rect 22298 12484 22354 12540
rect 22354 12484 22358 12540
rect 22294 12480 22358 12484
rect 30495 12540 30559 12544
rect 30495 12484 30499 12540
rect 30499 12484 30555 12540
rect 30555 12484 30559 12540
rect 30495 12480 30559 12484
rect 30575 12540 30639 12544
rect 30575 12484 30579 12540
rect 30579 12484 30635 12540
rect 30635 12484 30639 12540
rect 30575 12480 30639 12484
rect 30655 12540 30719 12544
rect 30655 12484 30659 12540
rect 30659 12484 30715 12540
rect 30715 12484 30719 12540
rect 30655 12480 30719 12484
rect 30735 12540 30799 12544
rect 30735 12484 30739 12540
rect 30739 12484 30795 12540
rect 30795 12484 30799 12540
rect 30735 12480 30799 12484
rect 9392 11996 9456 12000
rect 9392 11940 9396 11996
rect 9396 11940 9452 11996
rect 9452 11940 9456 11996
rect 9392 11936 9456 11940
rect 9472 11996 9536 12000
rect 9472 11940 9476 11996
rect 9476 11940 9532 11996
rect 9532 11940 9536 11996
rect 9472 11936 9536 11940
rect 9552 11996 9616 12000
rect 9552 11940 9556 11996
rect 9556 11940 9612 11996
rect 9612 11940 9616 11996
rect 9552 11936 9616 11940
rect 9632 11996 9696 12000
rect 9632 11940 9636 11996
rect 9636 11940 9692 11996
rect 9692 11940 9696 11996
rect 9632 11936 9696 11940
rect 17833 11996 17897 12000
rect 17833 11940 17837 11996
rect 17837 11940 17893 11996
rect 17893 11940 17897 11996
rect 17833 11936 17897 11940
rect 17913 11996 17977 12000
rect 17913 11940 17917 11996
rect 17917 11940 17973 11996
rect 17973 11940 17977 11996
rect 17913 11936 17977 11940
rect 17993 11996 18057 12000
rect 17993 11940 17997 11996
rect 17997 11940 18053 11996
rect 18053 11940 18057 11996
rect 17993 11936 18057 11940
rect 18073 11996 18137 12000
rect 18073 11940 18077 11996
rect 18077 11940 18133 11996
rect 18133 11940 18137 11996
rect 18073 11936 18137 11940
rect 26274 11996 26338 12000
rect 26274 11940 26278 11996
rect 26278 11940 26334 11996
rect 26334 11940 26338 11996
rect 26274 11936 26338 11940
rect 26354 11996 26418 12000
rect 26354 11940 26358 11996
rect 26358 11940 26414 11996
rect 26414 11940 26418 11996
rect 26354 11936 26418 11940
rect 26434 11996 26498 12000
rect 26434 11940 26438 11996
rect 26438 11940 26494 11996
rect 26494 11940 26498 11996
rect 26434 11936 26498 11940
rect 26514 11996 26578 12000
rect 26514 11940 26518 11996
rect 26518 11940 26574 11996
rect 26574 11940 26578 11996
rect 26514 11936 26578 11940
rect 34715 11996 34779 12000
rect 34715 11940 34719 11996
rect 34719 11940 34775 11996
rect 34775 11940 34779 11996
rect 34715 11936 34779 11940
rect 34795 11996 34859 12000
rect 34795 11940 34799 11996
rect 34799 11940 34855 11996
rect 34855 11940 34859 11996
rect 34795 11936 34859 11940
rect 34875 11996 34939 12000
rect 34875 11940 34879 11996
rect 34879 11940 34935 11996
rect 34935 11940 34939 11996
rect 34875 11936 34939 11940
rect 34955 11996 35019 12000
rect 34955 11940 34959 11996
rect 34959 11940 35015 11996
rect 35015 11940 35019 11996
rect 34955 11936 35019 11940
rect 5172 11452 5236 11456
rect 5172 11396 5176 11452
rect 5176 11396 5232 11452
rect 5232 11396 5236 11452
rect 5172 11392 5236 11396
rect 5252 11452 5316 11456
rect 5252 11396 5256 11452
rect 5256 11396 5312 11452
rect 5312 11396 5316 11452
rect 5252 11392 5316 11396
rect 5332 11452 5396 11456
rect 5332 11396 5336 11452
rect 5336 11396 5392 11452
rect 5392 11396 5396 11452
rect 5332 11392 5396 11396
rect 5412 11452 5476 11456
rect 5412 11396 5416 11452
rect 5416 11396 5472 11452
rect 5472 11396 5476 11452
rect 5412 11392 5476 11396
rect 13613 11452 13677 11456
rect 13613 11396 13617 11452
rect 13617 11396 13673 11452
rect 13673 11396 13677 11452
rect 13613 11392 13677 11396
rect 13693 11452 13757 11456
rect 13693 11396 13697 11452
rect 13697 11396 13753 11452
rect 13753 11396 13757 11452
rect 13693 11392 13757 11396
rect 13773 11452 13837 11456
rect 13773 11396 13777 11452
rect 13777 11396 13833 11452
rect 13833 11396 13837 11452
rect 13773 11392 13837 11396
rect 13853 11452 13917 11456
rect 13853 11396 13857 11452
rect 13857 11396 13913 11452
rect 13913 11396 13917 11452
rect 13853 11392 13917 11396
rect 22054 11452 22118 11456
rect 22054 11396 22058 11452
rect 22058 11396 22114 11452
rect 22114 11396 22118 11452
rect 22054 11392 22118 11396
rect 22134 11452 22198 11456
rect 22134 11396 22138 11452
rect 22138 11396 22194 11452
rect 22194 11396 22198 11452
rect 22134 11392 22198 11396
rect 22214 11452 22278 11456
rect 22214 11396 22218 11452
rect 22218 11396 22274 11452
rect 22274 11396 22278 11452
rect 22214 11392 22278 11396
rect 22294 11452 22358 11456
rect 22294 11396 22298 11452
rect 22298 11396 22354 11452
rect 22354 11396 22358 11452
rect 22294 11392 22358 11396
rect 30495 11452 30559 11456
rect 30495 11396 30499 11452
rect 30499 11396 30555 11452
rect 30555 11396 30559 11452
rect 30495 11392 30559 11396
rect 30575 11452 30639 11456
rect 30575 11396 30579 11452
rect 30579 11396 30635 11452
rect 30635 11396 30639 11452
rect 30575 11392 30639 11396
rect 30655 11452 30719 11456
rect 30655 11396 30659 11452
rect 30659 11396 30715 11452
rect 30715 11396 30719 11452
rect 30655 11392 30719 11396
rect 30735 11452 30799 11456
rect 30735 11396 30739 11452
rect 30739 11396 30795 11452
rect 30795 11396 30799 11452
rect 30735 11392 30799 11396
rect 9392 10908 9456 10912
rect 9392 10852 9396 10908
rect 9396 10852 9452 10908
rect 9452 10852 9456 10908
rect 9392 10848 9456 10852
rect 9472 10908 9536 10912
rect 9472 10852 9476 10908
rect 9476 10852 9532 10908
rect 9532 10852 9536 10908
rect 9472 10848 9536 10852
rect 9552 10908 9616 10912
rect 9552 10852 9556 10908
rect 9556 10852 9612 10908
rect 9612 10852 9616 10908
rect 9552 10848 9616 10852
rect 9632 10908 9696 10912
rect 9632 10852 9636 10908
rect 9636 10852 9692 10908
rect 9692 10852 9696 10908
rect 9632 10848 9696 10852
rect 17833 10908 17897 10912
rect 17833 10852 17837 10908
rect 17837 10852 17893 10908
rect 17893 10852 17897 10908
rect 17833 10848 17897 10852
rect 17913 10908 17977 10912
rect 17913 10852 17917 10908
rect 17917 10852 17973 10908
rect 17973 10852 17977 10908
rect 17913 10848 17977 10852
rect 17993 10908 18057 10912
rect 17993 10852 17997 10908
rect 17997 10852 18053 10908
rect 18053 10852 18057 10908
rect 17993 10848 18057 10852
rect 18073 10908 18137 10912
rect 18073 10852 18077 10908
rect 18077 10852 18133 10908
rect 18133 10852 18137 10908
rect 18073 10848 18137 10852
rect 26274 10908 26338 10912
rect 26274 10852 26278 10908
rect 26278 10852 26334 10908
rect 26334 10852 26338 10908
rect 26274 10848 26338 10852
rect 26354 10908 26418 10912
rect 26354 10852 26358 10908
rect 26358 10852 26414 10908
rect 26414 10852 26418 10908
rect 26354 10848 26418 10852
rect 26434 10908 26498 10912
rect 26434 10852 26438 10908
rect 26438 10852 26494 10908
rect 26494 10852 26498 10908
rect 26434 10848 26498 10852
rect 26514 10908 26578 10912
rect 26514 10852 26518 10908
rect 26518 10852 26574 10908
rect 26574 10852 26578 10908
rect 26514 10848 26578 10852
rect 34715 10908 34779 10912
rect 34715 10852 34719 10908
rect 34719 10852 34775 10908
rect 34775 10852 34779 10908
rect 34715 10848 34779 10852
rect 34795 10908 34859 10912
rect 34795 10852 34799 10908
rect 34799 10852 34855 10908
rect 34855 10852 34859 10908
rect 34795 10848 34859 10852
rect 34875 10908 34939 10912
rect 34875 10852 34879 10908
rect 34879 10852 34935 10908
rect 34935 10852 34939 10908
rect 34875 10848 34939 10852
rect 34955 10908 35019 10912
rect 34955 10852 34959 10908
rect 34959 10852 35015 10908
rect 35015 10852 35019 10908
rect 34955 10848 35019 10852
rect 5172 10364 5236 10368
rect 5172 10308 5176 10364
rect 5176 10308 5232 10364
rect 5232 10308 5236 10364
rect 5172 10304 5236 10308
rect 5252 10364 5316 10368
rect 5252 10308 5256 10364
rect 5256 10308 5312 10364
rect 5312 10308 5316 10364
rect 5252 10304 5316 10308
rect 5332 10364 5396 10368
rect 5332 10308 5336 10364
rect 5336 10308 5392 10364
rect 5392 10308 5396 10364
rect 5332 10304 5396 10308
rect 5412 10364 5476 10368
rect 5412 10308 5416 10364
rect 5416 10308 5472 10364
rect 5472 10308 5476 10364
rect 5412 10304 5476 10308
rect 13613 10364 13677 10368
rect 13613 10308 13617 10364
rect 13617 10308 13673 10364
rect 13673 10308 13677 10364
rect 13613 10304 13677 10308
rect 13693 10364 13757 10368
rect 13693 10308 13697 10364
rect 13697 10308 13753 10364
rect 13753 10308 13757 10364
rect 13693 10304 13757 10308
rect 13773 10364 13837 10368
rect 13773 10308 13777 10364
rect 13777 10308 13833 10364
rect 13833 10308 13837 10364
rect 13773 10304 13837 10308
rect 13853 10364 13917 10368
rect 13853 10308 13857 10364
rect 13857 10308 13913 10364
rect 13913 10308 13917 10364
rect 13853 10304 13917 10308
rect 22054 10364 22118 10368
rect 22054 10308 22058 10364
rect 22058 10308 22114 10364
rect 22114 10308 22118 10364
rect 22054 10304 22118 10308
rect 22134 10364 22198 10368
rect 22134 10308 22138 10364
rect 22138 10308 22194 10364
rect 22194 10308 22198 10364
rect 22134 10304 22198 10308
rect 22214 10364 22278 10368
rect 22214 10308 22218 10364
rect 22218 10308 22274 10364
rect 22274 10308 22278 10364
rect 22214 10304 22278 10308
rect 22294 10364 22358 10368
rect 22294 10308 22298 10364
rect 22298 10308 22354 10364
rect 22354 10308 22358 10364
rect 22294 10304 22358 10308
rect 30495 10364 30559 10368
rect 30495 10308 30499 10364
rect 30499 10308 30555 10364
rect 30555 10308 30559 10364
rect 30495 10304 30559 10308
rect 30575 10364 30639 10368
rect 30575 10308 30579 10364
rect 30579 10308 30635 10364
rect 30635 10308 30639 10364
rect 30575 10304 30639 10308
rect 30655 10364 30719 10368
rect 30655 10308 30659 10364
rect 30659 10308 30715 10364
rect 30715 10308 30719 10364
rect 30655 10304 30719 10308
rect 30735 10364 30799 10368
rect 30735 10308 30739 10364
rect 30739 10308 30795 10364
rect 30795 10308 30799 10364
rect 30735 10304 30799 10308
rect 9392 9820 9456 9824
rect 9392 9764 9396 9820
rect 9396 9764 9452 9820
rect 9452 9764 9456 9820
rect 9392 9760 9456 9764
rect 9472 9820 9536 9824
rect 9472 9764 9476 9820
rect 9476 9764 9532 9820
rect 9532 9764 9536 9820
rect 9472 9760 9536 9764
rect 9552 9820 9616 9824
rect 9552 9764 9556 9820
rect 9556 9764 9612 9820
rect 9612 9764 9616 9820
rect 9552 9760 9616 9764
rect 9632 9820 9696 9824
rect 9632 9764 9636 9820
rect 9636 9764 9692 9820
rect 9692 9764 9696 9820
rect 9632 9760 9696 9764
rect 17833 9820 17897 9824
rect 17833 9764 17837 9820
rect 17837 9764 17893 9820
rect 17893 9764 17897 9820
rect 17833 9760 17897 9764
rect 17913 9820 17977 9824
rect 17913 9764 17917 9820
rect 17917 9764 17973 9820
rect 17973 9764 17977 9820
rect 17913 9760 17977 9764
rect 17993 9820 18057 9824
rect 17993 9764 17997 9820
rect 17997 9764 18053 9820
rect 18053 9764 18057 9820
rect 17993 9760 18057 9764
rect 18073 9820 18137 9824
rect 18073 9764 18077 9820
rect 18077 9764 18133 9820
rect 18133 9764 18137 9820
rect 18073 9760 18137 9764
rect 26274 9820 26338 9824
rect 26274 9764 26278 9820
rect 26278 9764 26334 9820
rect 26334 9764 26338 9820
rect 26274 9760 26338 9764
rect 26354 9820 26418 9824
rect 26354 9764 26358 9820
rect 26358 9764 26414 9820
rect 26414 9764 26418 9820
rect 26354 9760 26418 9764
rect 26434 9820 26498 9824
rect 26434 9764 26438 9820
rect 26438 9764 26494 9820
rect 26494 9764 26498 9820
rect 26434 9760 26498 9764
rect 26514 9820 26578 9824
rect 26514 9764 26518 9820
rect 26518 9764 26574 9820
rect 26574 9764 26578 9820
rect 26514 9760 26578 9764
rect 34715 9820 34779 9824
rect 34715 9764 34719 9820
rect 34719 9764 34775 9820
rect 34775 9764 34779 9820
rect 34715 9760 34779 9764
rect 34795 9820 34859 9824
rect 34795 9764 34799 9820
rect 34799 9764 34855 9820
rect 34855 9764 34859 9820
rect 34795 9760 34859 9764
rect 34875 9820 34939 9824
rect 34875 9764 34879 9820
rect 34879 9764 34935 9820
rect 34935 9764 34939 9820
rect 34875 9760 34939 9764
rect 34955 9820 35019 9824
rect 34955 9764 34959 9820
rect 34959 9764 35015 9820
rect 35015 9764 35019 9820
rect 34955 9760 35019 9764
rect 5172 9276 5236 9280
rect 5172 9220 5176 9276
rect 5176 9220 5232 9276
rect 5232 9220 5236 9276
rect 5172 9216 5236 9220
rect 5252 9276 5316 9280
rect 5252 9220 5256 9276
rect 5256 9220 5312 9276
rect 5312 9220 5316 9276
rect 5252 9216 5316 9220
rect 5332 9276 5396 9280
rect 5332 9220 5336 9276
rect 5336 9220 5392 9276
rect 5392 9220 5396 9276
rect 5332 9216 5396 9220
rect 5412 9276 5476 9280
rect 5412 9220 5416 9276
rect 5416 9220 5472 9276
rect 5472 9220 5476 9276
rect 5412 9216 5476 9220
rect 13613 9276 13677 9280
rect 13613 9220 13617 9276
rect 13617 9220 13673 9276
rect 13673 9220 13677 9276
rect 13613 9216 13677 9220
rect 13693 9276 13757 9280
rect 13693 9220 13697 9276
rect 13697 9220 13753 9276
rect 13753 9220 13757 9276
rect 13693 9216 13757 9220
rect 13773 9276 13837 9280
rect 13773 9220 13777 9276
rect 13777 9220 13833 9276
rect 13833 9220 13837 9276
rect 13773 9216 13837 9220
rect 13853 9276 13917 9280
rect 13853 9220 13857 9276
rect 13857 9220 13913 9276
rect 13913 9220 13917 9276
rect 13853 9216 13917 9220
rect 22054 9276 22118 9280
rect 22054 9220 22058 9276
rect 22058 9220 22114 9276
rect 22114 9220 22118 9276
rect 22054 9216 22118 9220
rect 22134 9276 22198 9280
rect 22134 9220 22138 9276
rect 22138 9220 22194 9276
rect 22194 9220 22198 9276
rect 22134 9216 22198 9220
rect 22214 9276 22278 9280
rect 22214 9220 22218 9276
rect 22218 9220 22274 9276
rect 22274 9220 22278 9276
rect 22214 9216 22278 9220
rect 22294 9276 22358 9280
rect 22294 9220 22298 9276
rect 22298 9220 22354 9276
rect 22354 9220 22358 9276
rect 22294 9216 22358 9220
rect 30495 9276 30559 9280
rect 30495 9220 30499 9276
rect 30499 9220 30555 9276
rect 30555 9220 30559 9276
rect 30495 9216 30559 9220
rect 30575 9276 30639 9280
rect 30575 9220 30579 9276
rect 30579 9220 30635 9276
rect 30635 9220 30639 9276
rect 30575 9216 30639 9220
rect 30655 9276 30719 9280
rect 30655 9220 30659 9276
rect 30659 9220 30715 9276
rect 30715 9220 30719 9276
rect 30655 9216 30719 9220
rect 30735 9276 30799 9280
rect 30735 9220 30739 9276
rect 30739 9220 30795 9276
rect 30795 9220 30799 9276
rect 30735 9216 30799 9220
rect 9392 8732 9456 8736
rect 9392 8676 9396 8732
rect 9396 8676 9452 8732
rect 9452 8676 9456 8732
rect 9392 8672 9456 8676
rect 9472 8732 9536 8736
rect 9472 8676 9476 8732
rect 9476 8676 9532 8732
rect 9532 8676 9536 8732
rect 9472 8672 9536 8676
rect 9552 8732 9616 8736
rect 9552 8676 9556 8732
rect 9556 8676 9612 8732
rect 9612 8676 9616 8732
rect 9552 8672 9616 8676
rect 9632 8732 9696 8736
rect 9632 8676 9636 8732
rect 9636 8676 9692 8732
rect 9692 8676 9696 8732
rect 9632 8672 9696 8676
rect 17833 8732 17897 8736
rect 17833 8676 17837 8732
rect 17837 8676 17893 8732
rect 17893 8676 17897 8732
rect 17833 8672 17897 8676
rect 17913 8732 17977 8736
rect 17913 8676 17917 8732
rect 17917 8676 17973 8732
rect 17973 8676 17977 8732
rect 17913 8672 17977 8676
rect 17993 8732 18057 8736
rect 17993 8676 17997 8732
rect 17997 8676 18053 8732
rect 18053 8676 18057 8732
rect 17993 8672 18057 8676
rect 18073 8732 18137 8736
rect 18073 8676 18077 8732
rect 18077 8676 18133 8732
rect 18133 8676 18137 8732
rect 18073 8672 18137 8676
rect 26274 8732 26338 8736
rect 26274 8676 26278 8732
rect 26278 8676 26334 8732
rect 26334 8676 26338 8732
rect 26274 8672 26338 8676
rect 26354 8732 26418 8736
rect 26354 8676 26358 8732
rect 26358 8676 26414 8732
rect 26414 8676 26418 8732
rect 26354 8672 26418 8676
rect 26434 8732 26498 8736
rect 26434 8676 26438 8732
rect 26438 8676 26494 8732
rect 26494 8676 26498 8732
rect 26434 8672 26498 8676
rect 26514 8732 26578 8736
rect 26514 8676 26518 8732
rect 26518 8676 26574 8732
rect 26574 8676 26578 8732
rect 26514 8672 26578 8676
rect 34715 8732 34779 8736
rect 34715 8676 34719 8732
rect 34719 8676 34775 8732
rect 34775 8676 34779 8732
rect 34715 8672 34779 8676
rect 34795 8732 34859 8736
rect 34795 8676 34799 8732
rect 34799 8676 34855 8732
rect 34855 8676 34859 8732
rect 34795 8672 34859 8676
rect 34875 8732 34939 8736
rect 34875 8676 34879 8732
rect 34879 8676 34935 8732
rect 34935 8676 34939 8732
rect 34875 8672 34939 8676
rect 34955 8732 35019 8736
rect 34955 8676 34959 8732
rect 34959 8676 35015 8732
rect 35015 8676 35019 8732
rect 34955 8672 35019 8676
rect 5172 8188 5236 8192
rect 5172 8132 5176 8188
rect 5176 8132 5232 8188
rect 5232 8132 5236 8188
rect 5172 8128 5236 8132
rect 5252 8188 5316 8192
rect 5252 8132 5256 8188
rect 5256 8132 5312 8188
rect 5312 8132 5316 8188
rect 5252 8128 5316 8132
rect 5332 8188 5396 8192
rect 5332 8132 5336 8188
rect 5336 8132 5392 8188
rect 5392 8132 5396 8188
rect 5332 8128 5396 8132
rect 5412 8188 5476 8192
rect 5412 8132 5416 8188
rect 5416 8132 5472 8188
rect 5472 8132 5476 8188
rect 5412 8128 5476 8132
rect 13613 8188 13677 8192
rect 13613 8132 13617 8188
rect 13617 8132 13673 8188
rect 13673 8132 13677 8188
rect 13613 8128 13677 8132
rect 13693 8188 13757 8192
rect 13693 8132 13697 8188
rect 13697 8132 13753 8188
rect 13753 8132 13757 8188
rect 13693 8128 13757 8132
rect 13773 8188 13837 8192
rect 13773 8132 13777 8188
rect 13777 8132 13833 8188
rect 13833 8132 13837 8188
rect 13773 8128 13837 8132
rect 13853 8188 13917 8192
rect 13853 8132 13857 8188
rect 13857 8132 13913 8188
rect 13913 8132 13917 8188
rect 13853 8128 13917 8132
rect 22054 8188 22118 8192
rect 22054 8132 22058 8188
rect 22058 8132 22114 8188
rect 22114 8132 22118 8188
rect 22054 8128 22118 8132
rect 22134 8188 22198 8192
rect 22134 8132 22138 8188
rect 22138 8132 22194 8188
rect 22194 8132 22198 8188
rect 22134 8128 22198 8132
rect 22214 8188 22278 8192
rect 22214 8132 22218 8188
rect 22218 8132 22274 8188
rect 22274 8132 22278 8188
rect 22214 8128 22278 8132
rect 22294 8188 22358 8192
rect 22294 8132 22298 8188
rect 22298 8132 22354 8188
rect 22354 8132 22358 8188
rect 22294 8128 22358 8132
rect 30495 8188 30559 8192
rect 30495 8132 30499 8188
rect 30499 8132 30555 8188
rect 30555 8132 30559 8188
rect 30495 8128 30559 8132
rect 30575 8188 30639 8192
rect 30575 8132 30579 8188
rect 30579 8132 30635 8188
rect 30635 8132 30639 8188
rect 30575 8128 30639 8132
rect 30655 8188 30719 8192
rect 30655 8132 30659 8188
rect 30659 8132 30715 8188
rect 30715 8132 30719 8188
rect 30655 8128 30719 8132
rect 30735 8188 30799 8192
rect 30735 8132 30739 8188
rect 30739 8132 30795 8188
rect 30795 8132 30799 8188
rect 30735 8128 30799 8132
rect 9392 7644 9456 7648
rect 9392 7588 9396 7644
rect 9396 7588 9452 7644
rect 9452 7588 9456 7644
rect 9392 7584 9456 7588
rect 9472 7644 9536 7648
rect 9472 7588 9476 7644
rect 9476 7588 9532 7644
rect 9532 7588 9536 7644
rect 9472 7584 9536 7588
rect 9552 7644 9616 7648
rect 9552 7588 9556 7644
rect 9556 7588 9612 7644
rect 9612 7588 9616 7644
rect 9552 7584 9616 7588
rect 9632 7644 9696 7648
rect 9632 7588 9636 7644
rect 9636 7588 9692 7644
rect 9692 7588 9696 7644
rect 9632 7584 9696 7588
rect 17833 7644 17897 7648
rect 17833 7588 17837 7644
rect 17837 7588 17893 7644
rect 17893 7588 17897 7644
rect 17833 7584 17897 7588
rect 17913 7644 17977 7648
rect 17913 7588 17917 7644
rect 17917 7588 17973 7644
rect 17973 7588 17977 7644
rect 17913 7584 17977 7588
rect 17993 7644 18057 7648
rect 17993 7588 17997 7644
rect 17997 7588 18053 7644
rect 18053 7588 18057 7644
rect 17993 7584 18057 7588
rect 18073 7644 18137 7648
rect 18073 7588 18077 7644
rect 18077 7588 18133 7644
rect 18133 7588 18137 7644
rect 18073 7584 18137 7588
rect 26274 7644 26338 7648
rect 26274 7588 26278 7644
rect 26278 7588 26334 7644
rect 26334 7588 26338 7644
rect 26274 7584 26338 7588
rect 26354 7644 26418 7648
rect 26354 7588 26358 7644
rect 26358 7588 26414 7644
rect 26414 7588 26418 7644
rect 26354 7584 26418 7588
rect 26434 7644 26498 7648
rect 26434 7588 26438 7644
rect 26438 7588 26494 7644
rect 26494 7588 26498 7644
rect 26434 7584 26498 7588
rect 26514 7644 26578 7648
rect 26514 7588 26518 7644
rect 26518 7588 26574 7644
rect 26574 7588 26578 7644
rect 26514 7584 26578 7588
rect 34715 7644 34779 7648
rect 34715 7588 34719 7644
rect 34719 7588 34775 7644
rect 34775 7588 34779 7644
rect 34715 7584 34779 7588
rect 34795 7644 34859 7648
rect 34795 7588 34799 7644
rect 34799 7588 34855 7644
rect 34855 7588 34859 7644
rect 34795 7584 34859 7588
rect 34875 7644 34939 7648
rect 34875 7588 34879 7644
rect 34879 7588 34935 7644
rect 34935 7588 34939 7644
rect 34875 7584 34939 7588
rect 34955 7644 35019 7648
rect 34955 7588 34959 7644
rect 34959 7588 35015 7644
rect 35015 7588 35019 7644
rect 34955 7584 35019 7588
rect 5172 7100 5236 7104
rect 5172 7044 5176 7100
rect 5176 7044 5232 7100
rect 5232 7044 5236 7100
rect 5172 7040 5236 7044
rect 5252 7100 5316 7104
rect 5252 7044 5256 7100
rect 5256 7044 5312 7100
rect 5312 7044 5316 7100
rect 5252 7040 5316 7044
rect 5332 7100 5396 7104
rect 5332 7044 5336 7100
rect 5336 7044 5392 7100
rect 5392 7044 5396 7100
rect 5332 7040 5396 7044
rect 5412 7100 5476 7104
rect 5412 7044 5416 7100
rect 5416 7044 5472 7100
rect 5472 7044 5476 7100
rect 5412 7040 5476 7044
rect 13613 7100 13677 7104
rect 13613 7044 13617 7100
rect 13617 7044 13673 7100
rect 13673 7044 13677 7100
rect 13613 7040 13677 7044
rect 13693 7100 13757 7104
rect 13693 7044 13697 7100
rect 13697 7044 13753 7100
rect 13753 7044 13757 7100
rect 13693 7040 13757 7044
rect 13773 7100 13837 7104
rect 13773 7044 13777 7100
rect 13777 7044 13833 7100
rect 13833 7044 13837 7100
rect 13773 7040 13837 7044
rect 13853 7100 13917 7104
rect 13853 7044 13857 7100
rect 13857 7044 13913 7100
rect 13913 7044 13917 7100
rect 13853 7040 13917 7044
rect 22054 7100 22118 7104
rect 22054 7044 22058 7100
rect 22058 7044 22114 7100
rect 22114 7044 22118 7100
rect 22054 7040 22118 7044
rect 22134 7100 22198 7104
rect 22134 7044 22138 7100
rect 22138 7044 22194 7100
rect 22194 7044 22198 7100
rect 22134 7040 22198 7044
rect 22214 7100 22278 7104
rect 22214 7044 22218 7100
rect 22218 7044 22274 7100
rect 22274 7044 22278 7100
rect 22214 7040 22278 7044
rect 22294 7100 22358 7104
rect 22294 7044 22298 7100
rect 22298 7044 22354 7100
rect 22354 7044 22358 7100
rect 22294 7040 22358 7044
rect 30495 7100 30559 7104
rect 30495 7044 30499 7100
rect 30499 7044 30555 7100
rect 30555 7044 30559 7100
rect 30495 7040 30559 7044
rect 30575 7100 30639 7104
rect 30575 7044 30579 7100
rect 30579 7044 30635 7100
rect 30635 7044 30639 7100
rect 30575 7040 30639 7044
rect 30655 7100 30719 7104
rect 30655 7044 30659 7100
rect 30659 7044 30715 7100
rect 30715 7044 30719 7100
rect 30655 7040 30719 7044
rect 30735 7100 30799 7104
rect 30735 7044 30739 7100
rect 30739 7044 30795 7100
rect 30795 7044 30799 7100
rect 30735 7040 30799 7044
rect 9392 6556 9456 6560
rect 9392 6500 9396 6556
rect 9396 6500 9452 6556
rect 9452 6500 9456 6556
rect 9392 6496 9456 6500
rect 9472 6556 9536 6560
rect 9472 6500 9476 6556
rect 9476 6500 9532 6556
rect 9532 6500 9536 6556
rect 9472 6496 9536 6500
rect 9552 6556 9616 6560
rect 9552 6500 9556 6556
rect 9556 6500 9612 6556
rect 9612 6500 9616 6556
rect 9552 6496 9616 6500
rect 9632 6556 9696 6560
rect 9632 6500 9636 6556
rect 9636 6500 9692 6556
rect 9692 6500 9696 6556
rect 9632 6496 9696 6500
rect 17833 6556 17897 6560
rect 17833 6500 17837 6556
rect 17837 6500 17893 6556
rect 17893 6500 17897 6556
rect 17833 6496 17897 6500
rect 17913 6556 17977 6560
rect 17913 6500 17917 6556
rect 17917 6500 17973 6556
rect 17973 6500 17977 6556
rect 17913 6496 17977 6500
rect 17993 6556 18057 6560
rect 17993 6500 17997 6556
rect 17997 6500 18053 6556
rect 18053 6500 18057 6556
rect 17993 6496 18057 6500
rect 18073 6556 18137 6560
rect 18073 6500 18077 6556
rect 18077 6500 18133 6556
rect 18133 6500 18137 6556
rect 18073 6496 18137 6500
rect 26274 6556 26338 6560
rect 26274 6500 26278 6556
rect 26278 6500 26334 6556
rect 26334 6500 26338 6556
rect 26274 6496 26338 6500
rect 26354 6556 26418 6560
rect 26354 6500 26358 6556
rect 26358 6500 26414 6556
rect 26414 6500 26418 6556
rect 26354 6496 26418 6500
rect 26434 6556 26498 6560
rect 26434 6500 26438 6556
rect 26438 6500 26494 6556
rect 26494 6500 26498 6556
rect 26434 6496 26498 6500
rect 26514 6556 26578 6560
rect 26514 6500 26518 6556
rect 26518 6500 26574 6556
rect 26574 6500 26578 6556
rect 26514 6496 26578 6500
rect 34715 6556 34779 6560
rect 34715 6500 34719 6556
rect 34719 6500 34775 6556
rect 34775 6500 34779 6556
rect 34715 6496 34779 6500
rect 34795 6556 34859 6560
rect 34795 6500 34799 6556
rect 34799 6500 34855 6556
rect 34855 6500 34859 6556
rect 34795 6496 34859 6500
rect 34875 6556 34939 6560
rect 34875 6500 34879 6556
rect 34879 6500 34935 6556
rect 34935 6500 34939 6556
rect 34875 6496 34939 6500
rect 34955 6556 35019 6560
rect 34955 6500 34959 6556
rect 34959 6500 35015 6556
rect 35015 6500 35019 6556
rect 34955 6496 35019 6500
rect 5172 6012 5236 6016
rect 5172 5956 5176 6012
rect 5176 5956 5232 6012
rect 5232 5956 5236 6012
rect 5172 5952 5236 5956
rect 5252 6012 5316 6016
rect 5252 5956 5256 6012
rect 5256 5956 5312 6012
rect 5312 5956 5316 6012
rect 5252 5952 5316 5956
rect 5332 6012 5396 6016
rect 5332 5956 5336 6012
rect 5336 5956 5392 6012
rect 5392 5956 5396 6012
rect 5332 5952 5396 5956
rect 5412 6012 5476 6016
rect 5412 5956 5416 6012
rect 5416 5956 5472 6012
rect 5472 5956 5476 6012
rect 5412 5952 5476 5956
rect 13613 6012 13677 6016
rect 13613 5956 13617 6012
rect 13617 5956 13673 6012
rect 13673 5956 13677 6012
rect 13613 5952 13677 5956
rect 13693 6012 13757 6016
rect 13693 5956 13697 6012
rect 13697 5956 13753 6012
rect 13753 5956 13757 6012
rect 13693 5952 13757 5956
rect 13773 6012 13837 6016
rect 13773 5956 13777 6012
rect 13777 5956 13833 6012
rect 13833 5956 13837 6012
rect 13773 5952 13837 5956
rect 13853 6012 13917 6016
rect 13853 5956 13857 6012
rect 13857 5956 13913 6012
rect 13913 5956 13917 6012
rect 13853 5952 13917 5956
rect 22054 6012 22118 6016
rect 22054 5956 22058 6012
rect 22058 5956 22114 6012
rect 22114 5956 22118 6012
rect 22054 5952 22118 5956
rect 22134 6012 22198 6016
rect 22134 5956 22138 6012
rect 22138 5956 22194 6012
rect 22194 5956 22198 6012
rect 22134 5952 22198 5956
rect 22214 6012 22278 6016
rect 22214 5956 22218 6012
rect 22218 5956 22274 6012
rect 22274 5956 22278 6012
rect 22214 5952 22278 5956
rect 22294 6012 22358 6016
rect 22294 5956 22298 6012
rect 22298 5956 22354 6012
rect 22354 5956 22358 6012
rect 22294 5952 22358 5956
rect 30495 6012 30559 6016
rect 30495 5956 30499 6012
rect 30499 5956 30555 6012
rect 30555 5956 30559 6012
rect 30495 5952 30559 5956
rect 30575 6012 30639 6016
rect 30575 5956 30579 6012
rect 30579 5956 30635 6012
rect 30635 5956 30639 6012
rect 30575 5952 30639 5956
rect 30655 6012 30719 6016
rect 30655 5956 30659 6012
rect 30659 5956 30715 6012
rect 30715 5956 30719 6012
rect 30655 5952 30719 5956
rect 30735 6012 30799 6016
rect 30735 5956 30739 6012
rect 30739 5956 30795 6012
rect 30795 5956 30799 6012
rect 30735 5952 30799 5956
rect 9392 5468 9456 5472
rect 9392 5412 9396 5468
rect 9396 5412 9452 5468
rect 9452 5412 9456 5468
rect 9392 5408 9456 5412
rect 9472 5468 9536 5472
rect 9472 5412 9476 5468
rect 9476 5412 9532 5468
rect 9532 5412 9536 5468
rect 9472 5408 9536 5412
rect 9552 5468 9616 5472
rect 9552 5412 9556 5468
rect 9556 5412 9612 5468
rect 9612 5412 9616 5468
rect 9552 5408 9616 5412
rect 9632 5468 9696 5472
rect 9632 5412 9636 5468
rect 9636 5412 9692 5468
rect 9692 5412 9696 5468
rect 9632 5408 9696 5412
rect 17833 5468 17897 5472
rect 17833 5412 17837 5468
rect 17837 5412 17893 5468
rect 17893 5412 17897 5468
rect 17833 5408 17897 5412
rect 17913 5468 17977 5472
rect 17913 5412 17917 5468
rect 17917 5412 17973 5468
rect 17973 5412 17977 5468
rect 17913 5408 17977 5412
rect 17993 5468 18057 5472
rect 17993 5412 17997 5468
rect 17997 5412 18053 5468
rect 18053 5412 18057 5468
rect 17993 5408 18057 5412
rect 18073 5468 18137 5472
rect 18073 5412 18077 5468
rect 18077 5412 18133 5468
rect 18133 5412 18137 5468
rect 18073 5408 18137 5412
rect 26274 5468 26338 5472
rect 26274 5412 26278 5468
rect 26278 5412 26334 5468
rect 26334 5412 26338 5468
rect 26274 5408 26338 5412
rect 26354 5468 26418 5472
rect 26354 5412 26358 5468
rect 26358 5412 26414 5468
rect 26414 5412 26418 5468
rect 26354 5408 26418 5412
rect 26434 5468 26498 5472
rect 26434 5412 26438 5468
rect 26438 5412 26494 5468
rect 26494 5412 26498 5468
rect 26434 5408 26498 5412
rect 26514 5468 26578 5472
rect 26514 5412 26518 5468
rect 26518 5412 26574 5468
rect 26574 5412 26578 5468
rect 26514 5408 26578 5412
rect 34715 5468 34779 5472
rect 34715 5412 34719 5468
rect 34719 5412 34775 5468
rect 34775 5412 34779 5468
rect 34715 5408 34779 5412
rect 34795 5468 34859 5472
rect 34795 5412 34799 5468
rect 34799 5412 34855 5468
rect 34855 5412 34859 5468
rect 34795 5408 34859 5412
rect 34875 5468 34939 5472
rect 34875 5412 34879 5468
rect 34879 5412 34935 5468
rect 34935 5412 34939 5468
rect 34875 5408 34939 5412
rect 34955 5468 35019 5472
rect 34955 5412 34959 5468
rect 34959 5412 35015 5468
rect 35015 5412 35019 5468
rect 34955 5408 35019 5412
rect 5172 4924 5236 4928
rect 5172 4868 5176 4924
rect 5176 4868 5232 4924
rect 5232 4868 5236 4924
rect 5172 4864 5236 4868
rect 5252 4924 5316 4928
rect 5252 4868 5256 4924
rect 5256 4868 5312 4924
rect 5312 4868 5316 4924
rect 5252 4864 5316 4868
rect 5332 4924 5396 4928
rect 5332 4868 5336 4924
rect 5336 4868 5392 4924
rect 5392 4868 5396 4924
rect 5332 4864 5396 4868
rect 5412 4924 5476 4928
rect 5412 4868 5416 4924
rect 5416 4868 5472 4924
rect 5472 4868 5476 4924
rect 5412 4864 5476 4868
rect 13613 4924 13677 4928
rect 13613 4868 13617 4924
rect 13617 4868 13673 4924
rect 13673 4868 13677 4924
rect 13613 4864 13677 4868
rect 13693 4924 13757 4928
rect 13693 4868 13697 4924
rect 13697 4868 13753 4924
rect 13753 4868 13757 4924
rect 13693 4864 13757 4868
rect 13773 4924 13837 4928
rect 13773 4868 13777 4924
rect 13777 4868 13833 4924
rect 13833 4868 13837 4924
rect 13773 4864 13837 4868
rect 13853 4924 13917 4928
rect 13853 4868 13857 4924
rect 13857 4868 13913 4924
rect 13913 4868 13917 4924
rect 13853 4864 13917 4868
rect 22054 4924 22118 4928
rect 22054 4868 22058 4924
rect 22058 4868 22114 4924
rect 22114 4868 22118 4924
rect 22054 4864 22118 4868
rect 22134 4924 22198 4928
rect 22134 4868 22138 4924
rect 22138 4868 22194 4924
rect 22194 4868 22198 4924
rect 22134 4864 22198 4868
rect 22214 4924 22278 4928
rect 22214 4868 22218 4924
rect 22218 4868 22274 4924
rect 22274 4868 22278 4924
rect 22214 4864 22278 4868
rect 22294 4924 22358 4928
rect 22294 4868 22298 4924
rect 22298 4868 22354 4924
rect 22354 4868 22358 4924
rect 22294 4864 22358 4868
rect 30495 4924 30559 4928
rect 30495 4868 30499 4924
rect 30499 4868 30555 4924
rect 30555 4868 30559 4924
rect 30495 4864 30559 4868
rect 30575 4924 30639 4928
rect 30575 4868 30579 4924
rect 30579 4868 30635 4924
rect 30635 4868 30639 4924
rect 30575 4864 30639 4868
rect 30655 4924 30719 4928
rect 30655 4868 30659 4924
rect 30659 4868 30715 4924
rect 30715 4868 30719 4924
rect 30655 4864 30719 4868
rect 30735 4924 30799 4928
rect 30735 4868 30739 4924
rect 30739 4868 30795 4924
rect 30795 4868 30799 4924
rect 30735 4864 30799 4868
rect 9392 4380 9456 4384
rect 9392 4324 9396 4380
rect 9396 4324 9452 4380
rect 9452 4324 9456 4380
rect 9392 4320 9456 4324
rect 9472 4380 9536 4384
rect 9472 4324 9476 4380
rect 9476 4324 9532 4380
rect 9532 4324 9536 4380
rect 9472 4320 9536 4324
rect 9552 4380 9616 4384
rect 9552 4324 9556 4380
rect 9556 4324 9612 4380
rect 9612 4324 9616 4380
rect 9552 4320 9616 4324
rect 9632 4380 9696 4384
rect 9632 4324 9636 4380
rect 9636 4324 9692 4380
rect 9692 4324 9696 4380
rect 9632 4320 9696 4324
rect 17833 4380 17897 4384
rect 17833 4324 17837 4380
rect 17837 4324 17893 4380
rect 17893 4324 17897 4380
rect 17833 4320 17897 4324
rect 17913 4380 17977 4384
rect 17913 4324 17917 4380
rect 17917 4324 17973 4380
rect 17973 4324 17977 4380
rect 17913 4320 17977 4324
rect 17993 4380 18057 4384
rect 17993 4324 17997 4380
rect 17997 4324 18053 4380
rect 18053 4324 18057 4380
rect 17993 4320 18057 4324
rect 18073 4380 18137 4384
rect 18073 4324 18077 4380
rect 18077 4324 18133 4380
rect 18133 4324 18137 4380
rect 18073 4320 18137 4324
rect 26274 4380 26338 4384
rect 26274 4324 26278 4380
rect 26278 4324 26334 4380
rect 26334 4324 26338 4380
rect 26274 4320 26338 4324
rect 26354 4380 26418 4384
rect 26354 4324 26358 4380
rect 26358 4324 26414 4380
rect 26414 4324 26418 4380
rect 26354 4320 26418 4324
rect 26434 4380 26498 4384
rect 26434 4324 26438 4380
rect 26438 4324 26494 4380
rect 26494 4324 26498 4380
rect 26434 4320 26498 4324
rect 26514 4380 26578 4384
rect 26514 4324 26518 4380
rect 26518 4324 26574 4380
rect 26574 4324 26578 4380
rect 26514 4320 26578 4324
rect 34715 4380 34779 4384
rect 34715 4324 34719 4380
rect 34719 4324 34775 4380
rect 34775 4324 34779 4380
rect 34715 4320 34779 4324
rect 34795 4380 34859 4384
rect 34795 4324 34799 4380
rect 34799 4324 34855 4380
rect 34855 4324 34859 4380
rect 34795 4320 34859 4324
rect 34875 4380 34939 4384
rect 34875 4324 34879 4380
rect 34879 4324 34935 4380
rect 34935 4324 34939 4380
rect 34875 4320 34939 4324
rect 34955 4380 35019 4384
rect 34955 4324 34959 4380
rect 34959 4324 35015 4380
rect 35015 4324 35019 4380
rect 34955 4320 35019 4324
rect 5172 3836 5236 3840
rect 5172 3780 5176 3836
rect 5176 3780 5232 3836
rect 5232 3780 5236 3836
rect 5172 3776 5236 3780
rect 5252 3836 5316 3840
rect 5252 3780 5256 3836
rect 5256 3780 5312 3836
rect 5312 3780 5316 3836
rect 5252 3776 5316 3780
rect 5332 3836 5396 3840
rect 5332 3780 5336 3836
rect 5336 3780 5392 3836
rect 5392 3780 5396 3836
rect 5332 3776 5396 3780
rect 5412 3836 5476 3840
rect 5412 3780 5416 3836
rect 5416 3780 5472 3836
rect 5472 3780 5476 3836
rect 5412 3776 5476 3780
rect 13613 3836 13677 3840
rect 13613 3780 13617 3836
rect 13617 3780 13673 3836
rect 13673 3780 13677 3836
rect 13613 3776 13677 3780
rect 13693 3836 13757 3840
rect 13693 3780 13697 3836
rect 13697 3780 13753 3836
rect 13753 3780 13757 3836
rect 13693 3776 13757 3780
rect 13773 3836 13837 3840
rect 13773 3780 13777 3836
rect 13777 3780 13833 3836
rect 13833 3780 13837 3836
rect 13773 3776 13837 3780
rect 13853 3836 13917 3840
rect 13853 3780 13857 3836
rect 13857 3780 13913 3836
rect 13913 3780 13917 3836
rect 13853 3776 13917 3780
rect 22054 3836 22118 3840
rect 22054 3780 22058 3836
rect 22058 3780 22114 3836
rect 22114 3780 22118 3836
rect 22054 3776 22118 3780
rect 22134 3836 22198 3840
rect 22134 3780 22138 3836
rect 22138 3780 22194 3836
rect 22194 3780 22198 3836
rect 22134 3776 22198 3780
rect 22214 3836 22278 3840
rect 22214 3780 22218 3836
rect 22218 3780 22274 3836
rect 22274 3780 22278 3836
rect 22214 3776 22278 3780
rect 22294 3836 22358 3840
rect 22294 3780 22298 3836
rect 22298 3780 22354 3836
rect 22354 3780 22358 3836
rect 22294 3776 22358 3780
rect 30495 3836 30559 3840
rect 30495 3780 30499 3836
rect 30499 3780 30555 3836
rect 30555 3780 30559 3836
rect 30495 3776 30559 3780
rect 30575 3836 30639 3840
rect 30575 3780 30579 3836
rect 30579 3780 30635 3836
rect 30635 3780 30639 3836
rect 30575 3776 30639 3780
rect 30655 3836 30719 3840
rect 30655 3780 30659 3836
rect 30659 3780 30715 3836
rect 30715 3780 30719 3836
rect 30655 3776 30719 3780
rect 30735 3836 30799 3840
rect 30735 3780 30739 3836
rect 30739 3780 30795 3836
rect 30795 3780 30799 3836
rect 30735 3776 30799 3780
rect 9392 3292 9456 3296
rect 9392 3236 9396 3292
rect 9396 3236 9452 3292
rect 9452 3236 9456 3292
rect 9392 3232 9456 3236
rect 9472 3292 9536 3296
rect 9472 3236 9476 3292
rect 9476 3236 9532 3292
rect 9532 3236 9536 3292
rect 9472 3232 9536 3236
rect 9552 3292 9616 3296
rect 9552 3236 9556 3292
rect 9556 3236 9612 3292
rect 9612 3236 9616 3292
rect 9552 3232 9616 3236
rect 9632 3292 9696 3296
rect 9632 3236 9636 3292
rect 9636 3236 9692 3292
rect 9692 3236 9696 3292
rect 9632 3232 9696 3236
rect 17833 3292 17897 3296
rect 17833 3236 17837 3292
rect 17837 3236 17893 3292
rect 17893 3236 17897 3292
rect 17833 3232 17897 3236
rect 17913 3292 17977 3296
rect 17913 3236 17917 3292
rect 17917 3236 17973 3292
rect 17973 3236 17977 3292
rect 17913 3232 17977 3236
rect 17993 3292 18057 3296
rect 17993 3236 17997 3292
rect 17997 3236 18053 3292
rect 18053 3236 18057 3292
rect 17993 3232 18057 3236
rect 18073 3292 18137 3296
rect 18073 3236 18077 3292
rect 18077 3236 18133 3292
rect 18133 3236 18137 3292
rect 18073 3232 18137 3236
rect 26274 3292 26338 3296
rect 26274 3236 26278 3292
rect 26278 3236 26334 3292
rect 26334 3236 26338 3292
rect 26274 3232 26338 3236
rect 26354 3292 26418 3296
rect 26354 3236 26358 3292
rect 26358 3236 26414 3292
rect 26414 3236 26418 3292
rect 26354 3232 26418 3236
rect 26434 3292 26498 3296
rect 26434 3236 26438 3292
rect 26438 3236 26494 3292
rect 26494 3236 26498 3292
rect 26434 3232 26498 3236
rect 26514 3292 26578 3296
rect 26514 3236 26518 3292
rect 26518 3236 26574 3292
rect 26574 3236 26578 3292
rect 26514 3232 26578 3236
rect 34715 3292 34779 3296
rect 34715 3236 34719 3292
rect 34719 3236 34775 3292
rect 34775 3236 34779 3292
rect 34715 3232 34779 3236
rect 34795 3292 34859 3296
rect 34795 3236 34799 3292
rect 34799 3236 34855 3292
rect 34855 3236 34859 3292
rect 34795 3232 34859 3236
rect 34875 3292 34939 3296
rect 34875 3236 34879 3292
rect 34879 3236 34935 3292
rect 34935 3236 34939 3292
rect 34875 3232 34939 3236
rect 34955 3292 35019 3296
rect 34955 3236 34959 3292
rect 34959 3236 35015 3292
rect 35015 3236 35019 3292
rect 34955 3232 35019 3236
rect 5172 2748 5236 2752
rect 5172 2692 5176 2748
rect 5176 2692 5232 2748
rect 5232 2692 5236 2748
rect 5172 2688 5236 2692
rect 5252 2748 5316 2752
rect 5252 2692 5256 2748
rect 5256 2692 5312 2748
rect 5312 2692 5316 2748
rect 5252 2688 5316 2692
rect 5332 2748 5396 2752
rect 5332 2692 5336 2748
rect 5336 2692 5392 2748
rect 5392 2692 5396 2748
rect 5332 2688 5396 2692
rect 5412 2748 5476 2752
rect 5412 2692 5416 2748
rect 5416 2692 5472 2748
rect 5472 2692 5476 2748
rect 5412 2688 5476 2692
rect 13613 2748 13677 2752
rect 13613 2692 13617 2748
rect 13617 2692 13673 2748
rect 13673 2692 13677 2748
rect 13613 2688 13677 2692
rect 13693 2748 13757 2752
rect 13693 2692 13697 2748
rect 13697 2692 13753 2748
rect 13753 2692 13757 2748
rect 13693 2688 13757 2692
rect 13773 2748 13837 2752
rect 13773 2692 13777 2748
rect 13777 2692 13833 2748
rect 13833 2692 13837 2748
rect 13773 2688 13837 2692
rect 13853 2748 13917 2752
rect 13853 2692 13857 2748
rect 13857 2692 13913 2748
rect 13913 2692 13917 2748
rect 13853 2688 13917 2692
rect 22054 2748 22118 2752
rect 22054 2692 22058 2748
rect 22058 2692 22114 2748
rect 22114 2692 22118 2748
rect 22054 2688 22118 2692
rect 22134 2748 22198 2752
rect 22134 2692 22138 2748
rect 22138 2692 22194 2748
rect 22194 2692 22198 2748
rect 22134 2688 22198 2692
rect 22214 2748 22278 2752
rect 22214 2692 22218 2748
rect 22218 2692 22274 2748
rect 22274 2692 22278 2748
rect 22214 2688 22278 2692
rect 22294 2748 22358 2752
rect 22294 2692 22298 2748
rect 22298 2692 22354 2748
rect 22354 2692 22358 2748
rect 22294 2688 22358 2692
rect 30495 2748 30559 2752
rect 30495 2692 30499 2748
rect 30499 2692 30555 2748
rect 30555 2692 30559 2748
rect 30495 2688 30559 2692
rect 30575 2748 30639 2752
rect 30575 2692 30579 2748
rect 30579 2692 30635 2748
rect 30635 2692 30639 2748
rect 30575 2688 30639 2692
rect 30655 2748 30719 2752
rect 30655 2692 30659 2748
rect 30659 2692 30715 2748
rect 30715 2692 30719 2748
rect 30655 2688 30719 2692
rect 30735 2748 30799 2752
rect 30735 2692 30739 2748
rect 30739 2692 30795 2748
rect 30795 2692 30799 2748
rect 30735 2688 30799 2692
rect 9392 2204 9456 2208
rect 9392 2148 9396 2204
rect 9396 2148 9452 2204
rect 9452 2148 9456 2204
rect 9392 2144 9456 2148
rect 9472 2204 9536 2208
rect 9472 2148 9476 2204
rect 9476 2148 9532 2204
rect 9532 2148 9536 2204
rect 9472 2144 9536 2148
rect 9552 2204 9616 2208
rect 9552 2148 9556 2204
rect 9556 2148 9612 2204
rect 9612 2148 9616 2204
rect 9552 2144 9616 2148
rect 9632 2204 9696 2208
rect 9632 2148 9636 2204
rect 9636 2148 9692 2204
rect 9692 2148 9696 2204
rect 9632 2144 9696 2148
rect 17833 2204 17897 2208
rect 17833 2148 17837 2204
rect 17837 2148 17893 2204
rect 17893 2148 17897 2204
rect 17833 2144 17897 2148
rect 17913 2204 17977 2208
rect 17913 2148 17917 2204
rect 17917 2148 17973 2204
rect 17973 2148 17977 2204
rect 17913 2144 17977 2148
rect 17993 2204 18057 2208
rect 17993 2148 17997 2204
rect 17997 2148 18053 2204
rect 18053 2148 18057 2204
rect 17993 2144 18057 2148
rect 18073 2204 18137 2208
rect 18073 2148 18077 2204
rect 18077 2148 18133 2204
rect 18133 2148 18137 2204
rect 18073 2144 18137 2148
rect 26274 2204 26338 2208
rect 26274 2148 26278 2204
rect 26278 2148 26334 2204
rect 26334 2148 26338 2204
rect 26274 2144 26338 2148
rect 26354 2204 26418 2208
rect 26354 2148 26358 2204
rect 26358 2148 26414 2204
rect 26414 2148 26418 2204
rect 26354 2144 26418 2148
rect 26434 2204 26498 2208
rect 26434 2148 26438 2204
rect 26438 2148 26494 2204
rect 26494 2148 26498 2204
rect 26434 2144 26498 2148
rect 26514 2204 26578 2208
rect 26514 2148 26518 2204
rect 26518 2148 26574 2204
rect 26574 2148 26578 2204
rect 26514 2144 26578 2148
rect 34715 2204 34779 2208
rect 34715 2148 34719 2204
rect 34719 2148 34775 2204
rect 34775 2148 34779 2204
rect 34715 2144 34779 2148
rect 34795 2204 34859 2208
rect 34795 2148 34799 2204
rect 34799 2148 34855 2204
rect 34855 2148 34859 2204
rect 34795 2144 34859 2148
rect 34875 2204 34939 2208
rect 34875 2148 34879 2204
rect 34879 2148 34935 2204
rect 34935 2148 34939 2204
rect 34875 2144 34939 2148
rect 34955 2204 35019 2208
rect 34955 2148 34959 2204
rect 34959 2148 35015 2204
rect 35015 2148 35019 2204
rect 34955 2144 35019 2148
<< metal4 >>
rect 5164 39744 5484 39760
rect 5164 39680 5172 39744
rect 5236 39680 5252 39744
rect 5316 39680 5332 39744
rect 5396 39680 5412 39744
rect 5476 39680 5484 39744
rect 5164 38656 5484 39680
rect 5164 38592 5172 38656
rect 5236 38592 5252 38656
rect 5316 38592 5332 38656
rect 5396 38592 5412 38656
rect 5476 38592 5484 38656
rect 5164 37568 5484 38592
rect 5164 37504 5172 37568
rect 5236 37504 5252 37568
rect 5316 37504 5332 37568
rect 5396 37504 5412 37568
rect 5476 37504 5484 37568
rect 5164 36480 5484 37504
rect 5164 36416 5172 36480
rect 5236 36416 5252 36480
rect 5316 36416 5332 36480
rect 5396 36416 5412 36480
rect 5476 36416 5484 36480
rect 5164 35392 5484 36416
rect 5164 35328 5172 35392
rect 5236 35328 5252 35392
rect 5316 35328 5332 35392
rect 5396 35328 5412 35392
rect 5476 35328 5484 35392
rect 5164 34304 5484 35328
rect 5164 34240 5172 34304
rect 5236 34240 5252 34304
rect 5316 34240 5332 34304
rect 5396 34240 5412 34304
rect 5476 34240 5484 34304
rect 5164 33216 5484 34240
rect 5164 33152 5172 33216
rect 5236 33152 5252 33216
rect 5316 33152 5332 33216
rect 5396 33152 5412 33216
rect 5476 33152 5484 33216
rect 5164 32128 5484 33152
rect 5164 32064 5172 32128
rect 5236 32064 5252 32128
rect 5316 32064 5332 32128
rect 5396 32064 5412 32128
rect 5476 32064 5484 32128
rect 5164 31040 5484 32064
rect 5164 30976 5172 31040
rect 5236 30976 5252 31040
rect 5316 30976 5332 31040
rect 5396 30976 5412 31040
rect 5476 30976 5484 31040
rect 5164 29952 5484 30976
rect 5164 29888 5172 29952
rect 5236 29888 5252 29952
rect 5316 29888 5332 29952
rect 5396 29888 5412 29952
rect 5476 29888 5484 29952
rect 5164 28864 5484 29888
rect 5164 28800 5172 28864
rect 5236 28800 5252 28864
rect 5316 28800 5332 28864
rect 5396 28800 5412 28864
rect 5476 28800 5484 28864
rect 5164 27776 5484 28800
rect 5164 27712 5172 27776
rect 5236 27712 5252 27776
rect 5316 27712 5332 27776
rect 5396 27712 5412 27776
rect 5476 27712 5484 27776
rect 5164 26688 5484 27712
rect 5164 26624 5172 26688
rect 5236 26624 5252 26688
rect 5316 26624 5332 26688
rect 5396 26624 5412 26688
rect 5476 26624 5484 26688
rect 5164 25600 5484 26624
rect 5164 25536 5172 25600
rect 5236 25536 5252 25600
rect 5316 25536 5332 25600
rect 5396 25536 5412 25600
rect 5476 25536 5484 25600
rect 5164 24512 5484 25536
rect 5164 24448 5172 24512
rect 5236 24448 5252 24512
rect 5316 24448 5332 24512
rect 5396 24448 5412 24512
rect 5476 24448 5484 24512
rect 5164 23424 5484 24448
rect 5164 23360 5172 23424
rect 5236 23360 5252 23424
rect 5316 23360 5332 23424
rect 5396 23360 5412 23424
rect 5476 23360 5484 23424
rect 5164 22336 5484 23360
rect 5164 22272 5172 22336
rect 5236 22272 5252 22336
rect 5316 22272 5332 22336
rect 5396 22272 5412 22336
rect 5476 22272 5484 22336
rect 5164 21248 5484 22272
rect 5164 21184 5172 21248
rect 5236 21184 5252 21248
rect 5316 21184 5332 21248
rect 5396 21184 5412 21248
rect 5476 21184 5484 21248
rect 5164 20160 5484 21184
rect 5164 20096 5172 20160
rect 5236 20096 5252 20160
rect 5316 20096 5332 20160
rect 5396 20096 5412 20160
rect 5476 20096 5484 20160
rect 5164 19072 5484 20096
rect 5164 19008 5172 19072
rect 5236 19008 5252 19072
rect 5316 19008 5332 19072
rect 5396 19008 5412 19072
rect 5476 19008 5484 19072
rect 5164 17984 5484 19008
rect 5164 17920 5172 17984
rect 5236 17920 5252 17984
rect 5316 17920 5332 17984
rect 5396 17920 5412 17984
rect 5476 17920 5484 17984
rect 5164 16896 5484 17920
rect 5164 16832 5172 16896
rect 5236 16832 5252 16896
rect 5316 16832 5332 16896
rect 5396 16832 5412 16896
rect 5476 16832 5484 16896
rect 5164 15808 5484 16832
rect 5164 15744 5172 15808
rect 5236 15744 5252 15808
rect 5316 15744 5332 15808
rect 5396 15744 5412 15808
rect 5476 15744 5484 15808
rect 5164 14720 5484 15744
rect 5164 14656 5172 14720
rect 5236 14656 5252 14720
rect 5316 14656 5332 14720
rect 5396 14656 5412 14720
rect 5476 14656 5484 14720
rect 5164 13632 5484 14656
rect 5164 13568 5172 13632
rect 5236 13568 5252 13632
rect 5316 13568 5332 13632
rect 5396 13568 5412 13632
rect 5476 13568 5484 13632
rect 5164 12544 5484 13568
rect 5164 12480 5172 12544
rect 5236 12480 5252 12544
rect 5316 12480 5332 12544
rect 5396 12480 5412 12544
rect 5476 12480 5484 12544
rect 5164 11456 5484 12480
rect 5164 11392 5172 11456
rect 5236 11392 5252 11456
rect 5316 11392 5332 11456
rect 5396 11392 5412 11456
rect 5476 11392 5484 11456
rect 5164 10368 5484 11392
rect 5164 10304 5172 10368
rect 5236 10304 5252 10368
rect 5316 10304 5332 10368
rect 5396 10304 5412 10368
rect 5476 10304 5484 10368
rect 5164 9280 5484 10304
rect 5164 9216 5172 9280
rect 5236 9216 5252 9280
rect 5316 9216 5332 9280
rect 5396 9216 5412 9280
rect 5476 9216 5484 9280
rect 5164 8192 5484 9216
rect 5164 8128 5172 8192
rect 5236 8128 5252 8192
rect 5316 8128 5332 8192
rect 5396 8128 5412 8192
rect 5476 8128 5484 8192
rect 5164 7104 5484 8128
rect 5164 7040 5172 7104
rect 5236 7040 5252 7104
rect 5316 7040 5332 7104
rect 5396 7040 5412 7104
rect 5476 7040 5484 7104
rect 5164 6016 5484 7040
rect 5164 5952 5172 6016
rect 5236 5952 5252 6016
rect 5316 5952 5332 6016
rect 5396 5952 5412 6016
rect 5476 5952 5484 6016
rect 5164 4928 5484 5952
rect 5164 4864 5172 4928
rect 5236 4864 5252 4928
rect 5316 4864 5332 4928
rect 5396 4864 5412 4928
rect 5476 4864 5484 4928
rect 5164 3840 5484 4864
rect 5164 3776 5172 3840
rect 5236 3776 5252 3840
rect 5316 3776 5332 3840
rect 5396 3776 5412 3840
rect 5476 3776 5484 3840
rect 5164 2752 5484 3776
rect 5164 2688 5172 2752
rect 5236 2688 5252 2752
rect 5316 2688 5332 2752
rect 5396 2688 5412 2752
rect 5476 2688 5484 2752
rect 5164 2128 5484 2688
rect 9384 39200 9704 39760
rect 9384 39136 9392 39200
rect 9456 39136 9472 39200
rect 9536 39136 9552 39200
rect 9616 39136 9632 39200
rect 9696 39136 9704 39200
rect 9384 38112 9704 39136
rect 9384 38048 9392 38112
rect 9456 38048 9472 38112
rect 9536 38048 9552 38112
rect 9616 38048 9632 38112
rect 9696 38048 9704 38112
rect 9384 37024 9704 38048
rect 9384 36960 9392 37024
rect 9456 36960 9472 37024
rect 9536 36960 9552 37024
rect 9616 36960 9632 37024
rect 9696 36960 9704 37024
rect 9384 35936 9704 36960
rect 9384 35872 9392 35936
rect 9456 35872 9472 35936
rect 9536 35872 9552 35936
rect 9616 35872 9632 35936
rect 9696 35872 9704 35936
rect 9384 34848 9704 35872
rect 9384 34784 9392 34848
rect 9456 34784 9472 34848
rect 9536 34784 9552 34848
rect 9616 34784 9632 34848
rect 9696 34784 9704 34848
rect 9384 33760 9704 34784
rect 9384 33696 9392 33760
rect 9456 33696 9472 33760
rect 9536 33696 9552 33760
rect 9616 33696 9632 33760
rect 9696 33696 9704 33760
rect 9384 32672 9704 33696
rect 9384 32608 9392 32672
rect 9456 32608 9472 32672
rect 9536 32608 9552 32672
rect 9616 32608 9632 32672
rect 9696 32608 9704 32672
rect 9384 31584 9704 32608
rect 9384 31520 9392 31584
rect 9456 31520 9472 31584
rect 9536 31520 9552 31584
rect 9616 31520 9632 31584
rect 9696 31520 9704 31584
rect 9384 30496 9704 31520
rect 9384 30432 9392 30496
rect 9456 30432 9472 30496
rect 9536 30432 9552 30496
rect 9616 30432 9632 30496
rect 9696 30432 9704 30496
rect 9384 29408 9704 30432
rect 9384 29344 9392 29408
rect 9456 29344 9472 29408
rect 9536 29344 9552 29408
rect 9616 29344 9632 29408
rect 9696 29344 9704 29408
rect 9384 28320 9704 29344
rect 9384 28256 9392 28320
rect 9456 28256 9472 28320
rect 9536 28256 9552 28320
rect 9616 28256 9632 28320
rect 9696 28256 9704 28320
rect 9384 27232 9704 28256
rect 9384 27168 9392 27232
rect 9456 27168 9472 27232
rect 9536 27168 9552 27232
rect 9616 27168 9632 27232
rect 9696 27168 9704 27232
rect 9384 26144 9704 27168
rect 9384 26080 9392 26144
rect 9456 26080 9472 26144
rect 9536 26080 9552 26144
rect 9616 26080 9632 26144
rect 9696 26080 9704 26144
rect 9384 25056 9704 26080
rect 9384 24992 9392 25056
rect 9456 24992 9472 25056
rect 9536 24992 9552 25056
rect 9616 24992 9632 25056
rect 9696 24992 9704 25056
rect 9384 23968 9704 24992
rect 9384 23904 9392 23968
rect 9456 23904 9472 23968
rect 9536 23904 9552 23968
rect 9616 23904 9632 23968
rect 9696 23904 9704 23968
rect 9384 22880 9704 23904
rect 9384 22816 9392 22880
rect 9456 22816 9472 22880
rect 9536 22816 9552 22880
rect 9616 22816 9632 22880
rect 9696 22816 9704 22880
rect 9384 21792 9704 22816
rect 9384 21728 9392 21792
rect 9456 21728 9472 21792
rect 9536 21728 9552 21792
rect 9616 21728 9632 21792
rect 9696 21728 9704 21792
rect 9384 20704 9704 21728
rect 9384 20640 9392 20704
rect 9456 20640 9472 20704
rect 9536 20640 9552 20704
rect 9616 20640 9632 20704
rect 9696 20640 9704 20704
rect 9384 19616 9704 20640
rect 9384 19552 9392 19616
rect 9456 19552 9472 19616
rect 9536 19552 9552 19616
rect 9616 19552 9632 19616
rect 9696 19552 9704 19616
rect 9384 18528 9704 19552
rect 9384 18464 9392 18528
rect 9456 18464 9472 18528
rect 9536 18464 9552 18528
rect 9616 18464 9632 18528
rect 9696 18464 9704 18528
rect 9384 17440 9704 18464
rect 9384 17376 9392 17440
rect 9456 17376 9472 17440
rect 9536 17376 9552 17440
rect 9616 17376 9632 17440
rect 9696 17376 9704 17440
rect 9384 16352 9704 17376
rect 9384 16288 9392 16352
rect 9456 16288 9472 16352
rect 9536 16288 9552 16352
rect 9616 16288 9632 16352
rect 9696 16288 9704 16352
rect 9384 15264 9704 16288
rect 9384 15200 9392 15264
rect 9456 15200 9472 15264
rect 9536 15200 9552 15264
rect 9616 15200 9632 15264
rect 9696 15200 9704 15264
rect 9384 14176 9704 15200
rect 9384 14112 9392 14176
rect 9456 14112 9472 14176
rect 9536 14112 9552 14176
rect 9616 14112 9632 14176
rect 9696 14112 9704 14176
rect 9384 13088 9704 14112
rect 9384 13024 9392 13088
rect 9456 13024 9472 13088
rect 9536 13024 9552 13088
rect 9616 13024 9632 13088
rect 9696 13024 9704 13088
rect 9384 12000 9704 13024
rect 9384 11936 9392 12000
rect 9456 11936 9472 12000
rect 9536 11936 9552 12000
rect 9616 11936 9632 12000
rect 9696 11936 9704 12000
rect 9384 10912 9704 11936
rect 9384 10848 9392 10912
rect 9456 10848 9472 10912
rect 9536 10848 9552 10912
rect 9616 10848 9632 10912
rect 9696 10848 9704 10912
rect 9384 9824 9704 10848
rect 9384 9760 9392 9824
rect 9456 9760 9472 9824
rect 9536 9760 9552 9824
rect 9616 9760 9632 9824
rect 9696 9760 9704 9824
rect 9384 8736 9704 9760
rect 9384 8672 9392 8736
rect 9456 8672 9472 8736
rect 9536 8672 9552 8736
rect 9616 8672 9632 8736
rect 9696 8672 9704 8736
rect 9384 7648 9704 8672
rect 9384 7584 9392 7648
rect 9456 7584 9472 7648
rect 9536 7584 9552 7648
rect 9616 7584 9632 7648
rect 9696 7584 9704 7648
rect 9384 6560 9704 7584
rect 9384 6496 9392 6560
rect 9456 6496 9472 6560
rect 9536 6496 9552 6560
rect 9616 6496 9632 6560
rect 9696 6496 9704 6560
rect 9384 5472 9704 6496
rect 9384 5408 9392 5472
rect 9456 5408 9472 5472
rect 9536 5408 9552 5472
rect 9616 5408 9632 5472
rect 9696 5408 9704 5472
rect 9384 4384 9704 5408
rect 9384 4320 9392 4384
rect 9456 4320 9472 4384
rect 9536 4320 9552 4384
rect 9616 4320 9632 4384
rect 9696 4320 9704 4384
rect 9384 3296 9704 4320
rect 9384 3232 9392 3296
rect 9456 3232 9472 3296
rect 9536 3232 9552 3296
rect 9616 3232 9632 3296
rect 9696 3232 9704 3296
rect 9384 2208 9704 3232
rect 9384 2144 9392 2208
rect 9456 2144 9472 2208
rect 9536 2144 9552 2208
rect 9616 2144 9632 2208
rect 9696 2144 9704 2208
rect 9384 2128 9704 2144
rect 13605 39744 13925 39760
rect 13605 39680 13613 39744
rect 13677 39680 13693 39744
rect 13757 39680 13773 39744
rect 13837 39680 13853 39744
rect 13917 39680 13925 39744
rect 13605 38656 13925 39680
rect 13605 38592 13613 38656
rect 13677 38592 13693 38656
rect 13757 38592 13773 38656
rect 13837 38592 13853 38656
rect 13917 38592 13925 38656
rect 13605 37568 13925 38592
rect 13605 37504 13613 37568
rect 13677 37504 13693 37568
rect 13757 37504 13773 37568
rect 13837 37504 13853 37568
rect 13917 37504 13925 37568
rect 13605 36480 13925 37504
rect 13605 36416 13613 36480
rect 13677 36416 13693 36480
rect 13757 36416 13773 36480
rect 13837 36416 13853 36480
rect 13917 36416 13925 36480
rect 13605 35392 13925 36416
rect 13605 35328 13613 35392
rect 13677 35328 13693 35392
rect 13757 35328 13773 35392
rect 13837 35328 13853 35392
rect 13917 35328 13925 35392
rect 13605 34304 13925 35328
rect 13605 34240 13613 34304
rect 13677 34240 13693 34304
rect 13757 34240 13773 34304
rect 13837 34240 13853 34304
rect 13917 34240 13925 34304
rect 13605 33216 13925 34240
rect 13605 33152 13613 33216
rect 13677 33152 13693 33216
rect 13757 33152 13773 33216
rect 13837 33152 13853 33216
rect 13917 33152 13925 33216
rect 13605 32128 13925 33152
rect 13605 32064 13613 32128
rect 13677 32064 13693 32128
rect 13757 32064 13773 32128
rect 13837 32064 13853 32128
rect 13917 32064 13925 32128
rect 13605 31040 13925 32064
rect 13605 30976 13613 31040
rect 13677 30976 13693 31040
rect 13757 30976 13773 31040
rect 13837 30976 13853 31040
rect 13917 30976 13925 31040
rect 13605 29952 13925 30976
rect 13605 29888 13613 29952
rect 13677 29888 13693 29952
rect 13757 29888 13773 29952
rect 13837 29888 13853 29952
rect 13917 29888 13925 29952
rect 13605 28864 13925 29888
rect 13605 28800 13613 28864
rect 13677 28800 13693 28864
rect 13757 28800 13773 28864
rect 13837 28800 13853 28864
rect 13917 28800 13925 28864
rect 13605 27776 13925 28800
rect 13605 27712 13613 27776
rect 13677 27712 13693 27776
rect 13757 27712 13773 27776
rect 13837 27712 13853 27776
rect 13917 27712 13925 27776
rect 13605 26688 13925 27712
rect 13605 26624 13613 26688
rect 13677 26624 13693 26688
rect 13757 26624 13773 26688
rect 13837 26624 13853 26688
rect 13917 26624 13925 26688
rect 13605 25600 13925 26624
rect 13605 25536 13613 25600
rect 13677 25536 13693 25600
rect 13757 25536 13773 25600
rect 13837 25536 13853 25600
rect 13917 25536 13925 25600
rect 13605 24512 13925 25536
rect 13605 24448 13613 24512
rect 13677 24448 13693 24512
rect 13757 24448 13773 24512
rect 13837 24448 13853 24512
rect 13917 24448 13925 24512
rect 13605 23424 13925 24448
rect 13605 23360 13613 23424
rect 13677 23360 13693 23424
rect 13757 23360 13773 23424
rect 13837 23360 13853 23424
rect 13917 23360 13925 23424
rect 13605 22336 13925 23360
rect 13605 22272 13613 22336
rect 13677 22272 13693 22336
rect 13757 22272 13773 22336
rect 13837 22272 13853 22336
rect 13917 22272 13925 22336
rect 13605 21248 13925 22272
rect 13605 21184 13613 21248
rect 13677 21184 13693 21248
rect 13757 21184 13773 21248
rect 13837 21184 13853 21248
rect 13917 21184 13925 21248
rect 13605 20160 13925 21184
rect 13605 20096 13613 20160
rect 13677 20096 13693 20160
rect 13757 20096 13773 20160
rect 13837 20096 13853 20160
rect 13917 20096 13925 20160
rect 13605 19072 13925 20096
rect 13605 19008 13613 19072
rect 13677 19008 13693 19072
rect 13757 19008 13773 19072
rect 13837 19008 13853 19072
rect 13917 19008 13925 19072
rect 13605 17984 13925 19008
rect 13605 17920 13613 17984
rect 13677 17920 13693 17984
rect 13757 17920 13773 17984
rect 13837 17920 13853 17984
rect 13917 17920 13925 17984
rect 13605 16896 13925 17920
rect 13605 16832 13613 16896
rect 13677 16832 13693 16896
rect 13757 16832 13773 16896
rect 13837 16832 13853 16896
rect 13917 16832 13925 16896
rect 13605 15808 13925 16832
rect 13605 15744 13613 15808
rect 13677 15744 13693 15808
rect 13757 15744 13773 15808
rect 13837 15744 13853 15808
rect 13917 15744 13925 15808
rect 13605 14720 13925 15744
rect 13605 14656 13613 14720
rect 13677 14656 13693 14720
rect 13757 14656 13773 14720
rect 13837 14656 13853 14720
rect 13917 14656 13925 14720
rect 13605 13632 13925 14656
rect 13605 13568 13613 13632
rect 13677 13568 13693 13632
rect 13757 13568 13773 13632
rect 13837 13568 13853 13632
rect 13917 13568 13925 13632
rect 13605 12544 13925 13568
rect 13605 12480 13613 12544
rect 13677 12480 13693 12544
rect 13757 12480 13773 12544
rect 13837 12480 13853 12544
rect 13917 12480 13925 12544
rect 13605 11456 13925 12480
rect 13605 11392 13613 11456
rect 13677 11392 13693 11456
rect 13757 11392 13773 11456
rect 13837 11392 13853 11456
rect 13917 11392 13925 11456
rect 13605 10368 13925 11392
rect 13605 10304 13613 10368
rect 13677 10304 13693 10368
rect 13757 10304 13773 10368
rect 13837 10304 13853 10368
rect 13917 10304 13925 10368
rect 13605 9280 13925 10304
rect 13605 9216 13613 9280
rect 13677 9216 13693 9280
rect 13757 9216 13773 9280
rect 13837 9216 13853 9280
rect 13917 9216 13925 9280
rect 13605 8192 13925 9216
rect 13605 8128 13613 8192
rect 13677 8128 13693 8192
rect 13757 8128 13773 8192
rect 13837 8128 13853 8192
rect 13917 8128 13925 8192
rect 13605 7104 13925 8128
rect 13605 7040 13613 7104
rect 13677 7040 13693 7104
rect 13757 7040 13773 7104
rect 13837 7040 13853 7104
rect 13917 7040 13925 7104
rect 13605 6016 13925 7040
rect 13605 5952 13613 6016
rect 13677 5952 13693 6016
rect 13757 5952 13773 6016
rect 13837 5952 13853 6016
rect 13917 5952 13925 6016
rect 13605 4928 13925 5952
rect 13605 4864 13613 4928
rect 13677 4864 13693 4928
rect 13757 4864 13773 4928
rect 13837 4864 13853 4928
rect 13917 4864 13925 4928
rect 13605 3840 13925 4864
rect 13605 3776 13613 3840
rect 13677 3776 13693 3840
rect 13757 3776 13773 3840
rect 13837 3776 13853 3840
rect 13917 3776 13925 3840
rect 13605 2752 13925 3776
rect 13605 2688 13613 2752
rect 13677 2688 13693 2752
rect 13757 2688 13773 2752
rect 13837 2688 13853 2752
rect 13917 2688 13925 2752
rect 13605 2128 13925 2688
rect 17825 39200 18145 39760
rect 17825 39136 17833 39200
rect 17897 39136 17913 39200
rect 17977 39136 17993 39200
rect 18057 39136 18073 39200
rect 18137 39136 18145 39200
rect 17825 38112 18145 39136
rect 17825 38048 17833 38112
rect 17897 38048 17913 38112
rect 17977 38048 17993 38112
rect 18057 38048 18073 38112
rect 18137 38048 18145 38112
rect 17825 37024 18145 38048
rect 17825 36960 17833 37024
rect 17897 36960 17913 37024
rect 17977 36960 17993 37024
rect 18057 36960 18073 37024
rect 18137 36960 18145 37024
rect 17825 35936 18145 36960
rect 17825 35872 17833 35936
rect 17897 35872 17913 35936
rect 17977 35872 17993 35936
rect 18057 35872 18073 35936
rect 18137 35872 18145 35936
rect 17825 34848 18145 35872
rect 17825 34784 17833 34848
rect 17897 34784 17913 34848
rect 17977 34784 17993 34848
rect 18057 34784 18073 34848
rect 18137 34784 18145 34848
rect 17825 33760 18145 34784
rect 17825 33696 17833 33760
rect 17897 33696 17913 33760
rect 17977 33696 17993 33760
rect 18057 33696 18073 33760
rect 18137 33696 18145 33760
rect 17825 32672 18145 33696
rect 17825 32608 17833 32672
rect 17897 32608 17913 32672
rect 17977 32608 17993 32672
rect 18057 32608 18073 32672
rect 18137 32608 18145 32672
rect 17825 31584 18145 32608
rect 17825 31520 17833 31584
rect 17897 31520 17913 31584
rect 17977 31520 17993 31584
rect 18057 31520 18073 31584
rect 18137 31520 18145 31584
rect 17825 30496 18145 31520
rect 17825 30432 17833 30496
rect 17897 30432 17913 30496
rect 17977 30432 17993 30496
rect 18057 30432 18073 30496
rect 18137 30432 18145 30496
rect 17825 29408 18145 30432
rect 17825 29344 17833 29408
rect 17897 29344 17913 29408
rect 17977 29344 17993 29408
rect 18057 29344 18073 29408
rect 18137 29344 18145 29408
rect 17825 28320 18145 29344
rect 17825 28256 17833 28320
rect 17897 28256 17913 28320
rect 17977 28256 17993 28320
rect 18057 28256 18073 28320
rect 18137 28256 18145 28320
rect 17825 27232 18145 28256
rect 17825 27168 17833 27232
rect 17897 27168 17913 27232
rect 17977 27168 17993 27232
rect 18057 27168 18073 27232
rect 18137 27168 18145 27232
rect 17825 26144 18145 27168
rect 17825 26080 17833 26144
rect 17897 26080 17913 26144
rect 17977 26080 17993 26144
rect 18057 26080 18073 26144
rect 18137 26080 18145 26144
rect 17825 25056 18145 26080
rect 17825 24992 17833 25056
rect 17897 24992 17913 25056
rect 17977 24992 17993 25056
rect 18057 24992 18073 25056
rect 18137 24992 18145 25056
rect 17825 23968 18145 24992
rect 17825 23904 17833 23968
rect 17897 23904 17913 23968
rect 17977 23904 17993 23968
rect 18057 23904 18073 23968
rect 18137 23904 18145 23968
rect 17825 22880 18145 23904
rect 17825 22816 17833 22880
rect 17897 22816 17913 22880
rect 17977 22816 17993 22880
rect 18057 22816 18073 22880
rect 18137 22816 18145 22880
rect 17825 21792 18145 22816
rect 17825 21728 17833 21792
rect 17897 21728 17913 21792
rect 17977 21728 17993 21792
rect 18057 21728 18073 21792
rect 18137 21728 18145 21792
rect 17825 20704 18145 21728
rect 17825 20640 17833 20704
rect 17897 20640 17913 20704
rect 17977 20640 17993 20704
rect 18057 20640 18073 20704
rect 18137 20640 18145 20704
rect 17825 19616 18145 20640
rect 17825 19552 17833 19616
rect 17897 19552 17913 19616
rect 17977 19552 17993 19616
rect 18057 19552 18073 19616
rect 18137 19552 18145 19616
rect 17825 18528 18145 19552
rect 17825 18464 17833 18528
rect 17897 18464 17913 18528
rect 17977 18464 17993 18528
rect 18057 18464 18073 18528
rect 18137 18464 18145 18528
rect 17825 17440 18145 18464
rect 17825 17376 17833 17440
rect 17897 17376 17913 17440
rect 17977 17376 17993 17440
rect 18057 17376 18073 17440
rect 18137 17376 18145 17440
rect 17825 16352 18145 17376
rect 17825 16288 17833 16352
rect 17897 16288 17913 16352
rect 17977 16288 17993 16352
rect 18057 16288 18073 16352
rect 18137 16288 18145 16352
rect 17825 15264 18145 16288
rect 17825 15200 17833 15264
rect 17897 15200 17913 15264
rect 17977 15200 17993 15264
rect 18057 15200 18073 15264
rect 18137 15200 18145 15264
rect 17825 14176 18145 15200
rect 17825 14112 17833 14176
rect 17897 14112 17913 14176
rect 17977 14112 17993 14176
rect 18057 14112 18073 14176
rect 18137 14112 18145 14176
rect 17825 13088 18145 14112
rect 17825 13024 17833 13088
rect 17897 13024 17913 13088
rect 17977 13024 17993 13088
rect 18057 13024 18073 13088
rect 18137 13024 18145 13088
rect 17825 12000 18145 13024
rect 17825 11936 17833 12000
rect 17897 11936 17913 12000
rect 17977 11936 17993 12000
rect 18057 11936 18073 12000
rect 18137 11936 18145 12000
rect 17825 10912 18145 11936
rect 17825 10848 17833 10912
rect 17897 10848 17913 10912
rect 17977 10848 17993 10912
rect 18057 10848 18073 10912
rect 18137 10848 18145 10912
rect 17825 9824 18145 10848
rect 17825 9760 17833 9824
rect 17897 9760 17913 9824
rect 17977 9760 17993 9824
rect 18057 9760 18073 9824
rect 18137 9760 18145 9824
rect 17825 8736 18145 9760
rect 17825 8672 17833 8736
rect 17897 8672 17913 8736
rect 17977 8672 17993 8736
rect 18057 8672 18073 8736
rect 18137 8672 18145 8736
rect 17825 7648 18145 8672
rect 17825 7584 17833 7648
rect 17897 7584 17913 7648
rect 17977 7584 17993 7648
rect 18057 7584 18073 7648
rect 18137 7584 18145 7648
rect 17825 6560 18145 7584
rect 17825 6496 17833 6560
rect 17897 6496 17913 6560
rect 17977 6496 17993 6560
rect 18057 6496 18073 6560
rect 18137 6496 18145 6560
rect 17825 5472 18145 6496
rect 17825 5408 17833 5472
rect 17897 5408 17913 5472
rect 17977 5408 17993 5472
rect 18057 5408 18073 5472
rect 18137 5408 18145 5472
rect 17825 4384 18145 5408
rect 17825 4320 17833 4384
rect 17897 4320 17913 4384
rect 17977 4320 17993 4384
rect 18057 4320 18073 4384
rect 18137 4320 18145 4384
rect 17825 3296 18145 4320
rect 17825 3232 17833 3296
rect 17897 3232 17913 3296
rect 17977 3232 17993 3296
rect 18057 3232 18073 3296
rect 18137 3232 18145 3296
rect 17825 2208 18145 3232
rect 17825 2144 17833 2208
rect 17897 2144 17913 2208
rect 17977 2144 17993 2208
rect 18057 2144 18073 2208
rect 18137 2144 18145 2208
rect 17825 2128 18145 2144
rect 22046 39744 22366 39760
rect 22046 39680 22054 39744
rect 22118 39680 22134 39744
rect 22198 39680 22214 39744
rect 22278 39680 22294 39744
rect 22358 39680 22366 39744
rect 22046 38656 22366 39680
rect 22046 38592 22054 38656
rect 22118 38592 22134 38656
rect 22198 38592 22214 38656
rect 22278 38592 22294 38656
rect 22358 38592 22366 38656
rect 22046 37568 22366 38592
rect 22046 37504 22054 37568
rect 22118 37504 22134 37568
rect 22198 37504 22214 37568
rect 22278 37504 22294 37568
rect 22358 37504 22366 37568
rect 22046 36480 22366 37504
rect 22046 36416 22054 36480
rect 22118 36416 22134 36480
rect 22198 36416 22214 36480
rect 22278 36416 22294 36480
rect 22358 36416 22366 36480
rect 22046 35392 22366 36416
rect 22046 35328 22054 35392
rect 22118 35328 22134 35392
rect 22198 35328 22214 35392
rect 22278 35328 22294 35392
rect 22358 35328 22366 35392
rect 22046 34304 22366 35328
rect 22046 34240 22054 34304
rect 22118 34240 22134 34304
rect 22198 34240 22214 34304
rect 22278 34240 22294 34304
rect 22358 34240 22366 34304
rect 22046 33216 22366 34240
rect 22046 33152 22054 33216
rect 22118 33152 22134 33216
rect 22198 33152 22214 33216
rect 22278 33152 22294 33216
rect 22358 33152 22366 33216
rect 22046 32128 22366 33152
rect 22046 32064 22054 32128
rect 22118 32064 22134 32128
rect 22198 32064 22214 32128
rect 22278 32064 22294 32128
rect 22358 32064 22366 32128
rect 22046 31040 22366 32064
rect 22046 30976 22054 31040
rect 22118 30976 22134 31040
rect 22198 30976 22214 31040
rect 22278 30976 22294 31040
rect 22358 30976 22366 31040
rect 22046 29952 22366 30976
rect 22046 29888 22054 29952
rect 22118 29888 22134 29952
rect 22198 29888 22214 29952
rect 22278 29888 22294 29952
rect 22358 29888 22366 29952
rect 22046 28864 22366 29888
rect 22046 28800 22054 28864
rect 22118 28800 22134 28864
rect 22198 28800 22214 28864
rect 22278 28800 22294 28864
rect 22358 28800 22366 28864
rect 22046 27776 22366 28800
rect 22046 27712 22054 27776
rect 22118 27712 22134 27776
rect 22198 27712 22214 27776
rect 22278 27712 22294 27776
rect 22358 27712 22366 27776
rect 22046 26688 22366 27712
rect 22046 26624 22054 26688
rect 22118 26624 22134 26688
rect 22198 26624 22214 26688
rect 22278 26624 22294 26688
rect 22358 26624 22366 26688
rect 22046 25600 22366 26624
rect 22046 25536 22054 25600
rect 22118 25536 22134 25600
rect 22198 25536 22214 25600
rect 22278 25536 22294 25600
rect 22358 25536 22366 25600
rect 22046 24512 22366 25536
rect 22046 24448 22054 24512
rect 22118 24448 22134 24512
rect 22198 24448 22214 24512
rect 22278 24448 22294 24512
rect 22358 24448 22366 24512
rect 22046 23424 22366 24448
rect 22046 23360 22054 23424
rect 22118 23360 22134 23424
rect 22198 23360 22214 23424
rect 22278 23360 22294 23424
rect 22358 23360 22366 23424
rect 22046 22336 22366 23360
rect 22046 22272 22054 22336
rect 22118 22272 22134 22336
rect 22198 22272 22214 22336
rect 22278 22272 22294 22336
rect 22358 22272 22366 22336
rect 22046 21248 22366 22272
rect 22046 21184 22054 21248
rect 22118 21184 22134 21248
rect 22198 21184 22214 21248
rect 22278 21184 22294 21248
rect 22358 21184 22366 21248
rect 22046 20160 22366 21184
rect 22046 20096 22054 20160
rect 22118 20096 22134 20160
rect 22198 20096 22214 20160
rect 22278 20096 22294 20160
rect 22358 20096 22366 20160
rect 22046 19072 22366 20096
rect 22046 19008 22054 19072
rect 22118 19008 22134 19072
rect 22198 19008 22214 19072
rect 22278 19008 22294 19072
rect 22358 19008 22366 19072
rect 22046 17984 22366 19008
rect 22046 17920 22054 17984
rect 22118 17920 22134 17984
rect 22198 17920 22214 17984
rect 22278 17920 22294 17984
rect 22358 17920 22366 17984
rect 22046 16896 22366 17920
rect 22046 16832 22054 16896
rect 22118 16832 22134 16896
rect 22198 16832 22214 16896
rect 22278 16832 22294 16896
rect 22358 16832 22366 16896
rect 22046 15808 22366 16832
rect 22046 15744 22054 15808
rect 22118 15744 22134 15808
rect 22198 15744 22214 15808
rect 22278 15744 22294 15808
rect 22358 15744 22366 15808
rect 22046 14720 22366 15744
rect 22046 14656 22054 14720
rect 22118 14656 22134 14720
rect 22198 14656 22214 14720
rect 22278 14656 22294 14720
rect 22358 14656 22366 14720
rect 22046 13632 22366 14656
rect 22046 13568 22054 13632
rect 22118 13568 22134 13632
rect 22198 13568 22214 13632
rect 22278 13568 22294 13632
rect 22358 13568 22366 13632
rect 22046 12544 22366 13568
rect 22046 12480 22054 12544
rect 22118 12480 22134 12544
rect 22198 12480 22214 12544
rect 22278 12480 22294 12544
rect 22358 12480 22366 12544
rect 22046 11456 22366 12480
rect 22046 11392 22054 11456
rect 22118 11392 22134 11456
rect 22198 11392 22214 11456
rect 22278 11392 22294 11456
rect 22358 11392 22366 11456
rect 22046 10368 22366 11392
rect 22046 10304 22054 10368
rect 22118 10304 22134 10368
rect 22198 10304 22214 10368
rect 22278 10304 22294 10368
rect 22358 10304 22366 10368
rect 22046 9280 22366 10304
rect 22046 9216 22054 9280
rect 22118 9216 22134 9280
rect 22198 9216 22214 9280
rect 22278 9216 22294 9280
rect 22358 9216 22366 9280
rect 22046 8192 22366 9216
rect 22046 8128 22054 8192
rect 22118 8128 22134 8192
rect 22198 8128 22214 8192
rect 22278 8128 22294 8192
rect 22358 8128 22366 8192
rect 22046 7104 22366 8128
rect 22046 7040 22054 7104
rect 22118 7040 22134 7104
rect 22198 7040 22214 7104
rect 22278 7040 22294 7104
rect 22358 7040 22366 7104
rect 22046 6016 22366 7040
rect 22046 5952 22054 6016
rect 22118 5952 22134 6016
rect 22198 5952 22214 6016
rect 22278 5952 22294 6016
rect 22358 5952 22366 6016
rect 22046 4928 22366 5952
rect 22046 4864 22054 4928
rect 22118 4864 22134 4928
rect 22198 4864 22214 4928
rect 22278 4864 22294 4928
rect 22358 4864 22366 4928
rect 22046 3840 22366 4864
rect 22046 3776 22054 3840
rect 22118 3776 22134 3840
rect 22198 3776 22214 3840
rect 22278 3776 22294 3840
rect 22358 3776 22366 3840
rect 22046 2752 22366 3776
rect 22046 2688 22054 2752
rect 22118 2688 22134 2752
rect 22198 2688 22214 2752
rect 22278 2688 22294 2752
rect 22358 2688 22366 2752
rect 22046 2128 22366 2688
rect 26266 39200 26586 39760
rect 26266 39136 26274 39200
rect 26338 39136 26354 39200
rect 26418 39136 26434 39200
rect 26498 39136 26514 39200
rect 26578 39136 26586 39200
rect 26266 38112 26586 39136
rect 26266 38048 26274 38112
rect 26338 38048 26354 38112
rect 26418 38048 26434 38112
rect 26498 38048 26514 38112
rect 26578 38048 26586 38112
rect 26266 37024 26586 38048
rect 26266 36960 26274 37024
rect 26338 36960 26354 37024
rect 26418 36960 26434 37024
rect 26498 36960 26514 37024
rect 26578 36960 26586 37024
rect 26266 35936 26586 36960
rect 26266 35872 26274 35936
rect 26338 35872 26354 35936
rect 26418 35872 26434 35936
rect 26498 35872 26514 35936
rect 26578 35872 26586 35936
rect 26266 34848 26586 35872
rect 26266 34784 26274 34848
rect 26338 34784 26354 34848
rect 26418 34784 26434 34848
rect 26498 34784 26514 34848
rect 26578 34784 26586 34848
rect 26266 33760 26586 34784
rect 26266 33696 26274 33760
rect 26338 33696 26354 33760
rect 26418 33696 26434 33760
rect 26498 33696 26514 33760
rect 26578 33696 26586 33760
rect 26266 32672 26586 33696
rect 26266 32608 26274 32672
rect 26338 32608 26354 32672
rect 26418 32608 26434 32672
rect 26498 32608 26514 32672
rect 26578 32608 26586 32672
rect 26266 31584 26586 32608
rect 26266 31520 26274 31584
rect 26338 31520 26354 31584
rect 26418 31520 26434 31584
rect 26498 31520 26514 31584
rect 26578 31520 26586 31584
rect 26266 30496 26586 31520
rect 26266 30432 26274 30496
rect 26338 30432 26354 30496
rect 26418 30432 26434 30496
rect 26498 30432 26514 30496
rect 26578 30432 26586 30496
rect 26266 29408 26586 30432
rect 26266 29344 26274 29408
rect 26338 29344 26354 29408
rect 26418 29344 26434 29408
rect 26498 29344 26514 29408
rect 26578 29344 26586 29408
rect 26266 28320 26586 29344
rect 26266 28256 26274 28320
rect 26338 28256 26354 28320
rect 26418 28256 26434 28320
rect 26498 28256 26514 28320
rect 26578 28256 26586 28320
rect 26266 27232 26586 28256
rect 26266 27168 26274 27232
rect 26338 27168 26354 27232
rect 26418 27168 26434 27232
rect 26498 27168 26514 27232
rect 26578 27168 26586 27232
rect 26266 26144 26586 27168
rect 26266 26080 26274 26144
rect 26338 26080 26354 26144
rect 26418 26080 26434 26144
rect 26498 26080 26514 26144
rect 26578 26080 26586 26144
rect 26266 25056 26586 26080
rect 26266 24992 26274 25056
rect 26338 24992 26354 25056
rect 26418 24992 26434 25056
rect 26498 24992 26514 25056
rect 26578 24992 26586 25056
rect 26266 23968 26586 24992
rect 26266 23904 26274 23968
rect 26338 23904 26354 23968
rect 26418 23904 26434 23968
rect 26498 23904 26514 23968
rect 26578 23904 26586 23968
rect 26266 22880 26586 23904
rect 26266 22816 26274 22880
rect 26338 22816 26354 22880
rect 26418 22816 26434 22880
rect 26498 22816 26514 22880
rect 26578 22816 26586 22880
rect 26266 21792 26586 22816
rect 26266 21728 26274 21792
rect 26338 21728 26354 21792
rect 26418 21728 26434 21792
rect 26498 21728 26514 21792
rect 26578 21728 26586 21792
rect 26266 20704 26586 21728
rect 26266 20640 26274 20704
rect 26338 20640 26354 20704
rect 26418 20640 26434 20704
rect 26498 20640 26514 20704
rect 26578 20640 26586 20704
rect 26266 19616 26586 20640
rect 26266 19552 26274 19616
rect 26338 19552 26354 19616
rect 26418 19552 26434 19616
rect 26498 19552 26514 19616
rect 26578 19552 26586 19616
rect 26266 18528 26586 19552
rect 26266 18464 26274 18528
rect 26338 18464 26354 18528
rect 26418 18464 26434 18528
rect 26498 18464 26514 18528
rect 26578 18464 26586 18528
rect 26266 17440 26586 18464
rect 26266 17376 26274 17440
rect 26338 17376 26354 17440
rect 26418 17376 26434 17440
rect 26498 17376 26514 17440
rect 26578 17376 26586 17440
rect 26266 16352 26586 17376
rect 26266 16288 26274 16352
rect 26338 16288 26354 16352
rect 26418 16288 26434 16352
rect 26498 16288 26514 16352
rect 26578 16288 26586 16352
rect 26266 15264 26586 16288
rect 26266 15200 26274 15264
rect 26338 15200 26354 15264
rect 26418 15200 26434 15264
rect 26498 15200 26514 15264
rect 26578 15200 26586 15264
rect 26266 14176 26586 15200
rect 26266 14112 26274 14176
rect 26338 14112 26354 14176
rect 26418 14112 26434 14176
rect 26498 14112 26514 14176
rect 26578 14112 26586 14176
rect 26266 13088 26586 14112
rect 26266 13024 26274 13088
rect 26338 13024 26354 13088
rect 26418 13024 26434 13088
rect 26498 13024 26514 13088
rect 26578 13024 26586 13088
rect 26266 12000 26586 13024
rect 26266 11936 26274 12000
rect 26338 11936 26354 12000
rect 26418 11936 26434 12000
rect 26498 11936 26514 12000
rect 26578 11936 26586 12000
rect 26266 10912 26586 11936
rect 26266 10848 26274 10912
rect 26338 10848 26354 10912
rect 26418 10848 26434 10912
rect 26498 10848 26514 10912
rect 26578 10848 26586 10912
rect 26266 9824 26586 10848
rect 26266 9760 26274 9824
rect 26338 9760 26354 9824
rect 26418 9760 26434 9824
rect 26498 9760 26514 9824
rect 26578 9760 26586 9824
rect 26266 8736 26586 9760
rect 26266 8672 26274 8736
rect 26338 8672 26354 8736
rect 26418 8672 26434 8736
rect 26498 8672 26514 8736
rect 26578 8672 26586 8736
rect 26266 7648 26586 8672
rect 26266 7584 26274 7648
rect 26338 7584 26354 7648
rect 26418 7584 26434 7648
rect 26498 7584 26514 7648
rect 26578 7584 26586 7648
rect 26266 6560 26586 7584
rect 26266 6496 26274 6560
rect 26338 6496 26354 6560
rect 26418 6496 26434 6560
rect 26498 6496 26514 6560
rect 26578 6496 26586 6560
rect 26266 5472 26586 6496
rect 26266 5408 26274 5472
rect 26338 5408 26354 5472
rect 26418 5408 26434 5472
rect 26498 5408 26514 5472
rect 26578 5408 26586 5472
rect 26266 4384 26586 5408
rect 26266 4320 26274 4384
rect 26338 4320 26354 4384
rect 26418 4320 26434 4384
rect 26498 4320 26514 4384
rect 26578 4320 26586 4384
rect 26266 3296 26586 4320
rect 26266 3232 26274 3296
rect 26338 3232 26354 3296
rect 26418 3232 26434 3296
rect 26498 3232 26514 3296
rect 26578 3232 26586 3296
rect 26266 2208 26586 3232
rect 26266 2144 26274 2208
rect 26338 2144 26354 2208
rect 26418 2144 26434 2208
rect 26498 2144 26514 2208
rect 26578 2144 26586 2208
rect 26266 2128 26586 2144
rect 30487 39744 30807 39760
rect 30487 39680 30495 39744
rect 30559 39680 30575 39744
rect 30639 39680 30655 39744
rect 30719 39680 30735 39744
rect 30799 39680 30807 39744
rect 30487 38656 30807 39680
rect 30487 38592 30495 38656
rect 30559 38592 30575 38656
rect 30639 38592 30655 38656
rect 30719 38592 30735 38656
rect 30799 38592 30807 38656
rect 30487 37568 30807 38592
rect 30487 37504 30495 37568
rect 30559 37504 30575 37568
rect 30639 37504 30655 37568
rect 30719 37504 30735 37568
rect 30799 37504 30807 37568
rect 30487 36480 30807 37504
rect 30487 36416 30495 36480
rect 30559 36416 30575 36480
rect 30639 36416 30655 36480
rect 30719 36416 30735 36480
rect 30799 36416 30807 36480
rect 30487 35392 30807 36416
rect 30487 35328 30495 35392
rect 30559 35328 30575 35392
rect 30639 35328 30655 35392
rect 30719 35328 30735 35392
rect 30799 35328 30807 35392
rect 30487 34304 30807 35328
rect 30487 34240 30495 34304
rect 30559 34240 30575 34304
rect 30639 34240 30655 34304
rect 30719 34240 30735 34304
rect 30799 34240 30807 34304
rect 30487 33216 30807 34240
rect 30487 33152 30495 33216
rect 30559 33152 30575 33216
rect 30639 33152 30655 33216
rect 30719 33152 30735 33216
rect 30799 33152 30807 33216
rect 30487 32128 30807 33152
rect 30487 32064 30495 32128
rect 30559 32064 30575 32128
rect 30639 32064 30655 32128
rect 30719 32064 30735 32128
rect 30799 32064 30807 32128
rect 30487 31040 30807 32064
rect 30487 30976 30495 31040
rect 30559 30976 30575 31040
rect 30639 30976 30655 31040
rect 30719 30976 30735 31040
rect 30799 30976 30807 31040
rect 30487 29952 30807 30976
rect 30487 29888 30495 29952
rect 30559 29888 30575 29952
rect 30639 29888 30655 29952
rect 30719 29888 30735 29952
rect 30799 29888 30807 29952
rect 30487 28864 30807 29888
rect 30487 28800 30495 28864
rect 30559 28800 30575 28864
rect 30639 28800 30655 28864
rect 30719 28800 30735 28864
rect 30799 28800 30807 28864
rect 30487 27776 30807 28800
rect 30487 27712 30495 27776
rect 30559 27712 30575 27776
rect 30639 27712 30655 27776
rect 30719 27712 30735 27776
rect 30799 27712 30807 27776
rect 30487 26688 30807 27712
rect 30487 26624 30495 26688
rect 30559 26624 30575 26688
rect 30639 26624 30655 26688
rect 30719 26624 30735 26688
rect 30799 26624 30807 26688
rect 30487 25600 30807 26624
rect 30487 25536 30495 25600
rect 30559 25536 30575 25600
rect 30639 25536 30655 25600
rect 30719 25536 30735 25600
rect 30799 25536 30807 25600
rect 30487 24512 30807 25536
rect 30487 24448 30495 24512
rect 30559 24448 30575 24512
rect 30639 24448 30655 24512
rect 30719 24448 30735 24512
rect 30799 24448 30807 24512
rect 30487 23424 30807 24448
rect 30487 23360 30495 23424
rect 30559 23360 30575 23424
rect 30639 23360 30655 23424
rect 30719 23360 30735 23424
rect 30799 23360 30807 23424
rect 30487 22336 30807 23360
rect 30487 22272 30495 22336
rect 30559 22272 30575 22336
rect 30639 22272 30655 22336
rect 30719 22272 30735 22336
rect 30799 22272 30807 22336
rect 30487 21248 30807 22272
rect 30487 21184 30495 21248
rect 30559 21184 30575 21248
rect 30639 21184 30655 21248
rect 30719 21184 30735 21248
rect 30799 21184 30807 21248
rect 30487 20160 30807 21184
rect 30487 20096 30495 20160
rect 30559 20096 30575 20160
rect 30639 20096 30655 20160
rect 30719 20096 30735 20160
rect 30799 20096 30807 20160
rect 30487 19072 30807 20096
rect 30487 19008 30495 19072
rect 30559 19008 30575 19072
rect 30639 19008 30655 19072
rect 30719 19008 30735 19072
rect 30799 19008 30807 19072
rect 30487 17984 30807 19008
rect 30487 17920 30495 17984
rect 30559 17920 30575 17984
rect 30639 17920 30655 17984
rect 30719 17920 30735 17984
rect 30799 17920 30807 17984
rect 30487 16896 30807 17920
rect 30487 16832 30495 16896
rect 30559 16832 30575 16896
rect 30639 16832 30655 16896
rect 30719 16832 30735 16896
rect 30799 16832 30807 16896
rect 30487 15808 30807 16832
rect 30487 15744 30495 15808
rect 30559 15744 30575 15808
rect 30639 15744 30655 15808
rect 30719 15744 30735 15808
rect 30799 15744 30807 15808
rect 30487 14720 30807 15744
rect 30487 14656 30495 14720
rect 30559 14656 30575 14720
rect 30639 14656 30655 14720
rect 30719 14656 30735 14720
rect 30799 14656 30807 14720
rect 30487 13632 30807 14656
rect 30487 13568 30495 13632
rect 30559 13568 30575 13632
rect 30639 13568 30655 13632
rect 30719 13568 30735 13632
rect 30799 13568 30807 13632
rect 30487 12544 30807 13568
rect 30487 12480 30495 12544
rect 30559 12480 30575 12544
rect 30639 12480 30655 12544
rect 30719 12480 30735 12544
rect 30799 12480 30807 12544
rect 30487 11456 30807 12480
rect 30487 11392 30495 11456
rect 30559 11392 30575 11456
rect 30639 11392 30655 11456
rect 30719 11392 30735 11456
rect 30799 11392 30807 11456
rect 30487 10368 30807 11392
rect 30487 10304 30495 10368
rect 30559 10304 30575 10368
rect 30639 10304 30655 10368
rect 30719 10304 30735 10368
rect 30799 10304 30807 10368
rect 30487 9280 30807 10304
rect 30487 9216 30495 9280
rect 30559 9216 30575 9280
rect 30639 9216 30655 9280
rect 30719 9216 30735 9280
rect 30799 9216 30807 9280
rect 30487 8192 30807 9216
rect 30487 8128 30495 8192
rect 30559 8128 30575 8192
rect 30639 8128 30655 8192
rect 30719 8128 30735 8192
rect 30799 8128 30807 8192
rect 30487 7104 30807 8128
rect 30487 7040 30495 7104
rect 30559 7040 30575 7104
rect 30639 7040 30655 7104
rect 30719 7040 30735 7104
rect 30799 7040 30807 7104
rect 30487 6016 30807 7040
rect 30487 5952 30495 6016
rect 30559 5952 30575 6016
rect 30639 5952 30655 6016
rect 30719 5952 30735 6016
rect 30799 5952 30807 6016
rect 30487 4928 30807 5952
rect 30487 4864 30495 4928
rect 30559 4864 30575 4928
rect 30639 4864 30655 4928
rect 30719 4864 30735 4928
rect 30799 4864 30807 4928
rect 30487 3840 30807 4864
rect 30487 3776 30495 3840
rect 30559 3776 30575 3840
rect 30639 3776 30655 3840
rect 30719 3776 30735 3840
rect 30799 3776 30807 3840
rect 30487 2752 30807 3776
rect 30487 2688 30495 2752
rect 30559 2688 30575 2752
rect 30639 2688 30655 2752
rect 30719 2688 30735 2752
rect 30799 2688 30807 2752
rect 30487 2128 30807 2688
rect 34707 39200 35027 39760
rect 34707 39136 34715 39200
rect 34779 39136 34795 39200
rect 34859 39136 34875 39200
rect 34939 39136 34955 39200
rect 35019 39136 35027 39200
rect 34707 38112 35027 39136
rect 34707 38048 34715 38112
rect 34779 38048 34795 38112
rect 34859 38048 34875 38112
rect 34939 38048 34955 38112
rect 35019 38048 35027 38112
rect 34707 37024 35027 38048
rect 34707 36960 34715 37024
rect 34779 36960 34795 37024
rect 34859 36960 34875 37024
rect 34939 36960 34955 37024
rect 35019 36960 35027 37024
rect 34707 35936 35027 36960
rect 34707 35872 34715 35936
rect 34779 35872 34795 35936
rect 34859 35872 34875 35936
rect 34939 35872 34955 35936
rect 35019 35872 35027 35936
rect 34707 34848 35027 35872
rect 34707 34784 34715 34848
rect 34779 34784 34795 34848
rect 34859 34784 34875 34848
rect 34939 34784 34955 34848
rect 35019 34784 35027 34848
rect 34707 33760 35027 34784
rect 34707 33696 34715 33760
rect 34779 33696 34795 33760
rect 34859 33696 34875 33760
rect 34939 33696 34955 33760
rect 35019 33696 35027 33760
rect 34707 32672 35027 33696
rect 34707 32608 34715 32672
rect 34779 32608 34795 32672
rect 34859 32608 34875 32672
rect 34939 32608 34955 32672
rect 35019 32608 35027 32672
rect 34707 31584 35027 32608
rect 34707 31520 34715 31584
rect 34779 31520 34795 31584
rect 34859 31520 34875 31584
rect 34939 31520 34955 31584
rect 35019 31520 35027 31584
rect 34707 30496 35027 31520
rect 34707 30432 34715 30496
rect 34779 30432 34795 30496
rect 34859 30432 34875 30496
rect 34939 30432 34955 30496
rect 35019 30432 35027 30496
rect 34707 29408 35027 30432
rect 34707 29344 34715 29408
rect 34779 29344 34795 29408
rect 34859 29344 34875 29408
rect 34939 29344 34955 29408
rect 35019 29344 35027 29408
rect 34707 28320 35027 29344
rect 34707 28256 34715 28320
rect 34779 28256 34795 28320
rect 34859 28256 34875 28320
rect 34939 28256 34955 28320
rect 35019 28256 35027 28320
rect 34707 27232 35027 28256
rect 34707 27168 34715 27232
rect 34779 27168 34795 27232
rect 34859 27168 34875 27232
rect 34939 27168 34955 27232
rect 35019 27168 35027 27232
rect 34707 26144 35027 27168
rect 34707 26080 34715 26144
rect 34779 26080 34795 26144
rect 34859 26080 34875 26144
rect 34939 26080 34955 26144
rect 35019 26080 35027 26144
rect 34707 25056 35027 26080
rect 34707 24992 34715 25056
rect 34779 24992 34795 25056
rect 34859 24992 34875 25056
rect 34939 24992 34955 25056
rect 35019 24992 35027 25056
rect 34707 23968 35027 24992
rect 34707 23904 34715 23968
rect 34779 23904 34795 23968
rect 34859 23904 34875 23968
rect 34939 23904 34955 23968
rect 35019 23904 35027 23968
rect 34707 22880 35027 23904
rect 34707 22816 34715 22880
rect 34779 22816 34795 22880
rect 34859 22816 34875 22880
rect 34939 22816 34955 22880
rect 35019 22816 35027 22880
rect 34707 21792 35027 22816
rect 34707 21728 34715 21792
rect 34779 21728 34795 21792
rect 34859 21728 34875 21792
rect 34939 21728 34955 21792
rect 35019 21728 35027 21792
rect 34707 20704 35027 21728
rect 34707 20640 34715 20704
rect 34779 20640 34795 20704
rect 34859 20640 34875 20704
rect 34939 20640 34955 20704
rect 35019 20640 35027 20704
rect 34707 19616 35027 20640
rect 34707 19552 34715 19616
rect 34779 19552 34795 19616
rect 34859 19552 34875 19616
rect 34939 19552 34955 19616
rect 35019 19552 35027 19616
rect 34707 18528 35027 19552
rect 34707 18464 34715 18528
rect 34779 18464 34795 18528
rect 34859 18464 34875 18528
rect 34939 18464 34955 18528
rect 35019 18464 35027 18528
rect 34707 17440 35027 18464
rect 34707 17376 34715 17440
rect 34779 17376 34795 17440
rect 34859 17376 34875 17440
rect 34939 17376 34955 17440
rect 35019 17376 35027 17440
rect 34707 16352 35027 17376
rect 34707 16288 34715 16352
rect 34779 16288 34795 16352
rect 34859 16288 34875 16352
rect 34939 16288 34955 16352
rect 35019 16288 35027 16352
rect 34707 15264 35027 16288
rect 34707 15200 34715 15264
rect 34779 15200 34795 15264
rect 34859 15200 34875 15264
rect 34939 15200 34955 15264
rect 35019 15200 35027 15264
rect 34707 14176 35027 15200
rect 34707 14112 34715 14176
rect 34779 14112 34795 14176
rect 34859 14112 34875 14176
rect 34939 14112 34955 14176
rect 35019 14112 35027 14176
rect 34707 13088 35027 14112
rect 34707 13024 34715 13088
rect 34779 13024 34795 13088
rect 34859 13024 34875 13088
rect 34939 13024 34955 13088
rect 35019 13024 35027 13088
rect 34707 12000 35027 13024
rect 34707 11936 34715 12000
rect 34779 11936 34795 12000
rect 34859 11936 34875 12000
rect 34939 11936 34955 12000
rect 35019 11936 35027 12000
rect 34707 10912 35027 11936
rect 34707 10848 34715 10912
rect 34779 10848 34795 10912
rect 34859 10848 34875 10912
rect 34939 10848 34955 10912
rect 35019 10848 35027 10912
rect 34707 9824 35027 10848
rect 34707 9760 34715 9824
rect 34779 9760 34795 9824
rect 34859 9760 34875 9824
rect 34939 9760 34955 9824
rect 35019 9760 35027 9824
rect 34707 8736 35027 9760
rect 34707 8672 34715 8736
rect 34779 8672 34795 8736
rect 34859 8672 34875 8736
rect 34939 8672 34955 8736
rect 35019 8672 35027 8736
rect 34707 7648 35027 8672
rect 34707 7584 34715 7648
rect 34779 7584 34795 7648
rect 34859 7584 34875 7648
rect 34939 7584 34955 7648
rect 35019 7584 35027 7648
rect 34707 6560 35027 7584
rect 34707 6496 34715 6560
rect 34779 6496 34795 6560
rect 34859 6496 34875 6560
rect 34939 6496 34955 6560
rect 35019 6496 35027 6560
rect 34707 5472 35027 6496
rect 34707 5408 34715 5472
rect 34779 5408 34795 5472
rect 34859 5408 34875 5472
rect 34939 5408 34955 5472
rect 35019 5408 35027 5472
rect 34707 4384 35027 5408
rect 34707 4320 34715 4384
rect 34779 4320 34795 4384
rect 34859 4320 34875 4384
rect 34939 4320 34955 4384
rect 35019 4320 35027 4384
rect 34707 3296 35027 4320
rect 34707 3232 34715 3296
rect 34779 3232 34795 3296
rect 34859 3232 34875 3296
rect 34939 3232 34955 3296
rect 35019 3232 35027 3296
rect 34707 2208 35027 3232
rect 34707 2144 34715 2208
rect 34779 2144 34795 2208
rect 34859 2144 34875 2208
rect 34939 2144 34955 2208
rect 35019 2144 35027 2208
rect 34707 2128 35027 2144
use sky130_fd_sc_hd__inv_2  _427_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 25392 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _428_
timestamp 1688980957
transform 1 0 24840 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _429_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 24840 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _430_
timestamp 1688980957
transform 1 0 24748 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _431_
timestamp 1688980957
transform 1 0 24656 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _432_
timestamp 1688980957
transform 1 0 25024 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _433_
timestamp 1688980957
transform 1 0 24840 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _434_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 24748 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _435_
timestamp 1688980957
transform 1 0 26312 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _436_
timestamp 1688980957
transform -1 0 26312 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _437_
timestamp 1688980957
transform 1 0 24840 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _438_
timestamp 1688980957
transform -1 0 25852 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _439_
timestamp 1688980957
transform 1 0 25300 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _440_
timestamp 1688980957
transform -1 0 25852 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _441_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 25116 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _442_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 25852 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _443_
timestamp 1688980957
transform 1 0 25116 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  _444_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 17664 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _445_
timestamp 1688980957
transform 1 0 24472 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _446_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 26036 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _447_
timestamp 1688980957
transform -1 0 26312 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _448_
timestamp 1688980957
transform 1 0 25484 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _449_
timestamp 1688980957
transform -1 0 20516 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _450_
timestamp 1688980957
transform -1 0 20240 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _451_
timestamp 1688980957
transform -1 0 19504 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _452_
timestamp 1688980957
transform -1 0 19136 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _453_
timestamp 1688980957
transform -1 0 20148 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _454_
timestamp 1688980957
transform -1 0 19688 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _455_
timestamp 1688980957
transform -1 0 20424 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _456_
timestamp 1688980957
transform -1 0 20332 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _457_
timestamp 1688980957
transform -1 0 20608 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _458_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 19136 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _459_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 19136 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _460_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 20332 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _461_
timestamp 1688980957
transform -1 0 20148 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _462_
timestamp 1688980957
transform -1 0 19320 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _463_
timestamp 1688980957
transform 1 0 19228 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _464_
timestamp 1688980957
transform -1 0 19228 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _465_
timestamp 1688980957
transform 1 0 18584 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  _466_
timestamp 1688980957
transform 1 0 21620 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__a211oi_1  _467_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 19228 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _468_
timestamp 1688980957
transform -1 0 20148 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _469_
timestamp 1688980957
transform -1 0 19688 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _470_
timestamp 1688980957
transform -1 0 19320 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _471_
timestamp 1688980957
transform -1 0 19228 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _472_
timestamp 1688980957
transform -1 0 19136 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _473_
timestamp 1688980957
transform 1 0 18216 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _474_
timestamp 1688980957
transform -1 0 19504 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _475_
timestamp 1688980957
transform -1 0 19136 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _476_
timestamp 1688980957
transform -1 0 19964 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _477_
timestamp 1688980957
transform 1 0 18676 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _478_
timestamp 1688980957
transform -1 0 18676 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _479_
timestamp 1688980957
transform 1 0 18032 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _480_
timestamp 1688980957
transform 1 0 17572 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _481_
timestamp 1688980957
transform 1 0 18216 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _482_
timestamp 1688980957
transform -1 0 18952 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _483_
timestamp 1688980957
transform 1 0 18308 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _484_
timestamp 1688980957
transform 1 0 19228 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__a211oi_2  _485_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 18216 0 1 30464
box -38 -48 958 592
use sky130_fd_sc_hd__inv_2  _486_
timestamp 1688980957
transform 1 0 16100 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _487_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 29808 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__o41a_1  _488_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 30084 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__and4_1  _489_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 29716 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__a41o_1  _490_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 30912 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  _491_
timestamp 1688980957
transform 1 0 29440 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _492_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 29808 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  _493_
timestamp 1688980957
transform 1 0 25300 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _494_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 22908 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _495_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 23828 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _496_
timestamp 1688980957
transform 1 0 28704 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _497_
timestamp 1688980957
transform 1 0 29164 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _498_
timestamp 1688980957
transform 1 0 28704 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _499_
timestamp 1688980957
transform 1 0 29532 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _500_
timestamp 1688980957
transform 1 0 30360 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _501_
timestamp 1688980957
transform 1 0 31280 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _502_
timestamp 1688980957
transform 1 0 29808 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _503_
timestamp 1688980957
transform 1 0 30728 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _504_
timestamp 1688980957
transform 1 0 30820 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _505_
timestamp 1688980957
transform -1 0 30728 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _506_
timestamp 1688980957
transform 1 0 29716 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _507_
timestamp 1688980957
transform 1 0 30544 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _508_
timestamp 1688980957
transform -1 0 31464 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _509_
timestamp 1688980957
transform 1 0 31372 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _510_
timestamp 1688980957
transform -1 0 32752 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _511_
timestamp 1688980957
transform 1 0 31464 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__o41a_1  _512_
timestamp 1688980957
transform 1 0 32108 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__and4_1  _513_
timestamp 1688980957
transform 1 0 32108 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a41o_1  _514_
timestamp 1688980957
transform 1 0 32108 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _515_
timestamp 1688980957
transform -1 0 31832 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _516_
timestamp 1688980957
transform -1 0 32292 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _517_
timestamp 1688980957
transform 1 0 31648 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _518_
timestamp 1688980957
transform -1 0 32568 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _519_
timestamp 1688980957
transform -1 0 31832 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _520_
timestamp 1688980957
transform -1 0 31096 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _521_
timestamp 1688980957
transform 1 0 30360 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _522_
timestamp 1688980957
transform 1 0 30820 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _523_
timestamp 1688980957
transform -1 0 31372 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _524_
timestamp 1688980957
transform 1 0 31556 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _525_
timestamp 1688980957
transform 1 0 32292 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _526_
timestamp 1688980957
transform -1 0 31464 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _527_
timestamp 1688980957
transform 1 0 30728 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _528_
timestamp 1688980957
transform 1 0 30636 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _529_
timestamp 1688980957
transform 1 0 31280 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _530_
timestamp 1688980957
transform 1 0 26496 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _531_
timestamp 1688980957
transform 1 0 32108 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _532_
timestamp 1688980957
transform 1 0 32568 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _533_
timestamp 1688980957
transform 1 0 32108 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__o41a_1  _534_
timestamp 1688980957
transform 1 0 32108 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__and4_1  _535_
timestamp 1688980957
transform 1 0 32476 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a41o_1  _536_
timestamp 1688980957
transform 1 0 32936 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _537_
timestamp 1688980957
transform 1 0 30728 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _538_
timestamp 1688980957
transform 1 0 31280 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _539_
timestamp 1688980957
transform 1 0 31464 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _540_
timestamp 1688980957
transform 1 0 30912 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _541_
timestamp 1688980957
transform 1 0 31372 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _542_
timestamp 1688980957
transform -1 0 31648 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _543_
timestamp 1688980957
transform -1 0 30544 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _544_
timestamp 1688980957
transform 1 0 32200 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _545_
timestamp 1688980957
transform 1 0 33028 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _546_
timestamp 1688980957
transform 1 0 33120 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _547_
timestamp 1688980957
transform 1 0 33304 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _548_
timestamp 1688980957
transform -1 0 30452 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _549_
timestamp 1688980957
transform -1 0 30176 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _550_
timestamp 1688980957
transform 1 0 30268 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _551_
timestamp 1688980957
transform 1 0 31004 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _552_
timestamp 1688980957
transform 1 0 31648 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _553_
timestamp 1688980957
transform 1 0 33580 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _554_
timestamp 1688980957
transform -1 0 27876 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__o41a_1  _555_
timestamp 1688980957
transform 1 0 27140 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__and4_1  _556_
timestamp 1688980957
transform 1 0 27232 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a41o_1  _557_
timestamp 1688980957
transform 1 0 27232 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _558_
timestamp 1688980957
transform -1 0 27140 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _559_
timestamp 1688980957
transform 1 0 23000 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _560_
timestamp 1688980957
transform -1 0 24380 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _561_
timestamp 1688980957
transform 1 0 26128 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _562_
timestamp 1688980957
transform 1 0 26312 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _563_
timestamp 1688980957
transform -1 0 27416 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _564_
timestamp 1688980957
transform -1 0 26864 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _565_
timestamp 1688980957
transform -1 0 25668 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _566_
timestamp 1688980957
transform 1 0 27876 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _567_
timestamp 1688980957
transform -1 0 29072 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _568_
timestamp 1688980957
transform -1 0 28796 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _569_
timestamp 1688980957
transform -1 0 28428 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _570_
timestamp 1688980957
transform 1 0 25944 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _571_
timestamp 1688980957
transform 1 0 26404 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _572_
timestamp 1688980957
transform 1 0 26956 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _573_
timestamp 1688980957
transform 1 0 26956 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _574_
timestamp 1688980957
transform 1 0 27968 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _575_
timestamp 1688980957
transform -1 0 28796 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _576_
timestamp 1688980957
transform 1 0 25944 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__o41a_1  _577_
timestamp 1688980957
transform 1 0 25852 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__and4_1  _578_
timestamp 1688980957
transform 1 0 25576 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a41o_1  _579_
timestamp 1688980957
transform 1 0 25852 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _580_
timestamp 1688980957
transform 1 0 25484 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _581_
timestamp 1688980957
transform 1 0 22448 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _582_
timestamp 1688980957
transform -1 0 23460 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _583_
timestamp 1688980957
transform -1 0 24932 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _584_
timestamp 1688980957
transform -1 0 24656 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _585_
timestamp 1688980957
transform -1 0 25392 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _586_
timestamp 1688980957
transform -1 0 24288 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _587_
timestamp 1688980957
transform 1 0 25760 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _588_
timestamp 1688980957
transform -1 0 26772 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _589_
timestamp 1688980957
transform 1 0 26404 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _590_
timestamp 1688980957
transform -1 0 26864 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _591_
timestamp 1688980957
transform -1 0 25484 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _592_
timestamp 1688980957
transform 1 0 24748 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _593_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 26128 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _594_
timestamp 1688980957
transform -1 0 26680 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _595_
timestamp 1688980957
transform -1 0 25852 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _596_
timestamp 1688980957
transform -1 0 27416 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _597_
timestamp 1688980957
transform -1 0 27232 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _598_
timestamp 1688980957
transform -1 0 29440 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__o41a_1  _599_
timestamp 1688980957
transform 1 0 29532 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__and4_1  _600_
timestamp 1688980957
transform 1 0 29532 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a41o_1  _601_
timestamp 1688980957
transform 1 0 29256 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _602_
timestamp 1688980957
transform -1 0 29440 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _603_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 16836 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _604_
timestamp 1688980957
transform 1 0 25208 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _605_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 18492 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _606_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 17572 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _607_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 17940 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _608_
timestamp 1688980957
transform -1 0 17480 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_1  _609_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 17204 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _610_
timestamp 1688980957
transform -1 0 17848 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _611_
timestamp 1688980957
transform 1 0 18032 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _612_
timestamp 1688980957
transform -1 0 18124 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _613_
timestamp 1688980957
transform 1 0 24840 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _614_
timestamp 1688980957
transform -1 0 18216 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _615_
timestamp 1688980957
transform 1 0 17020 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _616_
timestamp 1688980957
transform 1 0 16836 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _617_
timestamp 1688980957
transform -1 0 17664 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _618_
timestamp 1688980957
transform -1 0 16560 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _619_
timestamp 1688980957
transform 1 0 16652 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _620_
timestamp 1688980957
transform 1 0 17388 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _621_
timestamp 1688980957
transform 1 0 17848 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _622_
timestamp 1688980957
transform 1 0 16744 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _623_
timestamp 1688980957
transform -1 0 18492 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _624_
timestamp 1688980957
transform 1 0 17388 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _625_
timestamp 1688980957
transform 1 0 29440 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _626_
timestamp 1688980957
transform 1 0 29900 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _627_
timestamp 1688980957
transform 1 0 27876 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _628_
timestamp 1688980957
transform 1 0 27968 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _629_
timestamp 1688980957
transform -1 0 28796 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _630_
timestamp 1688980957
transform -1 0 28520 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _631_
timestamp 1688980957
transform 1 0 28796 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _632_
timestamp 1688980957
transform -1 0 29808 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _633_
timestamp 1688980957
transform -1 0 31832 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _634_
timestamp 1688980957
transform -1 0 30084 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _635_
timestamp 1688980957
transform 1 0 30176 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _636_
timestamp 1688980957
transform -1 0 30912 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _637_
timestamp 1688980957
transform -1 0 28244 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _638_
timestamp 1688980957
transform 1 0 27508 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _639_
timestamp 1688980957
transform -1 0 29256 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _640_
timestamp 1688980957
transform -1 0 28520 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _641_
timestamp 1688980957
transform -1 0 30820 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _642_
timestamp 1688980957
transform -1 0 29900 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _643_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 29532 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _644_
timestamp 1688980957
transform 1 0 29532 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _645_
timestamp 1688980957
transform 1 0 30084 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _646_
timestamp 1688980957
transform -1 0 29440 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_2  _647_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 29256 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _648_
timestamp 1688980957
transform 1 0 28796 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _649_
timestamp 1688980957
transform 1 0 25944 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _650_
timestamp 1688980957
transform 1 0 25852 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _651_
timestamp 1688980957
transform 1 0 29992 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _652_
timestamp 1688980957
transform -1 0 28336 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _653_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 28888 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _654_
timestamp 1688980957
transform 1 0 26496 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _655_
timestamp 1688980957
transform -1 0 28612 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _656_
timestamp 1688980957
transform 1 0 26956 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _657_
timestamp 1688980957
transform -1 0 27876 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__a21boi_2  _658_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 27324 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _659_
timestamp 1688980957
transform 1 0 28704 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _660_
timestamp 1688980957
transform -1 0 28520 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _661_
timestamp 1688980957
transform 1 0 28888 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _662_
timestamp 1688980957
transform -1 0 29440 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _663_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 28244 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _664_
timestamp 1688980957
transform -1 0 29440 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _665_
timestamp 1688980957
transform -1 0 29440 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _666_
timestamp 1688980957
transform 1 0 26956 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _667_
timestamp 1688980957
transform 1 0 27784 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _668_
timestamp 1688980957
transform -1 0 27968 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _669_
timestamp 1688980957
transform 1 0 27048 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _670_
timestamp 1688980957
transform 1 0 25944 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _671_
timestamp 1688980957
transform 1 0 27232 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_1  _672_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 28244 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _673_
timestamp 1688980957
transform -1 0 28520 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _674_
timestamp 1688980957
transform -1 0 28980 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _675_
timestamp 1688980957
transform -1 0 28152 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _676_
timestamp 1688980957
transform -1 0 28612 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _677_
timestamp 1688980957
transform -1 0 28980 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _678_
timestamp 1688980957
transform 1 0 26404 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _679_
timestamp 1688980957
transform -1 0 28244 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _680_
timestamp 1688980957
transform 1 0 28612 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _681_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 27692 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _682_
timestamp 1688980957
transform 1 0 25944 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _683_
timestamp 1688980957
transform -1 0 26864 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _684_
timestamp 1688980957
transform -1 0 26588 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _685_
timestamp 1688980957
transform -1 0 27416 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _686_
timestamp 1688980957
transform 1 0 26956 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _687_
timestamp 1688980957
transform 1 0 27416 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_1  _688_
timestamp 1688980957
transform 1 0 27232 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _689_
timestamp 1688980957
transform 1 0 27416 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _690_
timestamp 1688980957
transform -1 0 27140 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__o22ai_1  _691_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 25944 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _692_
timestamp 1688980957
transform 1 0 23828 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _693_
timestamp 1688980957
transform -1 0 24196 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _694_
timestamp 1688980957
transform 1 0 25668 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _695_
timestamp 1688980957
transform 1 0 25852 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__o31ai_1  _696_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 26864 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _697_
timestamp 1688980957
transform 1 0 25760 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _698_
timestamp 1688980957
transform 1 0 24748 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _699_
timestamp 1688980957
transform -1 0 25944 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _700_
timestamp 1688980957
transform 1 0 28152 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _701_
timestamp 1688980957
transform 1 0 29072 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _702_
timestamp 1688980957
transform -1 0 25668 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _703_
timestamp 1688980957
transform -1 0 25116 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _704_
timestamp 1688980957
transform -1 0 25576 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _705_
timestamp 1688980957
transform 1 0 25944 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_2  _706_
timestamp 1688980957
transform 1 0 24380 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _707_
timestamp 1688980957
transform 1 0 20884 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _708_
timestamp 1688980957
transform 1 0 20884 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _709_
timestamp 1688980957
transform 1 0 20332 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _710_
timestamp 1688980957
transform 1 0 23644 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _711_
timestamp 1688980957
transform -1 0 23092 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _712_
timestamp 1688980957
transform -1 0 22080 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _713_
timestamp 1688980957
transform 1 0 21344 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _714_
timestamp 1688980957
transform 1 0 21252 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _715_
timestamp 1688980957
transform 1 0 21344 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _716_
timestamp 1688980957
transform 1 0 21804 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__a21boi_2  _717_
timestamp 1688980957
transform 1 0 21804 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _718_
timestamp 1688980957
transform 1 0 22356 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _719_
timestamp 1688980957
transform -1 0 23000 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _720_
timestamp 1688980957
transform -1 0 23092 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _721_
timestamp 1688980957
transform 1 0 22540 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _722_
timestamp 1688980957
transform 1 0 21896 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _723_
timestamp 1688980957
transform 1 0 23828 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _724_
timestamp 1688980957
transform 1 0 23092 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _725_
timestamp 1688980957
transform 1 0 21068 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _726_
timestamp 1688980957
transform -1 0 21896 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _727_
timestamp 1688980957
transform -1 0 21896 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _728_
timestamp 1688980957
transform 1 0 20976 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _729_
timestamp 1688980957
transform 1 0 20148 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _730_
timestamp 1688980957
transform 1 0 21160 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_1  _731_
timestamp 1688980957
transform -1 0 22448 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _732_
timestamp 1688980957
transform -1 0 22264 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _733_
timestamp 1688980957
transform -1 0 23828 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _734_
timestamp 1688980957
transform -1 0 22724 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _735_
timestamp 1688980957
transform 1 0 23276 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _736_
timestamp 1688980957
transform -1 0 22816 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _737_
timestamp 1688980957
transform 1 0 23736 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _738_
timestamp 1688980957
transform -1 0 23920 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _739_
timestamp 1688980957
transform 1 0 21804 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _740_
timestamp 1688980957
transform 1 0 22724 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__o31ai_1  _741_
timestamp 1688980957
transform -1 0 23368 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _742_
timestamp 1688980957
transform 1 0 22724 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _743_
timestamp 1688980957
transform -1 0 21620 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _744_
timestamp 1688980957
transform -1 0 21344 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _745_
timestamp 1688980957
transform 1 0 21344 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _746_
timestamp 1688980957
transform -1 0 22816 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_1  _747_
timestamp 1688980957
transform 1 0 21988 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _748_
timestamp 1688980957
transform -1 0 21896 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _749_
timestamp 1688980957
transform -1 0 21712 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _750_
timestamp 1688980957
transform 1 0 19504 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _751_
timestamp 1688980957
transform 1 0 19780 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _752_
timestamp 1688980957
transform 1 0 20240 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _753_
timestamp 1688980957
transform 1 0 20792 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__o31ai_1  _754_
timestamp 1688980957
transform -1 0 20792 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _755_
timestamp 1688980957
transform -1 0 20976 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _756_
timestamp 1688980957
transform 1 0 23736 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _757_
timestamp 1688980957
transform 1 0 24380 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _758_
timestamp 1688980957
transform 1 0 23644 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _759_
timestamp 1688980957
transform 1 0 24380 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _760_
timestamp 1688980957
transform -1 0 24104 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _761_
timestamp 1688980957
transform -1 0 23552 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _762_
timestamp 1688980957
transform -1 0 23092 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _763_
timestamp 1688980957
transform -1 0 22264 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_2  _764_
timestamp 1688980957
transform 1 0 22264 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _765_
timestamp 1688980957
transform 1 0 21804 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _766_
timestamp 1688980957
transform 1 0 19320 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _767_
timestamp 1688980957
transform 1 0 19228 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _768_
timestamp 1688980957
transform 1 0 23000 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _769_
timestamp 1688980957
transform -1 0 21160 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _770_
timestamp 1688980957
transform -1 0 20240 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _771_
timestamp 1688980957
transform -1 0 20700 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _772_
timestamp 1688980957
transform -1 0 21528 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _773_
timestamp 1688980957
transform 1 0 20884 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _774_
timestamp 1688980957
transform 1 0 20148 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__a21boi_2  _775_
timestamp 1688980957
transform 1 0 20240 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _776_
timestamp 1688980957
transform -1 0 21528 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _777_
timestamp 1688980957
transform -1 0 20424 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _778_
timestamp 1688980957
transform -1 0 21436 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _779_
timestamp 1688980957
transform -1 0 21344 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _780_
timestamp 1688980957
transform 1 0 20424 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _781_
timestamp 1688980957
transform -1 0 22356 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _782_
timestamp 1688980957
transform -1 0 22080 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _783_
timestamp 1688980957
transform 1 0 19136 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _784_
timestamp 1688980957
transform 1 0 20792 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _785_
timestamp 1688980957
transform 1 0 20700 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _786_
timestamp 1688980957
transform 1 0 20148 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _787_
timestamp 1688980957
transform 1 0 19412 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _788_
timestamp 1688980957
transform 1 0 19780 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_1  _789_
timestamp 1688980957
transform -1 0 20792 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _790_
timestamp 1688980957
transform -1 0 19872 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _791_
timestamp 1688980957
transform 1 0 19872 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _792_
timestamp 1688980957
transform 1 0 20240 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _793_
timestamp 1688980957
transform 1 0 20884 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _794_
timestamp 1688980957
transform 1 0 21804 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _795_
timestamp 1688980957
transform 1 0 21344 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _796_
timestamp 1688980957
transform -1 0 21252 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _797_
timestamp 1688980957
transform 1 0 19228 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _798_
timestamp 1688980957
transform -1 0 21252 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__o31ai_1  _799_
timestamp 1688980957
transform 1 0 20332 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _800_
timestamp 1688980957
transform 1 0 20700 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _801_
timestamp 1688980957
transform 1 0 21804 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _802_
timestamp 1688980957
transform 1 0 20056 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _803_
timestamp 1688980957
transform 1 0 21068 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _804_
timestamp 1688980957
transform -1 0 21620 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_1  _805_
timestamp 1688980957
transform 1 0 20056 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _806_
timestamp 1688980957
transform 1 0 20148 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _807_
timestamp 1688980957
transform -1 0 20424 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _808_
timestamp 1688980957
transform 1 0 19228 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _809_
timestamp 1688980957
transform -1 0 19044 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _810_
timestamp 1688980957
transform 1 0 20424 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _811_
timestamp 1688980957
transform -1 0 21252 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__o31ai_1  _812_
timestamp 1688980957
transform 1 0 20424 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _813_
timestamp 1688980957
transform 1 0 20976 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _814_
timestamp 1688980957
transform -1 0 23736 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _815_
timestamp 1688980957
transform 1 0 22264 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _816_
timestamp 1688980957
transform -1 0 22908 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _817_
timestamp 1688980957
transform -1 0 25944 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _818_
timestamp 1688980957
transform 1 0 24656 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _819_
timestamp 1688980957
transform -1 0 24840 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _820_
timestamp 1688980957
transform -1 0 24012 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_1  _821_
timestamp 1688980957
transform -1 0 22816 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _822_
timestamp 1688980957
transform -1 0 24012 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _823_
timestamp 1688980957
transform -1 0 24748 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _824_
timestamp 1688980957
transform -1 0 24288 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _825_
timestamp 1688980957
transform -1 0 24104 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _826_
timestamp 1688980957
transform -1 0 23276 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _827_
timestamp 1688980957
transform 1 0 22908 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _828_
timestamp 1688980957
transform -1 0 23920 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _829_
timestamp 1688980957
transform -1 0 23184 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _830_
timestamp 1688980957
transform 1 0 22632 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _831_
timestamp 1688980957
transform 1 0 23828 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _832_
timestamp 1688980957
transform -1 0 24196 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _833_
timestamp 1688980957
transform 1 0 23276 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _834_
timestamp 1688980957
transform -1 0 24748 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _835_
timestamp 1688980957
transform 1 0 24840 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _836_
timestamp 1688980957
transform -1 0 17572 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _837_
timestamp 1688980957
transform 1 0 18584 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _838_
timestamp 1688980957
transform -1 0 19320 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _839_
timestamp 1688980957
transform -1 0 18584 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _840_
timestamp 1688980957
transform 1 0 18584 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_1  _841_
timestamp 1688980957
transform -1 0 17756 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _842_
timestamp 1688980957
transform -1 0 17940 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _843_
timestamp 1688980957
transform 1 0 17848 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _844_
timestamp 1688980957
transform -1 0 17480 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _845_
timestamp 1688980957
transform -1 0 18768 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _846_
timestamp 1688980957
transform -1 0 17480 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _847_
timestamp 1688980957
transform 1 0 17756 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _848_
timestamp 1688980957
transform -1 0 17756 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _849_
timestamp 1688980957
transform -1 0 17296 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _850_
timestamp 1688980957
transform 1 0 17572 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _851_
timestamp 1688980957
transform 1 0 17756 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _852_
timestamp 1688980957
transform 1 0 18216 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _853_
timestamp 1688980957
transform 1 0 17112 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _854_
timestamp 1688980957
transform 1 0 18124 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _855_
timestamp 1688980957
transform 1 0 17848 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__dfstp_1  _856_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 15180 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _856__27 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 15824 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _857_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 29532 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _858_
timestamp 1688980957
transform 1 0 27232 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _859_
timestamp 1688980957
transform -1 0 29440 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _860_
timestamp 1688980957
transform 1 0 28336 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _861_
timestamp 1688980957
transform -1 0 31280 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _862_
timestamp 1688980957
transform 1 0 30452 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _863_
timestamp 1688980957
transform 1 0 29532 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _864_
timestamp 1688980957
transform 1 0 31004 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _865_
timestamp 1688980957
transform -1 0 33580 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _866_
timestamp 1688980957
transform 1 0 31648 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _867_
timestamp 1688980957
transform 1 0 31280 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _868_
timestamp 1688980957
transform 1 0 31556 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _869_
timestamp 1688980957
transform 1 0 29992 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _870_
timestamp 1688980957
transform 1 0 31004 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _871_
timestamp 1688980957
transform 1 0 31924 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _872_
timestamp 1688980957
transform 1 0 30176 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _873_
timestamp 1688980957
transform 1 0 30544 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _874_
timestamp 1688980957
transform 1 0 31924 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _875_
timestamp 1688980957
transform 1 0 30544 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _876_
timestamp 1688980957
transform 1 0 30728 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _877_
timestamp 1688980957
transform 1 0 31004 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _878_
timestamp 1688980957
transform 1 0 30544 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _879_
timestamp 1688980957
transform 1 0 32292 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _880_
timestamp 1688980957
transform 1 0 32476 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _881_
timestamp 1688980957
transform 1 0 29900 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _882_
timestamp 1688980957
transform 1 0 30452 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _883_
timestamp 1688980957
transform 1 0 32108 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _884_
timestamp 1688980957
transform -1 0 28428 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _885_
timestamp 1688980957
transform 1 0 24656 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _886_
timestamp 1688980957
transform 1 0 25852 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _887_
timestamp 1688980957
transform 1 0 26956 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _888_
timestamp 1688980957
transform -1 0 29348 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _889_
timestamp 1688980957
transform -1 0 29900 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _890_
timestamp 1688980957
transform 1 0 25392 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _891_
timestamp 1688980957
transform 1 0 26864 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _892_
timestamp 1688980957
transform -1 0 29440 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _893_
timestamp 1688980957
transform 1 0 24932 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _894_
timestamp 1688980957
transform 1 0 23000 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _895_
timestamp 1688980957
transform 1 0 24380 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _896_
timestamp 1688980957
transform 1 0 24472 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _897_
timestamp 1688980957
transform -1 0 27324 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _898_
timestamp 1688980957
transform -1 0 28428 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _899_
timestamp 1688980957
transform 1 0 24380 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _900_
timestamp 1688980957
transform 1 0 25852 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _901_
timestamp 1688980957
transform -1 0 28796 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _902_
timestamp 1688980957
transform -1 0 31004 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _903_
timestamp 1688980957
transform 1 0 16652 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _904_
timestamp 1688980957
transform 1 0 17020 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _905_
timestamp 1688980957
transform 1 0 16284 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _906_
timestamp 1688980957
transform 1 0 16560 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _907_
timestamp 1688980957
transform 1 0 16284 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _908_
timestamp 1688980957
transform 1 0 16652 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _909_
timestamp 1688980957
transform 1 0 16652 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _910_
timestamp 1688980957
transform 1 0 17020 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _911_
timestamp 1688980957
transform 1 0 29532 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _912_
timestamp 1688980957
transform 1 0 27600 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _913_
timestamp 1688980957
transform 1 0 28428 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _914_
timestamp 1688980957
transform 1 0 29900 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _915_
timestamp 1688980957
transform -1 0 31464 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _916_
timestamp 1688980957
transform -1 0 31556 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _917_
timestamp 1688980957
transform 1 0 27324 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _918_
timestamp 1688980957
transform 1 0 28244 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _919_
timestamp 1688980957
transform -1 0 31188 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _920_
timestamp 1688980957
transform 1 0 25668 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _921_
timestamp 1688980957
transform 1 0 27140 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _922_
timestamp 1688980957
transform -1 0 31004 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _923_
timestamp 1688980957
transform 1 0 25392 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _924_
timestamp 1688980957
transform -1 0 29440 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _925_
timestamp 1688980957
transform -1 0 27416 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _926_
timestamp 1688980957
transform 1 0 24380 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _927_
timestamp 1688980957
transform -1 0 25760 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _928_
timestamp 1688980957
transform -1 0 26128 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _929_
timestamp 1688980957
transform 1 0 28612 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _930_
timestamp 1688980957
transform 1 0 19688 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _931_
timestamp 1688980957
transform 1 0 21712 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _932_
timestamp 1688980957
transform 1 0 22816 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _933_
timestamp 1688980957
transform 1 0 19596 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _934_
timestamp 1688980957
transform -1 0 24932 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _935_
timestamp 1688980957
transform -1 0 25024 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _936_
timestamp 1688980957
transform 1 0 18768 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _937_
timestamp 1688980957
transform 1 0 19780 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _938_
timestamp 1688980957
transform 1 0 23736 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _939_
timestamp 1688980957
transform 1 0 23092 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _940_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 18492 0 -1 25024
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _941_
timestamp 1688980957
transform 1 0 20056 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _942_
timestamp 1688980957
transform -1 0 23276 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _943_
timestamp 1688980957
transform -1 0 19780 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _944_
timestamp 1688980957
transform -1 0 22724 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _945_
timestamp 1688980957
transform -1 0 23276 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _946_
timestamp 1688980957
transform 1 0 18400 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _947_
timestamp 1688980957
transform -1 0 23276 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _948_
timestamp 1688980957
transform 1 0 21804 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _949_
timestamp 1688980957
transform 1 0 22172 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _950_
timestamp 1688980957
transform -1 0 25576 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _951_
timestamp 1688980957
transform 1 0 22816 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _952_
timestamp 1688980957
transform 1 0 23736 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _953_
timestamp 1688980957
transform 1 0 22264 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _954_
timestamp 1688980957
transform 1 0 21988 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _955_
timestamp 1688980957
transform 1 0 23276 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _956_
timestamp 1688980957
transform 1 0 23368 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _957_
timestamp 1688980957
transform 1 0 16928 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _958_
timestamp 1688980957
transform -1 0 20700 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _959_
timestamp 1688980957
transform 1 0 17020 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _960_
timestamp 1688980957
transform 1 0 17940 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _961_
timestamp 1688980957
transform -1 0 17756 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _962_
timestamp 1688980957
transform 1 0 16100 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _963_
timestamp 1688980957
transform 1 0 16652 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _964_
timestamp 1688980957
transform 1 0 17480 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  _970_
timestamp 1688980957
transform -1 0 34224 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  fanout13
timestamp 1688980957
transform -1 0 23460 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout14
timestamp 1688980957
transform 1 0 23184 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout15
timestamp 1688980957
transform -1 0 24196 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout16
timestamp 1688980957
transform -1 0 27324 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout17
timestamp 1688980957
transform -1 0 33028 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout18
timestamp 1688980957
transform -1 0 31280 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout19
timestamp 1688980957
transform -1 0 33028 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout20
timestamp 1688980957
transform 1 0 32292 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout21
timestamp 1688980957
transform -1 0 23644 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout22
timestamp 1688980957
transform -1 0 23368 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout23 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 23920 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  fanout24
timestamp 1688980957
transform 1 0 31464 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout25
timestamp 1688980957
transform -1 0 32016 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout26
timestamp 1688980957
transform -1 0 33304 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_13 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2300 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_25 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3404 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_29
timestamp 1688980957
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_41
timestamp 1688980957
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_53
timestamp 1688980957
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_57
timestamp 1688980957
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_69
timestamp 1688980957
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_81
timestamp 1688980957
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_85 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 8924 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_90
timestamp 1688980957
transform 1 0 9384 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_102 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 10488 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_110
timestamp 1688980957
transform 1 0 11224 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_113
timestamp 1688980957
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_125
timestamp 1688980957
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_137
timestamp 1688980957
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_141
timestamp 1688980957
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_153
timestamp 1688980957
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_165
timestamp 1688980957
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_169
timestamp 1688980957
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_181
timestamp 1688980957
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_193
timestamp 1688980957
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_203
timestamp 1688980957
transform 1 0 19780 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_215
timestamp 1688980957
transform 1 0 20884 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_223 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 21620 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_225
timestamp 1688980957
transform 1 0 21804 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_237
timestamp 1688980957
transform 1 0 22908 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_249
timestamp 1688980957
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_253
timestamp 1688980957
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_265
timestamp 1688980957
transform 1 0 25484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_277
timestamp 1688980957
transform 1 0 26588 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_281
timestamp 1688980957
transform 1 0 26956 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_293 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 28060 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_300
timestamp 1688980957
transform 1 0 28704 0 1 2176
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_309
timestamp 1688980957
transform 1 0 29532 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_321
timestamp 1688980957
transform 1 0 30636 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_333
timestamp 1688980957
transform 1 0 31740 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_337
timestamp 1688980957
transform 1 0 32108 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_349
timestamp 1688980957
transform 1 0 33212 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 1688980957
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 1688980957
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp 1688980957
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_39
timestamp 1688980957
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_51
timestamp 1688980957
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 1688980957
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_57
timestamp 1688980957
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_69
timestamp 1688980957
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_81
timestamp 1688980957
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_93
timestamp 1688980957
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_105 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_111
timestamp 1688980957
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_113
timestamp 1688980957
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_125
timestamp 1688980957
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_137
timestamp 1688980957
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_149
timestamp 1688980957
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_161
timestamp 1688980957
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_167
timestamp 1688980957
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_169
timestamp 1688980957
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_181
timestamp 1688980957
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_193
timestamp 1688980957
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_205
timestamp 1688980957
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_217
timestamp 1688980957
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_223
timestamp 1688980957
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_225
timestamp 1688980957
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_237
timestamp 1688980957
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_249
timestamp 1688980957
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_261
timestamp 1688980957
transform 1 0 25116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_273
timestamp 1688980957
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_279
timestamp 1688980957
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_281
timestamp 1688980957
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_293
timestamp 1688980957
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_305
timestamp 1688980957
transform 1 0 29164 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_317
timestamp 1688980957
transform 1 0 30268 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_329
timestamp 1688980957
transform 1 0 31372 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_335
timestamp 1688980957
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_337
timestamp 1688980957
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_349
timestamp 1688980957
transform 1 0 33212 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_361
timestamp 1688980957
transform 1 0 34316 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1688980957
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1688980957
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1688980957
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 1688980957
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 1688980957
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_53
timestamp 1688980957
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_65
timestamp 1688980957
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_77
timestamp 1688980957
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 1688980957
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_85
timestamp 1688980957
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_97
timestamp 1688980957
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_109
timestamp 1688980957
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_121
timestamp 1688980957
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_133
timestamp 1688980957
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_139
timestamp 1688980957
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_141
timestamp 1688980957
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_153
timestamp 1688980957
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_165
timestamp 1688980957
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_177
timestamp 1688980957
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_189
timestamp 1688980957
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_195
timestamp 1688980957
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_197
timestamp 1688980957
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_209
timestamp 1688980957
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_221
timestamp 1688980957
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_233
timestamp 1688980957
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_245
timestamp 1688980957
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_251
timestamp 1688980957
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_253
timestamp 1688980957
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_265
timestamp 1688980957
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_277
timestamp 1688980957
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_289
timestamp 1688980957
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_301
timestamp 1688980957
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_307
timestamp 1688980957
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_309
timestamp 1688980957
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_321
timestamp 1688980957
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_333
timestamp 1688980957
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_345
timestamp 1688980957
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_357
timestamp 1688980957
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_363
timestamp 1688980957
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1688980957
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1688980957
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 1688980957
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 1688980957
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 1688980957
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1688980957
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 1688980957
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_69
timestamp 1688980957
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_81
timestamp 1688980957
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_93
timestamp 1688980957
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_105
timestamp 1688980957
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_111
timestamp 1688980957
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_113
timestamp 1688980957
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_125
timestamp 1688980957
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_137
timestamp 1688980957
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_149
timestamp 1688980957
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_161
timestamp 1688980957
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_167
timestamp 1688980957
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_169
timestamp 1688980957
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_181
timestamp 1688980957
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_193
timestamp 1688980957
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_205
timestamp 1688980957
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_217
timestamp 1688980957
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_223
timestamp 1688980957
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_225
timestamp 1688980957
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_237
timestamp 1688980957
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_249
timestamp 1688980957
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_261
timestamp 1688980957
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_273
timestamp 1688980957
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_279
timestamp 1688980957
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_281
timestamp 1688980957
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_293
timestamp 1688980957
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_305
timestamp 1688980957
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_317
timestamp 1688980957
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_329
timestamp 1688980957
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_335
timestamp 1688980957
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_337
timestamp 1688980957
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_349
timestamp 1688980957
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_361
timestamp 1688980957
transform 1 0 34316 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1688980957
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 1688980957
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1688980957
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1688980957
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 1688980957
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_53
timestamp 1688980957
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_65
timestamp 1688980957
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_77
timestamp 1688980957
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 1688980957
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_85
timestamp 1688980957
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_97
timestamp 1688980957
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_109
timestamp 1688980957
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_121
timestamp 1688980957
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_133
timestamp 1688980957
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_139
timestamp 1688980957
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_141
timestamp 1688980957
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_153
timestamp 1688980957
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_165
timestamp 1688980957
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_177
timestamp 1688980957
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_189
timestamp 1688980957
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_195
timestamp 1688980957
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_197
timestamp 1688980957
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_209
timestamp 1688980957
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_221
timestamp 1688980957
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_233
timestamp 1688980957
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_245
timestamp 1688980957
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_251
timestamp 1688980957
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_253
timestamp 1688980957
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_265
timestamp 1688980957
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_277
timestamp 1688980957
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_289
timestamp 1688980957
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_301
timestamp 1688980957
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_307
timestamp 1688980957
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_309
timestamp 1688980957
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_321
timestamp 1688980957
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_333
timestamp 1688980957
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_345
timestamp 1688980957
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_357
timestamp 1688980957
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_363
timestamp 1688980957
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 1688980957
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 1688980957
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_27
timestamp 1688980957
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_39
timestamp 1688980957
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_51
timestamp 1688980957
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 1688980957
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 1688980957
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_69
timestamp 1688980957
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_81
timestamp 1688980957
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_93
timestamp 1688980957
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_105
timestamp 1688980957
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_111
timestamp 1688980957
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_113
timestamp 1688980957
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_125
timestamp 1688980957
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_137
timestamp 1688980957
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_149
timestamp 1688980957
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_161
timestamp 1688980957
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_167
timestamp 1688980957
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_169
timestamp 1688980957
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_181
timestamp 1688980957
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_193
timestamp 1688980957
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_205
timestamp 1688980957
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_217
timestamp 1688980957
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_223
timestamp 1688980957
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_225
timestamp 1688980957
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_237
timestamp 1688980957
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_249
timestamp 1688980957
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_261
timestamp 1688980957
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_273
timestamp 1688980957
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_279
timestamp 1688980957
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_281
timestamp 1688980957
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_293
timestamp 1688980957
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_305
timestamp 1688980957
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_317
timestamp 1688980957
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_329
timestamp 1688980957
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_335
timestamp 1688980957
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_337
timestamp 1688980957
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_349
timestamp 1688980957
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_361
timestamp 1688980957
transform 1 0 34316 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 1688980957
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp 1688980957
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1688980957
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 1688980957
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_41
timestamp 1688980957
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_53
timestamp 1688980957
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_65
timestamp 1688980957
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_77
timestamp 1688980957
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp 1688980957
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_85
timestamp 1688980957
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_97
timestamp 1688980957
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_109
timestamp 1688980957
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_121
timestamp 1688980957
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_133
timestamp 1688980957
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_139
timestamp 1688980957
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_141
timestamp 1688980957
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_153
timestamp 1688980957
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_165
timestamp 1688980957
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_177
timestamp 1688980957
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_189
timestamp 1688980957
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_195
timestamp 1688980957
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_197
timestamp 1688980957
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_209
timestamp 1688980957
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_221
timestamp 1688980957
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_233
timestamp 1688980957
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_245
timestamp 1688980957
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_251
timestamp 1688980957
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_253
timestamp 1688980957
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_265
timestamp 1688980957
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_277
timestamp 1688980957
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_289
timestamp 1688980957
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_301
timestamp 1688980957
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_307
timestamp 1688980957
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_309
timestamp 1688980957
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_321
timestamp 1688980957
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_333
timestamp 1688980957
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_345
timestamp 1688980957
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_357
timestamp 1688980957
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_363
timestamp 1688980957
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 1688980957
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 1688980957
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_27
timestamp 1688980957
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_39
timestamp 1688980957
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_51
timestamp 1688980957
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 1688980957
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_57
timestamp 1688980957
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_69
timestamp 1688980957
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_81
timestamp 1688980957
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_93
timestamp 1688980957
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_105
timestamp 1688980957
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_111
timestamp 1688980957
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_113
timestamp 1688980957
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_125
timestamp 1688980957
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_137
timestamp 1688980957
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_149
timestamp 1688980957
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_161
timestamp 1688980957
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_167
timestamp 1688980957
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_169
timestamp 1688980957
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_181
timestamp 1688980957
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_193
timestamp 1688980957
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_205
timestamp 1688980957
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_217
timestamp 1688980957
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_223
timestamp 1688980957
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_225
timestamp 1688980957
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_237
timestamp 1688980957
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_249
timestamp 1688980957
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_261
timestamp 1688980957
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_273
timestamp 1688980957
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_279
timestamp 1688980957
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_281
timestamp 1688980957
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_293
timestamp 1688980957
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_305
timestamp 1688980957
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_317
timestamp 1688980957
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_329
timestamp 1688980957
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_335
timestamp 1688980957
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_337
timestamp 1688980957
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_349
timestamp 1688980957
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_361
timestamp 1688980957
transform 1 0 34316 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1688980957
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 1688980957
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1688980957
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 1688980957
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_41
timestamp 1688980957
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_53
timestamp 1688980957
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_65
timestamp 1688980957
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_77
timestamp 1688980957
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_83
timestamp 1688980957
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_85
timestamp 1688980957
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_97
timestamp 1688980957
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_109
timestamp 1688980957
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_121
timestamp 1688980957
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_133
timestamp 1688980957
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_139
timestamp 1688980957
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_141
timestamp 1688980957
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_153
timestamp 1688980957
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_165
timestamp 1688980957
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_177
timestamp 1688980957
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_189
timestamp 1688980957
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_195
timestamp 1688980957
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_197
timestamp 1688980957
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_209
timestamp 1688980957
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_221
timestamp 1688980957
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_233
timestamp 1688980957
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_245
timestamp 1688980957
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_251
timestamp 1688980957
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_253
timestamp 1688980957
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_265
timestamp 1688980957
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_277
timestamp 1688980957
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_289
timestamp 1688980957
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_301
timestamp 1688980957
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_307
timestamp 1688980957
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_309
timestamp 1688980957
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_321
timestamp 1688980957
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_333
timestamp 1688980957
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_345
timestamp 1688980957
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_357
timestamp 1688980957
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_363
timestamp 1688980957
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 1688980957
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_15
timestamp 1688980957
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_27
timestamp 1688980957
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_39
timestamp 1688980957
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_51
timestamp 1688980957
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_55
timestamp 1688980957
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_57
timestamp 1688980957
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_69
timestamp 1688980957
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_81
timestamp 1688980957
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_93
timestamp 1688980957
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_105
timestamp 1688980957
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_111
timestamp 1688980957
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_113
timestamp 1688980957
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_125
timestamp 1688980957
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_137
timestamp 1688980957
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_149
timestamp 1688980957
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_161
timestamp 1688980957
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_167
timestamp 1688980957
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_169
timestamp 1688980957
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_181
timestamp 1688980957
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_193
timestamp 1688980957
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_205
timestamp 1688980957
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_217
timestamp 1688980957
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_223
timestamp 1688980957
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_225
timestamp 1688980957
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_237
timestamp 1688980957
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_249
timestamp 1688980957
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_261
timestamp 1688980957
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_273
timestamp 1688980957
transform 1 0 26220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_279
timestamp 1688980957
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_281
timestamp 1688980957
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_293
timestamp 1688980957
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_305
timestamp 1688980957
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_317
timestamp 1688980957
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_329
timestamp 1688980957
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_335
timestamp 1688980957
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_337
timestamp 1688980957
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_349
timestamp 1688980957
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_361
timestamp 1688980957
transform 1 0 34316 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp 1688980957
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_15
timestamp 1688980957
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 1688980957
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_29
timestamp 1688980957
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_41
timestamp 1688980957
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_53
timestamp 1688980957
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_65
timestamp 1688980957
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_77
timestamp 1688980957
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_83
timestamp 1688980957
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_85
timestamp 1688980957
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_97
timestamp 1688980957
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_109
timestamp 1688980957
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_121
timestamp 1688980957
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_133
timestamp 1688980957
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_139
timestamp 1688980957
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_141
timestamp 1688980957
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_153
timestamp 1688980957
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_165
timestamp 1688980957
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_177
timestamp 1688980957
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_189
timestamp 1688980957
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_195
timestamp 1688980957
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_197
timestamp 1688980957
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_209
timestamp 1688980957
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_221
timestamp 1688980957
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_233
timestamp 1688980957
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_245
timestamp 1688980957
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_251
timestamp 1688980957
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_253
timestamp 1688980957
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_265
timestamp 1688980957
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_277
timestamp 1688980957
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_289
timestamp 1688980957
transform 1 0 27692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_301
timestamp 1688980957
transform 1 0 28796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_307
timestamp 1688980957
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_309
timestamp 1688980957
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_321
timestamp 1688980957
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_333
timestamp 1688980957
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_345
timestamp 1688980957
transform 1 0 32844 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_357
timestamp 1688980957
transform 1 0 33948 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_363
timestamp 1688980957
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_3
timestamp 1688980957
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_15
timestamp 1688980957
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_27
timestamp 1688980957
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_39
timestamp 1688980957
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_51
timestamp 1688980957
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_55
timestamp 1688980957
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_57
timestamp 1688980957
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_69
timestamp 1688980957
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_81
timestamp 1688980957
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_93
timestamp 1688980957
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_105
timestamp 1688980957
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_111
timestamp 1688980957
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_113
timestamp 1688980957
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_125
timestamp 1688980957
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_137
timestamp 1688980957
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_149
timestamp 1688980957
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_161
timestamp 1688980957
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_167
timestamp 1688980957
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_169
timestamp 1688980957
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_181
timestamp 1688980957
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_193
timestamp 1688980957
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_205
timestamp 1688980957
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_217
timestamp 1688980957
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_223
timestamp 1688980957
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_225
timestamp 1688980957
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_237
timestamp 1688980957
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_249
timestamp 1688980957
transform 1 0 24012 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_261
timestamp 1688980957
transform 1 0 25116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_273
timestamp 1688980957
transform 1 0 26220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_279
timestamp 1688980957
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_281
timestamp 1688980957
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_293
timestamp 1688980957
transform 1 0 28060 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_305
timestamp 1688980957
transform 1 0 29164 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_317
timestamp 1688980957
transform 1 0 30268 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_329
timestamp 1688980957
transform 1 0 31372 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_335
timestamp 1688980957
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_337
timestamp 1688980957
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_349
timestamp 1688980957
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_361
timestamp 1688980957
transform 1 0 34316 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_3
timestamp 1688980957
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_15
timestamp 1688980957
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 1688980957
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_29
timestamp 1688980957
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_41
timestamp 1688980957
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_53
timestamp 1688980957
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_65
timestamp 1688980957
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_77
timestamp 1688980957
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_83
timestamp 1688980957
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_85
timestamp 1688980957
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_97
timestamp 1688980957
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_109
timestamp 1688980957
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_121
timestamp 1688980957
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_133
timestamp 1688980957
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_139
timestamp 1688980957
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_141
timestamp 1688980957
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_153
timestamp 1688980957
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_165
timestamp 1688980957
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_177
timestamp 1688980957
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_189
timestamp 1688980957
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_195
timestamp 1688980957
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_197
timestamp 1688980957
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_209
timestamp 1688980957
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_221
timestamp 1688980957
transform 1 0 21436 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_233
timestamp 1688980957
transform 1 0 22540 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_245
timestamp 1688980957
transform 1 0 23644 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_251
timestamp 1688980957
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_253
timestamp 1688980957
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_265
timestamp 1688980957
transform 1 0 25484 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_277
timestamp 1688980957
transform 1 0 26588 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_289
timestamp 1688980957
transform 1 0 27692 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_301
timestamp 1688980957
transform 1 0 28796 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_307
timestamp 1688980957
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_309
timestamp 1688980957
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_321
timestamp 1688980957
transform 1 0 30636 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_333
timestamp 1688980957
transform 1 0 31740 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_345
timestamp 1688980957
transform 1 0 32844 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_357
timestamp 1688980957
transform 1 0 33948 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_363
timestamp 1688980957
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_3
timestamp 1688980957
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_15
timestamp 1688980957
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_27
timestamp 1688980957
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_39
timestamp 1688980957
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_51
timestamp 1688980957
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_55
timestamp 1688980957
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_57
timestamp 1688980957
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_69
timestamp 1688980957
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_81
timestamp 1688980957
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_93
timestamp 1688980957
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_105
timestamp 1688980957
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_111
timestamp 1688980957
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_113
timestamp 1688980957
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_125
timestamp 1688980957
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_137
timestamp 1688980957
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_149
timestamp 1688980957
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_161
timestamp 1688980957
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_167
timestamp 1688980957
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_169
timestamp 1688980957
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_181
timestamp 1688980957
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_193
timestamp 1688980957
transform 1 0 18860 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_205
timestamp 1688980957
transform 1 0 19964 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_217
timestamp 1688980957
transform 1 0 21068 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_223
timestamp 1688980957
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_225
timestamp 1688980957
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_237
timestamp 1688980957
transform 1 0 22908 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_249
timestamp 1688980957
transform 1 0 24012 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_261
timestamp 1688980957
transform 1 0 25116 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_273
timestamp 1688980957
transform 1 0 26220 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_279
timestamp 1688980957
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_281
timestamp 1688980957
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_293
timestamp 1688980957
transform 1 0 28060 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_305
timestamp 1688980957
transform 1 0 29164 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_317
timestamp 1688980957
transform 1 0 30268 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_329
timestamp 1688980957
transform 1 0 31372 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_335
timestamp 1688980957
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_337
timestamp 1688980957
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_349
timestamp 1688980957
transform 1 0 33212 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_361
timestamp 1688980957
transform 1 0 34316 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_6
timestamp 1688980957
transform 1 0 1656 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_18
timestamp 1688980957
transform 1 0 2760 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_26
timestamp 1688980957
transform 1 0 3496 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_29
timestamp 1688980957
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_41
timestamp 1688980957
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_53
timestamp 1688980957
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_65
timestamp 1688980957
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_77
timestamp 1688980957
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_83
timestamp 1688980957
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_85
timestamp 1688980957
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_97
timestamp 1688980957
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_109
timestamp 1688980957
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_121
timestamp 1688980957
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_133
timestamp 1688980957
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_139
timestamp 1688980957
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_141
timestamp 1688980957
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_153
timestamp 1688980957
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_165
timestamp 1688980957
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_177
timestamp 1688980957
transform 1 0 17388 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_189
timestamp 1688980957
transform 1 0 18492 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_195
timestamp 1688980957
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_197
timestamp 1688980957
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_209
timestamp 1688980957
transform 1 0 20332 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_221
timestamp 1688980957
transform 1 0 21436 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_233
timestamp 1688980957
transform 1 0 22540 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_245
timestamp 1688980957
transform 1 0 23644 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_251
timestamp 1688980957
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_253
timestamp 1688980957
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_265
timestamp 1688980957
transform 1 0 25484 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_277
timestamp 1688980957
transform 1 0 26588 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_289
timestamp 1688980957
transform 1 0 27692 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_301
timestamp 1688980957
transform 1 0 28796 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_307
timestamp 1688980957
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_309
timestamp 1688980957
transform 1 0 29532 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_321
timestamp 1688980957
transform 1 0 30636 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_333
timestamp 1688980957
transform 1 0 31740 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_345
timestamp 1688980957
transform 1 0 32844 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_357
timestamp 1688980957
transform 1 0 33948 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_363
timestamp 1688980957
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_3
timestamp 1688980957
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_15
timestamp 1688980957
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_27
timestamp 1688980957
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_39
timestamp 1688980957
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_51
timestamp 1688980957
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_55
timestamp 1688980957
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_57
timestamp 1688980957
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_69
timestamp 1688980957
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_81
timestamp 1688980957
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_93
timestamp 1688980957
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_105
timestamp 1688980957
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_111
timestamp 1688980957
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_113
timestamp 1688980957
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_125
timestamp 1688980957
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_137
timestamp 1688980957
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_149
timestamp 1688980957
transform 1 0 14812 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_161
timestamp 1688980957
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_167
timestamp 1688980957
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_169
timestamp 1688980957
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_181
timestamp 1688980957
transform 1 0 17756 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_193
timestamp 1688980957
transform 1 0 18860 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_205
timestamp 1688980957
transform 1 0 19964 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_217
timestamp 1688980957
transform 1 0 21068 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_223
timestamp 1688980957
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_225
timestamp 1688980957
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_237
timestamp 1688980957
transform 1 0 22908 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_249
timestamp 1688980957
transform 1 0 24012 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_261
timestamp 1688980957
transform 1 0 25116 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_273
timestamp 1688980957
transform 1 0 26220 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_279
timestamp 1688980957
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_281
timestamp 1688980957
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_293
timestamp 1688980957
transform 1 0 28060 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_305
timestamp 1688980957
transform 1 0 29164 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_317
timestamp 1688980957
transform 1 0 30268 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_329
timestamp 1688980957
transform 1 0 31372 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_335
timestamp 1688980957
transform 1 0 31924 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_337
timestamp 1688980957
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_349
timestamp 1688980957
transform 1 0 33212 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_361
timestamp 1688980957
transform 1 0 34316 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_3
timestamp 1688980957
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_15
timestamp 1688980957
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_27
timestamp 1688980957
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_29
timestamp 1688980957
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_41
timestamp 1688980957
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_53
timestamp 1688980957
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_65
timestamp 1688980957
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_77
timestamp 1688980957
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_83
timestamp 1688980957
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_85
timestamp 1688980957
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_97
timestamp 1688980957
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_109
timestamp 1688980957
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_121
timestamp 1688980957
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_133
timestamp 1688980957
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_139
timestamp 1688980957
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_141
timestamp 1688980957
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_153
timestamp 1688980957
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_165
timestamp 1688980957
transform 1 0 16284 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_177
timestamp 1688980957
transform 1 0 17388 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_189
timestamp 1688980957
transform 1 0 18492 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_195
timestamp 1688980957
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_197
timestamp 1688980957
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_209
timestamp 1688980957
transform 1 0 20332 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_221
timestamp 1688980957
transform 1 0 21436 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_233
timestamp 1688980957
transform 1 0 22540 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_245
timestamp 1688980957
transform 1 0 23644 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_251
timestamp 1688980957
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_253
timestamp 1688980957
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_265
timestamp 1688980957
transform 1 0 25484 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_277
timestamp 1688980957
transform 1 0 26588 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_289
timestamp 1688980957
transform 1 0 27692 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_301
timestamp 1688980957
transform 1 0 28796 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_307
timestamp 1688980957
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_309
timestamp 1688980957
transform 1 0 29532 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_321
timestamp 1688980957
transform 1 0 30636 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_333
timestamp 1688980957
transform 1 0 31740 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_345
timestamp 1688980957
transform 1 0 32844 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_357
timestamp 1688980957
transform 1 0 33948 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_363
timestamp 1688980957
transform 1 0 34500 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_3
timestamp 1688980957
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_15
timestamp 1688980957
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_27
timestamp 1688980957
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_39
timestamp 1688980957
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_51
timestamp 1688980957
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_55
timestamp 1688980957
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_57
timestamp 1688980957
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_69
timestamp 1688980957
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_81
timestamp 1688980957
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_93
timestamp 1688980957
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_105
timestamp 1688980957
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_111
timestamp 1688980957
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_113
timestamp 1688980957
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_125
timestamp 1688980957
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_137
timestamp 1688980957
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_149
timestamp 1688980957
transform 1 0 14812 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_161
timestamp 1688980957
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_167
timestamp 1688980957
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_169
timestamp 1688980957
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_181
timestamp 1688980957
transform 1 0 17756 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_193
timestamp 1688980957
transform 1 0 18860 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_205
timestamp 1688980957
transform 1 0 19964 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_217
timestamp 1688980957
transform 1 0 21068 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_223
timestamp 1688980957
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_225
timestamp 1688980957
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_237
timestamp 1688980957
transform 1 0 22908 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_249
timestamp 1688980957
transform 1 0 24012 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_261
timestamp 1688980957
transform 1 0 25116 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_273
timestamp 1688980957
transform 1 0 26220 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_279
timestamp 1688980957
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_281
timestamp 1688980957
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_293
timestamp 1688980957
transform 1 0 28060 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_305
timestamp 1688980957
transform 1 0 29164 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_317
timestamp 1688980957
transform 1 0 30268 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_329
timestamp 1688980957
transform 1 0 31372 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_335
timestamp 1688980957
transform 1 0 31924 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_337
timestamp 1688980957
transform 1 0 32108 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_349
timestamp 1688980957
transform 1 0 33212 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_357
timestamp 1688980957
transform 1 0 33948 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_3
timestamp 1688980957
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_15
timestamp 1688980957
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_27
timestamp 1688980957
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_29
timestamp 1688980957
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_41
timestamp 1688980957
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_53
timestamp 1688980957
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_65
timestamp 1688980957
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_77
timestamp 1688980957
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_83
timestamp 1688980957
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_85
timestamp 1688980957
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_97
timestamp 1688980957
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_109
timestamp 1688980957
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_121
timestamp 1688980957
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_133
timestamp 1688980957
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_139
timestamp 1688980957
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_141
timestamp 1688980957
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_153
timestamp 1688980957
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_165
timestamp 1688980957
transform 1 0 16284 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_177
timestamp 1688980957
transform 1 0 17388 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_189
timestamp 1688980957
transform 1 0 18492 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_195
timestamp 1688980957
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_197
timestamp 1688980957
transform 1 0 19228 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_209
timestamp 1688980957
transform 1 0 20332 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_221
timestamp 1688980957
transform 1 0 21436 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_233
timestamp 1688980957
transform 1 0 22540 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_245
timestamp 1688980957
transform 1 0 23644 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_251
timestamp 1688980957
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_253
timestamp 1688980957
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_265
timestamp 1688980957
transform 1 0 25484 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_277
timestamp 1688980957
transform 1 0 26588 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_289
timestamp 1688980957
transform 1 0 27692 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_301
timestamp 1688980957
transform 1 0 28796 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_307
timestamp 1688980957
transform 1 0 29348 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_309
timestamp 1688980957
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_321
timestamp 1688980957
transform 1 0 30636 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_333
timestamp 1688980957
transform 1 0 31740 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_345
timestamp 1688980957
transform 1 0 32844 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_360
timestamp 1688980957
transform 1 0 34224 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_3
timestamp 1688980957
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_15
timestamp 1688980957
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_27
timestamp 1688980957
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_39
timestamp 1688980957
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_51
timestamp 1688980957
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_55
timestamp 1688980957
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_57
timestamp 1688980957
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_69
timestamp 1688980957
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_81
timestamp 1688980957
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_93
timestamp 1688980957
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_105
timestamp 1688980957
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_111
timestamp 1688980957
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_113
timestamp 1688980957
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_125
timestamp 1688980957
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_137
timestamp 1688980957
transform 1 0 13708 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_149
timestamp 1688980957
transform 1 0 14812 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_161
timestamp 1688980957
transform 1 0 15916 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_167
timestamp 1688980957
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_169
timestamp 1688980957
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_181
timestamp 1688980957
transform 1 0 17756 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_193
timestamp 1688980957
transform 1 0 18860 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_205
timestamp 1688980957
transform 1 0 19964 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_217
timestamp 1688980957
transform 1 0 21068 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_223
timestamp 1688980957
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_225
timestamp 1688980957
transform 1 0 21804 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_237
timestamp 1688980957
transform 1 0 22908 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_249
timestamp 1688980957
transform 1 0 24012 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_261
timestamp 1688980957
transform 1 0 25116 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_273
timestamp 1688980957
transform 1 0 26220 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_279
timestamp 1688980957
transform 1 0 26772 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_281
timestamp 1688980957
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_293
timestamp 1688980957
transform 1 0 28060 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_305
timestamp 1688980957
transform 1 0 29164 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_317
timestamp 1688980957
transform 1 0 30268 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_329
timestamp 1688980957
transform 1 0 31372 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_335
timestamp 1688980957
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_337
timestamp 1688980957
transform 1 0 32108 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_349
timestamp 1688980957
transform 1 0 33212 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_361
timestamp 1688980957
transform 1 0 34316 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_3
timestamp 1688980957
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_15
timestamp 1688980957
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_27
timestamp 1688980957
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_29
timestamp 1688980957
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_41
timestamp 1688980957
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_53
timestamp 1688980957
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_65
timestamp 1688980957
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_77
timestamp 1688980957
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_83
timestamp 1688980957
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_85
timestamp 1688980957
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_97
timestamp 1688980957
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_109
timestamp 1688980957
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_121
timestamp 1688980957
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_133
timestamp 1688980957
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_139
timestamp 1688980957
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_141
timestamp 1688980957
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_153
timestamp 1688980957
transform 1 0 15180 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_165
timestamp 1688980957
transform 1 0 16284 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_177
timestamp 1688980957
transform 1 0 17388 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_189
timestamp 1688980957
transform 1 0 18492 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_195
timestamp 1688980957
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_197
timestamp 1688980957
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_209
timestamp 1688980957
transform 1 0 20332 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_221
timestamp 1688980957
transform 1 0 21436 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_233
timestamp 1688980957
transform 1 0 22540 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_245
timestamp 1688980957
transform 1 0 23644 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_251
timestamp 1688980957
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_253
timestamp 1688980957
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_265
timestamp 1688980957
transform 1 0 25484 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_277
timestamp 1688980957
transform 1 0 26588 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_289
timestamp 1688980957
transform 1 0 27692 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_301
timestamp 1688980957
transform 1 0 28796 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_307
timestamp 1688980957
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_309
timestamp 1688980957
transform 1 0 29532 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_321
timestamp 1688980957
transform 1 0 30636 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_333
timestamp 1688980957
transform 1 0 31740 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_345
timestamp 1688980957
transform 1 0 32844 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_357
timestamp 1688980957
transform 1 0 33948 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_363
timestamp 1688980957
transform 1 0 34500 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_3
timestamp 1688980957
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_15
timestamp 1688980957
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_27
timestamp 1688980957
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_39
timestamp 1688980957
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_51
timestamp 1688980957
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_55
timestamp 1688980957
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_57
timestamp 1688980957
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_69
timestamp 1688980957
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_81
timestamp 1688980957
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_93
timestamp 1688980957
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_105
timestamp 1688980957
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_111
timestamp 1688980957
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_113
timestamp 1688980957
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_125
timestamp 1688980957
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_137
timestamp 1688980957
transform 1 0 13708 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_149
timestamp 1688980957
transform 1 0 14812 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_161
timestamp 1688980957
transform 1 0 15916 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_167
timestamp 1688980957
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_169
timestamp 1688980957
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_181
timestamp 1688980957
transform 1 0 17756 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_193
timestamp 1688980957
transform 1 0 18860 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_205
timestamp 1688980957
transform 1 0 19964 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_217
timestamp 1688980957
transform 1 0 21068 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_223
timestamp 1688980957
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_225
timestamp 1688980957
transform 1 0 21804 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_237
timestamp 1688980957
transform 1 0 22908 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_249
timestamp 1688980957
transform 1 0 24012 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_261
timestamp 1688980957
transform 1 0 25116 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_273
timestamp 1688980957
transform 1 0 26220 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_279
timestamp 1688980957
transform 1 0 26772 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_281
timestamp 1688980957
transform 1 0 26956 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_293
timestamp 1688980957
transform 1 0 28060 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_305
timestamp 1688980957
transform 1 0 29164 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_317
timestamp 1688980957
transform 1 0 30268 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_329
timestamp 1688980957
transform 1 0 31372 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_335
timestamp 1688980957
transform 1 0 31924 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_337
timestamp 1688980957
transform 1 0 32108 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_349
timestamp 1688980957
transform 1 0 33212 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_361
timestamp 1688980957
transform 1 0 34316 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_3
timestamp 1688980957
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_15
timestamp 1688980957
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_27
timestamp 1688980957
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_29
timestamp 1688980957
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_41
timestamp 1688980957
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_53
timestamp 1688980957
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_65
timestamp 1688980957
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_77
timestamp 1688980957
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_83
timestamp 1688980957
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_85
timestamp 1688980957
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_97
timestamp 1688980957
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_109
timestamp 1688980957
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_121
timestamp 1688980957
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_133
timestamp 1688980957
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_139
timestamp 1688980957
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_141
timestamp 1688980957
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_153
timestamp 1688980957
transform 1 0 15180 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_165
timestamp 1688980957
transform 1 0 16284 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_177
timestamp 1688980957
transform 1 0 17388 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_189
timestamp 1688980957
transform 1 0 18492 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_195
timestamp 1688980957
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_197
timestamp 1688980957
transform 1 0 19228 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_209
timestamp 1688980957
transform 1 0 20332 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_221
timestamp 1688980957
transform 1 0 21436 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_229
timestamp 1688980957
transform 1 0 22172 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_237
timestamp 1688980957
transform 1 0 22908 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_243
timestamp 1688980957
transform 1 0 23460 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_251
timestamp 1688980957
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_256
timestamp 1688980957
transform 1 0 24656 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_273
timestamp 1688980957
transform 1 0 26220 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_285
timestamp 1688980957
transform 1 0 27324 0 1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_296
timestamp 1688980957
transform 1 0 28336 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_309
timestamp 1688980957
transform 1 0 29532 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_321
timestamp 1688980957
transform 1 0 30636 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_333
timestamp 1688980957
transform 1 0 31740 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_345
timestamp 1688980957
transform 1 0 32844 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_357
timestamp 1688980957
transform 1 0 33948 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_363
timestamp 1688980957
transform 1 0 34500 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_3
timestamp 1688980957
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_15
timestamp 1688980957
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_27
timestamp 1688980957
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_39
timestamp 1688980957
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_51
timestamp 1688980957
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_55
timestamp 1688980957
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_57
timestamp 1688980957
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_69
timestamp 1688980957
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_81
timestamp 1688980957
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_93
timestamp 1688980957
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_105
timestamp 1688980957
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_111
timestamp 1688980957
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_113
timestamp 1688980957
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_125
timestamp 1688980957
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_137
timestamp 1688980957
transform 1 0 13708 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_149
timestamp 1688980957
transform 1 0 14812 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_161
timestamp 1688980957
transform 1 0 15916 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_167
timestamp 1688980957
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_169
timestamp 1688980957
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_181
timestamp 1688980957
transform 1 0 17756 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_193
timestamp 1688980957
transform 1 0 18860 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_201
timestamp 1688980957
transform 1 0 19596 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_219
timestamp 1688980957
transform 1 0 21252 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_223
timestamp 1688980957
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_225
timestamp 1688980957
transform 1 0 21804 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_237
timestamp 1688980957
transform 1 0 22908 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_279
timestamp 1688980957
transform 1 0 26772 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_281
timestamp 1688980957
transform 1 0 26956 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_287
timestamp 1688980957
transform 1 0 27508 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_304
timestamp 1688980957
transform 1 0 29072 0 -1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_315
timestamp 1688980957
transform 1 0 30084 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_327
timestamp 1688980957
transform 1 0 31188 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_333
timestamp 1688980957
transform 1 0 31740 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_337
timestamp 1688980957
transform 1 0 32108 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_349
timestamp 1688980957
transform 1 0 33212 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_361
timestamp 1688980957
transform 1 0 34316 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_3
timestamp 1688980957
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_15
timestamp 1688980957
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_27
timestamp 1688980957
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_29
timestamp 1688980957
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_41
timestamp 1688980957
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_53
timestamp 1688980957
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_65
timestamp 1688980957
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_77
timestamp 1688980957
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_83
timestamp 1688980957
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_85
timestamp 1688980957
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_97
timestamp 1688980957
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_109
timestamp 1688980957
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_121
timestamp 1688980957
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_133
timestamp 1688980957
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_139
timestamp 1688980957
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_141
timestamp 1688980957
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_153
timestamp 1688980957
transform 1 0 15180 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_165
timestamp 1688980957
transform 1 0 16284 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_177
timestamp 1688980957
transform 1 0 17388 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_189
timestamp 1688980957
transform 1 0 18492 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_195
timestamp 1688980957
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_197
timestamp 1688980957
transform 1 0 19228 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_209
timestamp 1688980957
transform 1 0 20332 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_221
timestamp 1688980957
transform 1 0 21436 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_233
timestamp 1688980957
transform 1 0 22540 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_245
timestamp 1688980957
transform 1 0 23644 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_285
timestamp 1688980957
transform 1 0 27324 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_291
timestamp 1688980957
transform 1 0 27876 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_295
timestamp 1688980957
transform 1 0 28244 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_306
timestamp 1688980957
transform 1 0 29256 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_312
timestamp 1688980957
transform 1 0 29808 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_333
timestamp 1688980957
transform 1 0 31740 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_345
timestamp 1688980957
transform 1 0 32844 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_357
timestamp 1688980957
transform 1 0 33948 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_363
timestamp 1688980957
transform 1 0 34500 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_3
timestamp 1688980957
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_15
timestamp 1688980957
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_27
timestamp 1688980957
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_39
timestamp 1688980957
transform 1 0 4692 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_51
timestamp 1688980957
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_55
timestamp 1688980957
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_57
timestamp 1688980957
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_69
timestamp 1688980957
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_81
timestamp 1688980957
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_93
timestamp 1688980957
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_105
timestamp 1688980957
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_111
timestamp 1688980957
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_113
timestamp 1688980957
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_125
timestamp 1688980957
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_137
timestamp 1688980957
transform 1 0 13708 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_149
timestamp 1688980957
transform 1 0 14812 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_161
timestamp 1688980957
transform 1 0 15916 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_167
timestamp 1688980957
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_169
timestamp 1688980957
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_181
timestamp 1688980957
transform 1 0 17756 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_188
timestamp 1688980957
transform 1 0 18400 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_211
timestamp 1688980957
transform 1 0 20516 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_223
timestamp 1688980957
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_225
timestamp 1688980957
transform 1 0 21804 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_237
timestamp 1688980957
transform 1 0 22908 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_249
timestamp 1688980957
transform 1 0 24012 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_253
timestamp 1688980957
transform 1 0 24380 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_264
timestamp 1688980957
transform 1 0 25392 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_273
timestamp 1688980957
transform 1 0 26220 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_334
timestamp 1688980957
transform 1 0 31832 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_337
timestamp 1688980957
transform 1 0 32108 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_349
timestamp 1688980957
transform 1 0 33212 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_361
timestamp 1688980957
transform 1 0 34316 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_3
timestamp 1688980957
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_15
timestamp 1688980957
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_27
timestamp 1688980957
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_29
timestamp 1688980957
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_41
timestamp 1688980957
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_53
timestamp 1688980957
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_65
timestamp 1688980957
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_77
timestamp 1688980957
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_83
timestamp 1688980957
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_85
timestamp 1688980957
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_97
timestamp 1688980957
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_109
timestamp 1688980957
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_121
timestamp 1688980957
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_133
timestamp 1688980957
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_139
timestamp 1688980957
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_141
timestamp 1688980957
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_153
timestamp 1688980957
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_165
timestamp 1688980957
transform 1 0 16284 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_177
timestamp 1688980957
transform 1 0 17388 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_194
timestamp 1688980957
transform 1 0 18952 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_206
timestamp 1688980957
transform 1 0 20056 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_247
timestamp 1688980957
transform 1 0 23828 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_251
timestamp 1688980957
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_253
timestamp 1688980957
transform 1 0 24380 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_265
timestamp 1688980957
transform 1 0 25484 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_280
timestamp 1688980957
transform 1 0 26864 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_292
timestamp 1688980957
transform 1 0 27968 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_298
timestamp 1688980957
transform 1 0 28520 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_321
timestamp 1688980957
transform 1 0 30636 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_338
timestamp 1688980957
transform 1 0 32200 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_350
timestamp 1688980957
transform 1 0 33304 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_362
timestamp 1688980957
transform 1 0 34408 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_3
timestamp 1688980957
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_15
timestamp 1688980957
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_27
timestamp 1688980957
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_39
timestamp 1688980957
transform 1 0 4692 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_51
timestamp 1688980957
transform 1 0 5796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_55
timestamp 1688980957
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_57
timestamp 1688980957
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_69
timestamp 1688980957
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_81
timestamp 1688980957
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_93
timestamp 1688980957
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_105
timestamp 1688980957
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_111
timestamp 1688980957
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_113
timestamp 1688980957
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_125
timestamp 1688980957
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_137
timestamp 1688980957
transform 1 0 13708 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_149
timestamp 1688980957
transform 1 0 14812 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_160
timestamp 1688980957
transform 1 0 15824 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_166
timestamp 1688980957
transform 1 0 16376 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_189
timestamp 1688980957
transform 1 0 18492 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_199
timestamp 1688980957
transform 1 0 19412 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_225
timestamp 1688980957
transform 1 0 21804 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_234
timestamp 1688980957
transform 1 0 22632 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_265
timestamp 1688980957
transform 1 0 25484 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_278
timestamp 1688980957
transform 1 0 26680 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_286
timestamp 1688980957
transform 1 0 27416 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_298
timestamp 1688980957
transform 1 0 28520 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_314
timestamp 1688980957
transform 1 0 29992 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_320
timestamp 1688980957
transform 1 0 30544 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_324
timestamp 1688980957
transform 1 0 30912 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_337
timestamp 1688980957
transform 1 0 32108 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_349
timestamp 1688980957
transform 1 0 33212 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_361
timestamp 1688980957
transform 1 0 34316 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_3
timestamp 1688980957
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_15
timestamp 1688980957
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_27
timestamp 1688980957
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_29
timestamp 1688980957
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_41
timestamp 1688980957
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_53
timestamp 1688980957
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_65
timestamp 1688980957
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_77
timestamp 1688980957
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_83
timestamp 1688980957
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_85
timestamp 1688980957
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_97
timestamp 1688980957
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_109
timestamp 1688980957
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_121
timestamp 1688980957
transform 1 0 12236 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_133
timestamp 1688980957
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_139
timestamp 1688980957
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_141
timestamp 1688980957
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_189
timestamp 1688980957
transform 1 0 18492 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_195
timestamp 1688980957
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_200
timestamp 1688980957
transform 1 0 19504 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_204
timestamp 1688980957
transform 1 0 19872 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_226
timestamp 1688980957
transform 1 0 21896 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_250
timestamp 1688980957
transform 1 0 24104 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_301
timestamp 1688980957
transform 1 0 28796 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_307
timestamp 1688980957
transform 1 0 29348 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_309
timestamp 1688980957
transform 1 0 29532 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_313
timestamp 1688980957
transform 1 0 29900 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_331
timestamp 1688980957
transform 1 0 31556 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_343
timestamp 1688980957
transform 1 0 32660 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_355
timestamp 1688980957
transform 1 0 33764 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_363
timestamp 1688980957
transform 1 0 34500 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_3
timestamp 1688980957
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_15
timestamp 1688980957
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_27
timestamp 1688980957
transform 1 0 3588 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_39
timestamp 1688980957
transform 1 0 4692 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_51
timestamp 1688980957
transform 1 0 5796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_55
timestamp 1688980957
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_57
timestamp 1688980957
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_69
timestamp 1688980957
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_81
timestamp 1688980957
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_93
timestamp 1688980957
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_105
timestamp 1688980957
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_111
timestamp 1688980957
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_113
timestamp 1688980957
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_125
timestamp 1688980957
transform 1 0 12604 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_137
timestamp 1688980957
transform 1 0 13708 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_149
timestamp 1688980957
transform 1 0 14812 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_161
timestamp 1688980957
transform 1 0 15916 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_167
timestamp 1688980957
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_169
timestamp 1688980957
transform 1 0 16652 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_186
timestamp 1688980957
transform 1 0 18216 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_197
timestamp 1688980957
transform 1 0 19228 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_209
timestamp 1688980957
transform 1 0 20332 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_219
timestamp 1688980957
transform 1 0 21252 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_223
timestamp 1688980957
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_225
timestamp 1688980957
transform 1 0 21804 0 -1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_236
timestamp 1688980957
transform 1 0 22816 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_248
timestamp 1688980957
transform 1 0 23920 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_256
timestamp 1688980957
transform 1 0 24656 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_260
timestamp 1688980957
transform 1 0 25024 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_264
timestamp 1688980957
transform 1 0 25392 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_278
timestamp 1688980957
transform 1 0 26680 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_284
timestamp 1688980957
transform 1 0 27232 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_327
timestamp 1688980957
transform 1 0 31188 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_335
timestamp 1688980957
transform 1 0 31924 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_337
timestamp 1688980957
transform 1 0 32108 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_349
timestamp 1688980957
transform 1 0 33212 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_361
timestamp 1688980957
transform 1 0 34316 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_3
timestamp 1688980957
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_15
timestamp 1688980957
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_27
timestamp 1688980957
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_29
timestamp 1688980957
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_41
timestamp 1688980957
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_53
timestamp 1688980957
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_65
timestamp 1688980957
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_77
timestamp 1688980957
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_83
timestamp 1688980957
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_85
timestamp 1688980957
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_97
timestamp 1688980957
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_109
timestamp 1688980957
transform 1 0 11132 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_121
timestamp 1688980957
transform 1 0 12236 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_133
timestamp 1688980957
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_139
timestamp 1688980957
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_141
timestamp 1688980957
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_153
timestamp 1688980957
transform 1 0 15180 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_161
timestamp 1688980957
transform 1 0 15916 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_185
timestamp 1688980957
transform 1 0 18124 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_206
timestamp 1688980957
transform 1 0 20056 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_215
timestamp 1688980957
transform 1 0 20884 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_226
timestamp 1688980957
transform 1 0 21896 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_234
timestamp 1688980957
transform 1 0 22632 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_239
timestamp 1688980957
transform 1 0 23092 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_248
timestamp 1688980957
transform 1 0 23920 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_253
timestamp 1688980957
transform 1 0 24380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_265
timestamp 1688980957
transform 1 0 25484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_277
timestamp 1688980957
transform 1 0 26588 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_306
timestamp 1688980957
transform 1 0 29256 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_323
timestamp 1688980957
transform 1 0 30820 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_332
timestamp 1688980957
transform 1 0 31648 0 1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_343
timestamp 1688980957
transform 1 0 32660 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_355
timestamp 1688980957
transform 1 0 33764 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_363
timestamp 1688980957
transform 1 0 34500 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_3
timestamp 1688980957
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_15
timestamp 1688980957
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_27
timestamp 1688980957
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_39
timestamp 1688980957
transform 1 0 4692 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_51
timestamp 1688980957
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_55
timestamp 1688980957
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_57
timestamp 1688980957
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_69
timestamp 1688980957
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_81
timestamp 1688980957
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_93
timestamp 1688980957
transform 1 0 9660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_105
timestamp 1688980957
transform 1 0 10764 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_111
timestamp 1688980957
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_113
timestamp 1688980957
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_125
timestamp 1688980957
transform 1 0 12604 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_137
timestamp 1688980957
transform 1 0 13708 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_149
timestamp 1688980957
transform 1 0 14812 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_161
timestamp 1688980957
transform 1 0 15916 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_167
timestamp 1688980957
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_169
timestamp 1688980957
transform 1 0 16652 0 -1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_178
timestamp 1688980957
transform 1 0 17480 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_190
timestamp 1688980957
transform 1 0 18584 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_198
timestamp 1688980957
transform 1 0 19320 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_238
timestamp 1688980957
transform 1 0 23000 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_275
timestamp 1688980957
transform 1 0 26404 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_279
timestamp 1688980957
transform 1 0 26772 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_286
timestamp 1688980957
transform 1 0 27416 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_294
timestamp 1688980957
transform 1 0 28152 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_298
timestamp 1688980957
transform 1 0 28520 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_308
timestamp 1688980957
transform 1 0 29440 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_316
timestamp 1688980957
transform 1 0 30176 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_337
timestamp 1688980957
transform 1 0 32108 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_355
timestamp 1688980957
transform 1 0 33764 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_363
timestamp 1688980957
transform 1 0 34500 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_6
timestamp 1688980957
transform 1 0 1656 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_18
timestamp 1688980957
transform 1 0 2760 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_26
timestamp 1688980957
transform 1 0 3496 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_29
timestamp 1688980957
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_41
timestamp 1688980957
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_53
timestamp 1688980957
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_65
timestamp 1688980957
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_77
timestamp 1688980957
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_83
timestamp 1688980957
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_85
timestamp 1688980957
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_97
timestamp 1688980957
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_109
timestamp 1688980957
transform 1 0 11132 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_121
timestamp 1688980957
transform 1 0 12236 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_133
timestamp 1688980957
transform 1 0 13340 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_139
timestamp 1688980957
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_141
timestamp 1688980957
transform 1 0 14076 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_153
timestamp 1688980957
transform 1 0 15180 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_192
timestamp 1688980957
transform 1 0 18768 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_202
timestamp 1688980957
transform 1 0 19688 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_207
timestamp 1688980957
transform 1 0 20148 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_215
timestamp 1688980957
transform 1 0 20884 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_253
timestamp 1688980957
transform 1 0 24380 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_261
timestamp 1688980957
transform 1 0 25116 0 1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_296
timestamp 1688980957
transform 1 0 28336 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_353
timestamp 1688980957
transform 1 0 33580 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_361
timestamp 1688980957
transform 1 0 34316 0 1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_3
timestamp 1688980957
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_15
timestamp 1688980957
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_27
timestamp 1688980957
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_39
timestamp 1688980957
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_51
timestamp 1688980957
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_55
timestamp 1688980957
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_57
timestamp 1688980957
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_69
timestamp 1688980957
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_81
timestamp 1688980957
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_93
timestamp 1688980957
transform 1 0 9660 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_105
timestamp 1688980957
transform 1 0 10764 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_111
timestamp 1688980957
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_113
timestamp 1688980957
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_125
timestamp 1688980957
transform 1 0 12604 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_137
timestamp 1688980957
transform 1 0 13708 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_149
timestamp 1688980957
transform 1 0 14812 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_161
timestamp 1688980957
transform 1 0 15916 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_167
timestamp 1688980957
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_169
timestamp 1688980957
transform 1 0 16652 0 -1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_210
timestamp 1688980957
transform 1 0 20424 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_222
timestamp 1688980957
transform 1 0 21528 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_225
timestamp 1688980957
transform 1 0 21804 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_236
timestamp 1688980957
transform 1 0 22816 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_250
timestamp 1688980957
transform 1 0 24104 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_262
timestamp 1688980957
transform 1 0 25208 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_278
timestamp 1688980957
transform 1 0 26680 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_297
timestamp 1688980957
transform 1 0 28428 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_301
timestamp 1688980957
transform 1 0 28796 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_313
timestamp 1688980957
transform 1 0 29900 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_321
timestamp 1688980957
transform 1 0 30636 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_332
timestamp 1688980957
transform 1 0 31648 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_353
timestamp 1688980957
transform 1 0 33580 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_361
timestamp 1688980957
transform 1 0 34316 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_3
timestamp 1688980957
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_15
timestamp 1688980957
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_27
timestamp 1688980957
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_29
timestamp 1688980957
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_41
timestamp 1688980957
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_53
timestamp 1688980957
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_65
timestamp 1688980957
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_77
timestamp 1688980957
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_83
timestamp 1688980957
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_85
timestamp 1688980957
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_97
timestamp 1688980957
transform 1 0 10028 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_109
timestamp 1688980957
transform 1 0 11132 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_121
timestamp 1688980957
transform 1 0 12236 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_133
timestamp 1688980957
transform 1 0 13340 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_139
timestamp 1688980957
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_141
timestamp 1688980957
transform 1 0 14076 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_153
timestamp 1688980957
transform 1 0 15180 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_165
timestamp 1688980957
transform 1 0 16284 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_177
timestamp 1688980957
transform 1 0 17388 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_181
timestamp 1688980957
transform 1 0 17756 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_186
timestamp 1688980957
transform 1 0 18216 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_194
timestamp 1688980957
transform 1 0 18952 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_197
timestamp 1688980957
transform 1 0 19228 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_205
timestamp 1688980957
transform 1 0 19964 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_212
timestamp 1688980957
transform 1 0 20608 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_224
timestamp 1688980957
transform 1 0 21712 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_228
timestamp 1688980957
transform 1 0 22080 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_240
timestamp 1688980957
transform 1 0 23184 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_244
timestamp 1688980957
transform 1 0 23552 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_266
timestamp 1688980957
transform 1 0 25576 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_274
timestamp 1688980957
transform 1 0 26312 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_309
timestamp 1688980957
transform 1 0 29532 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_313
timestamp 1688980957
transform 1 0 29900 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_319
timestamp 1688980957
transform 1 0 30452 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_336
timestamp 1688980957
transform 1 0 32016 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_340
timestamp 1688980957
transform 1 0 32384 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_357
timestamp 1688980957
transform 1 0 33948 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_363
timestamp 1688980957
transform 1 0 34500 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_3
timestamp 1688980957
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_15
timestamp 1688980957
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_27
timestamp 1688980957
transform 1 0 3588 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_39
timestamp 1688980957
transform 1 0 4692 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_51
timestamp 1688980957
transform 1 0 5796 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_55
timestamp 1688980957
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_57
timestamp 1688980957
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_69
timestamp 1688980957
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_81
timestamp 1688980957
transform 1 0 8556 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_93
timestamp 1688980957
transform 1 0 9660 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_105
timestamp 1688980957
transform 1 0 10764 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_111
timestamp 1688980957
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_113
timestamp 1688980957
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_125
timestamp 1688980957
transform 1 0 12604 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_137
timestamp 1688980957
transform 1 0 13708 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_149
timestamp 1688980957
transform 1 0 14812 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_161
timestamp 1688980957
transform 1 0 15916 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_167
timestamp 1688980957
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_169
timestamp 1688980957
transform 1 0 16652 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_181
timestamp 1688980957
transform 1 0 17756 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_194
timestamp 1688980957
transform 1 0 18952 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_273
timestamp 1688980957
transform 1 0 26220 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_279
timestamp 1688980957
transform 1 0 26772 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_329
timestamp 1688980957
transform 1 0 31372 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_335
timestamp 1688980957
transform 1 0 31924 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_354
timestamp 1688980957
transform 1 0 33672 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_362
timestamp 1688980957
transform 1 0 34408 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_3
timestamp 1688980957
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_15
timestamp 1688980957
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_27
timestamp 1688980957
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_29
timestamp 1688980957
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_41
timestamp 1688980957
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_53
timestamp 1688980957
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_65
timestamp 1688980957
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_77
timestamp 1688980957
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_83
timestamp 1688980957
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_85
timestamp 1688980957
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_97
timestamp 1688980957
transform 1 0 10028 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_109
timestamp 1688980957
transform 1 0 11132 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_121
timestamp 1688980957
transform 1 0 12236 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_133
timestamp 1688980957
transform 1 0 13340 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_139
timestamp 1688980957
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_141
timestamp 1688980957
transform 1 0 14076 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_153
timestamp 1688980957
transform 1 0 15180 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_165
timestamp 1688980957
transform 1 0 16284 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_189
timestamp 1688980957
transform 1 0 18492 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_197
timestamp 1688980957
transform 1 0 19228 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_201
timestamp 1688980957
transform 1 0 19596 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_218
timestamp 1688980957
transform 1 0 21160 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_240
timestamp 1688980957
transform 1 0 23184 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_246
timestamp 1688980957
transform 1 0 23736 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_251
timestamp 1688980957
transform 1 0 24196 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_280
timestamp 1688980957
transform 1 0 26864 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_286
timestamp 1688980957
transform 1 0 27416 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_297
timestamp 1688980957
transform 1 0 28428 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_305
timestamp 1688980957
transform 1 0 29164 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_309
timestamp 1688980957
transform 1 0 29532 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_316
timestamp 1688980957
transform 1 0 30176 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_330
timestamp 1688980957
transform 1 0 31464 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_356
timestamp 1688980957
transform 1 0 33856 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_360
timestamp 1688980957
transform 1 0 34224 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_3
timestamp 1688980957
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_15
timestamp 1688980957
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_27
timestamp 1688980957
transform 1 0 3588 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_39
timestamp 1688980957
transform 1 0 4692 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_51
timestamp 1688980957
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_55
timestamp 1688980957
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_57
timestamp 1688980957
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_69
timestamp 1688980957
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_81
timestamp 1688980957
transform 1 0 8556 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_93
timestamp 1688980957
transform 1 0 9660 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_105
timestamp 1688980957
transform 1 0 10764 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_111
timestamp 1688980957
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_113
timestamp 1688980957
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_125
timestamp 1688980957
transform 1 0 12604 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_137
timestamp 1688980957
transform 1 0 13708 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_149
timestamp 1688980957
transform 1 0 14812 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_161
timestamp 1688980957
transform 1 0 15916 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_167
timestamp 1688980957
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_169
timestamp 1688980957
transform 1 0 16652 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_188
timestamp 1688980957
transform 1 0 18400 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_198
timestamp 1688980957
transform 1 0 19320 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_210
timestamp 1688980957
transform 1 0 20424 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_218
timestamp 1688980957
transform 1 0 21160 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_233
timestamp 1688980957
transform 1 0 22540 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_239
timestamp 1688980957
transform 1 0 23092 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_244
timestamp 1688980957
transform 1 0 23552 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_250
timestamp 1688980957
transform 1 0 24104 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_262
timestamp 1688980957
transform 1 0 25208 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_271
timestamp 1688980957
transform 1 0 26036 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_277
timestamp 1688980957
transform 1 0 26588 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_281
timestamp 1688980957
transform 1 0 26956 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_304
timestamp 1688980957
transform 1 0 29072 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_314
timestamp 1688980957
transform 1 0 29992 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_318
timestamp 1688980957
transform 1 0 30360 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_335
timestamp 1688980957
transform 1 0 31924 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_337
timestamp 1688980957
transform 1 0 32108 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_347
timestamp 1688980957
transform 1 0 33028 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_359
timestamp 1688980957
transform 1 0 34132 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_363
timestamp 1688980957
transform 1 0 34500 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_3
timestamp 1688980957
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_15
timestamp 1688980957
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_27
timestamp 1688980957
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_29
timestamp 1688980957
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_41
timestamp 1688980957
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_53
timestamp 1688980957
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_65
timestamp 1688980957
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_77
timestamp 1688980957
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_83
timestamp 1688980957
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_85
timestamp 1688980957
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_97
timestamp 1688980957
transform 1 0 10028 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_109
timestamp 1688980957
transform 1 0 11132 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_121
timestamp 1688980957
transform 1 0 12236 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_133
timestamp 1688980957
transform 1 0 13340 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_139
timestamp 1688980957
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_141
timestamp 1688980957
transform 1 0 14076 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_153
timestamp 1688980957
transform 1 0 15180 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_165
timestamp 1688980957
transform 1 0 16284 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_173
timestamp 1688980957
transform 1 0 17020 0 1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_179
timestamp 1688980957
transform 1 0 17572 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_191
timestamp 1688980957
transform 1 0 18676 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_195
timestamp 1688980957
transform 1 0 19044 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_213
timestamp 1688980957
transform 1 0 20700 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_221
timestamp 1688980957
transform 1 0 21436 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_229
timestamp 1688980957
transform 1 0 22172 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_233
timestamp 1688980957
transform 1 0 22540 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_237
timestamp 1688980957
transform 1 0 22908 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_250
timestamp 1688980957
transform 1 0 24104 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_256
timestamp 1688980957
transform 1 0 24656 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_262
timestamp 1688980957
transform 1 0 25208 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_307
timestamp 1688980957
transform 1 0 29348 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_328
timestamp 1688980957
transform 1 0 31280 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_340
timestamp 1688980957
transform 1 0 32384 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_352
timestamp 1688980957
transform 1 0 33488 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_3
timestamp 1688980957
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_15
timestamp 1688980957
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_27
timestamp 1688980957
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_39
timestamp 1688980957
transform 1 0 4692 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_51
timestamp 1688980957
transform 1 0 5796 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_55
timestamp 1688980957
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_57
timestamp 1688980957
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_69
timestamp 1688980957
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_81
timestamp 1688980957
transform 1 0 8556 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_93
timestamp 1688980957
transform 1 0 9660 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_105
timestamp 1688980957
transform 1 0 10764 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_111
timestamp 1688980957
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_113
timestamp 1688980957
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_125
timestamp 1688980957
transform 1 0 12604 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_137
timestamp 1688980957
transform 1 0 13708 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_149
timestamp 1688980957
transform 1 0 14812 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_161
timestamp 1688980957
transform 1 0 15916 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_167
timestamp 1688980957
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_169
timestamp 1688980957
transform 1 0 16652 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_181
timestamp 1688980957
transform 1 0 17756 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_193
timestamp 1688980957
transform 1 0 18860 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_205
timestamp 1688980957
transform 1 0 19964 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_222
timestamp 1688980957
transform 1 0 21528 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_297
timestamp 1688980957
transform 1 0 28428 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_305
timestamp 1688980957
transform 1 0 29164 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_316
timestamp 1688980957
transform 1 0 30176 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_345
timestamp 1688980957
transform 1 0 32844 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_357
timestamp 1688980957
transform 1 0 33948 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_363
timestamp 1688980957
transform 1 0 34500 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_3
timestamp 1688980957
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_15
timestamp 1688980957
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_27
timestamp 1688980957
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_29
timestamp 1688980957
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_41
timestamp 1688980957
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_53
timestamp 1688980957
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_65
timestamp 1688980957
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_77
timestamp 1688980957
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_83
timestamp 1688980957
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_85
timestamp 1688980957
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_97
timestamp 1688980957
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_109
timestamp 1688980957
transform 1 0 11132 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_121
timestamp 1688980957
transform 1 0 12236 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_133
timestamp 1688980957
transform 1 0 13340 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_139
timestamp 1688980957
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_141
timestamp 1688980957
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_153
timestamp 1688980957
transform 1 0 15180 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_165
timestamp 1688980957
transform 1 0 16284 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_189
timestamp 1688980957
transform 1 0 18492 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_195
timestamp 1688980957
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_203
timestamp 1688980957
transform 1 0 19780 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_219
timestamp 1688980957
transform 1 0 21252 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_245
timestamp 1688980957
transform 1 0 23644 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_251
timestamp 1688980957
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_253
timestamp 1688980957
transform 1 0 24380 0 1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_272
timestamp 1688980957
transform 1 0 26128 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_284
timestamp 1688980957
transform 1 0 27232 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_296
timestamp 1688980957
transform 1 0 28336 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_307
timestamp 1688980957
transform 1 0 29348 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_309
timestamp 1688980957
transform 1 0 29532 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_316
timestamp 1688980957
transform 1 0 30176 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_331
timestamp 1688980957
transform 1 0 31556 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_351
timestamp 1688980957
transform 1 0 33396 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_363
timestamp 1688980957
transform 1 0 34500 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_3
timestamp 1688980957
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_15
timestamp 1688980957
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_27
timestamp 1688980957
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_39
timestamp 1688980957
transform 1 0 4692 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_51
timestamp 1688980957
transform 1 0 5796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_55
timestamp 1688980957
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_57
timestamp 1688980957
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_69
timestamp 1688980957
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_81
timestamp 1688980957
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_93
timestamp 1688980957
transform 1 0 9660 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_105
timestamp 1688980957
transform 1 0 10764 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_111
timestamp 1688980957
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_113
timestamp 1688980957
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_125
timestamp 1688980957
transform 1 0 12604 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_137
timestamp 1688980957
transform 1 0 13708 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_149
timestamp 1688980957
transform 1 0 14812 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_161
timestamp 1688980957
transform 1 0 15916 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_167
timestamp 1688980957
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_206
timestamp 1688980957
transform 1 0 20056 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_222
timestamp 1688980957
transform 1 0 21528 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_229
timestamp 1688980957
transform 1 0 22172 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_233
timestamp 1688980957
transform 1 0 22540 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_239
timestamp 1688980957
transform 1 0 23092 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_247
timestamp 1688980957
transform 1 0 23828 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_253
timestamp 1688980957
transform 1 0 24380 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_257
timestamp 1688980957
transform 1 0 24748 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_264
timestamp 1688980957
transform 1 0 25392 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_268
timestamp 1688980957
transform 1 0 25760 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_275
timestamp 1688980957
transform 1 0 26404 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_279
timestamp 1688980957
transform 1 0 26772 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_281
timestamp 1688980957
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_293
timestamp 1688980957
transform 1 0 28060 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_320
timestamp 1688980957
transform 1 0 30544 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_334
timestamp 1688980957
transform 1 0 31832 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_350
timestamp 1688980957
transform 1 0 33304 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_362
timestamp 1688980957
transform 1 0 34408 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_3
timestamp 1688980957
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_15
timestamp 1688980957
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_27
timestamp 1688980957
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_29
timestamp 1688980957
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_41
timestamp 1688980957
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_53
timestamp 1688980957
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_65
timestamp 1688980957
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_77
timestamp 1688980957
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_83
timestamp 1688980957
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_85
timestamp 1688980957
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_97
timestamp 1688980957
transform 1 0 10028 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_109
timestamp 1688980957
transform 1 0 11132 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_121
timestamp 1688980957
transform 1 0 12236 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_133
timestamp 1688980957
transform 1 0 13340 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_139
timestamp 1688980957
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_141
timestamp 1688980957
transform 1 0 14076 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_153
timestamp 1688980957
transform 1 0 15180 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_165
timestamp 1688980957
transform 1 0 16284 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_174
timestamp 1688980957
transform 1 0 17112 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_179
timestamp 1688980957
transform 1 0 17572 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_183
timestamp 1688980957
transform 1 0 17940 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_190
timestamp 1688980957
transform 1 0 18584 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_197
timestamp 1688980957
transform 1 0 19228 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_208
timestamp 1688980957
transform 1 0 20240 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_218
timestamp 1688980957
transform 1 0 21160 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_230
timestamp 1688980957
transform 1 0 22264 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_237
timestamp 1688980957
transform 1 0 22908 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_243
timestamp 1688980957
transform 1 0 23460 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_251
timestamp 1688980957
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_253
timestamp 1688980957
transform 1 0 24380 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_262
timestamp 1688980957
transform 1 0 25208 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_266
timestamp 1688980957
transform 1 0 25576 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_299
timestamp 1688980957
transform 1 0 28612 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_315
timestamp 1688980957
transform 1 0 30084 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_348
timestamp 1688980957
transform 1 0 33120 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_360
timestamp 1688980957
transform 1 0 34224 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_3
timestamp 1688980957
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_15
timestamp 1688980957
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_27
timestamp 1688980957
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_39
timestamp 1688980957
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_51
timestamp 1688980957
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_55
timestamp 1688980957
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_57
timestamp 1688980957
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_69
timestamp 1688980957
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_81
timestamp 1688980957
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_93
timestamp 1688980957
transform 1 0 9660 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_105
timestamp 1688980957
transform 1 0 10764 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_111
timestamp 1688980957
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_113
timestamp 1688980957
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_125
timestamp 1688980957
transform 1 0 12604 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_137
timestamp 1688980957
transform 1 0 13708 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_149
timestamp 1688980957
transform 1 0 14812 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_161
timestamp 1688980957
transform 1 0 15916 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_167
timestamp 1688980957
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_169
timestamp 1688980957
transform 1 0 16652 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_173
timestamp 1688980957
transform 1 0 17020 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_183
timestamp 1688980957
transform 1 0 17940 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_197
timestamp 1688980957
transform 1 0 19228 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_209
timestamp 1688980957
transform 1 0 20332 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_222
timestamp 1688980957
transform 1 0 21528 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_225
timestamp 1688980957
transform 1 0 21804 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_249
timestamp 1688980957
transform 1 0 24012 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_274
timestamp 1688980957
transform 1 0 26312 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_302
timestamp 1688980957
transform 1 0 28888 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_321
timestamp 1688980957
transform 1 0 30636 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_334
timestamp 1688980957
transform 1 0 31832 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_345
timestamp 1688980957
transform 1 0 32844 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_357
timestamp 1688980957
transform 1 0 33948 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_363
timestamp 1688980957
transform 1 0 34500 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_3
timestamp 1688980957
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_15
timestamp 1688980957
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_27
timestamp 1688980957
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_29
timestamp 1688980957
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_41
timestamp 1688980957
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_53
timestamp 1688980957
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_65
timestamp 1688980957
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_77
timestamp 1688980957
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_83
timestamp 1688980957
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_85
timestamp 1688980957
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_97
timestamp 1688980957
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_109
timestamp 1688980957
transform 1 0 11132 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_121
timestamp 1688980957
transform 1 0 12236 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_133
timestamp 1688980957
transform 1 0 13340 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_139
timestamp 1688980957
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_141
timestamp 1688980957
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_153
timestamp 1688980957
transform 1 0 15180 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_181
timestamp 1688980957
transform 1 0 17756 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_193
timestamp 1688980957
transform 1 0 18860 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_200
timestamp 1688980957
transform 1 0 19504 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_231
timestamp 1688980957
transform 1 0 22356 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_261
timestamp 1688980957
transform 1 0 25116 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_277
timestamp 1688980957
transform 1 0 26588 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_296
timestamp 1688980957
transform 1 0 28336 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_300
timestamp 1688980957
transform 1 0 28704 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_305
timestamp 1688980957
transform 1 0 29164 0 1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_315
timestamp 1688980957
transform 1 0 30084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_327
timestamp 1688980957
transform 1 0 31188 0 1 26112
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_351
timestamp 1688980957
transform 1 0 33396 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_363
timestamp 1688980957
transform 1 0 34500 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_3
timestamp 1688980957
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_15
timestamp 1688980957
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_27
timestamp 1688980957
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_39
timestamp 1688980957
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_51
timestamp 1688980957
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_55
timestamp 1688980957
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_57
timestamp 1688980957
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_69
timestamp 1688980957
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_81
timestamp 1688980957
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_93
timestamp 1688980957
transform 1 0 9660 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_105
timestamp 1688980957
transform 1 0 10764 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_111
timestamp 1688980957
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_113
timestamp 1688980957
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_125
timestamp 1688980957
transform 1 0 12604 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_137
timestamp 1688980957
transform 1 0 13708 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_149
timestamp 1688980957
transform 1 0 14812 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_161
timestamp 1688980957
transform 1 0 15916 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_167
timestamp 1688980957
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_169
timestamp 1688980957
transform 1 0 16652 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_175
timestamp 1688980957
transform 1 0 17204 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_221
timestamp 1688980957
transform 1 0 21436 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_248
timestamp 1688980957
transform 1 0 23920 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_256
timestamp 1688980957
transform 1 0 24656 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_261
timestamp 1688980957
transform 1 0 25116 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_270
timestamp 1688980957
transform 1 0 25944 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_278
timestamp 1688980957
transform 1 0 26680 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_281
timestamp 1688980957
transform 1 0 26956 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_293
timestamp 1688980957
transform 1 0 28060 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_299
timestamp 1688980957
transform 1 0 28612 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_308
timestamp 1688980957
transform 1 0 29440 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_320
timestamp 1688980957
transform 1 0 30544 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_328
timestamp 1688980957
transform 1 0 31280 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_337
timestamp 1688980957
transform 1 0 32108 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_342
timestamp 1688980957
transform 1 0 32568 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_354
timestamp 1688980957
transform 1 0 33672 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_362
timestamp 1688980957
transform 1 0 34408 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_3
timestamp 1688980957
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_15
timestamp 1688980957
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_27
timestamp 1688980957
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_29
timestamp 1688980957
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_41
timestamp 1688980957
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_53
timestamp 1688980957
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_65
timestamp 1688980957
transform 1 0 7084 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_77
timestamp 1688980957
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_83
timestamp 1688980957
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_85
timestamp 1688980957
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_97
timestamp 1688980957
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_109
timestamp 1688980957
transform 1 0 11132 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_121
timestamp 1688980957
transform 1 0 12236 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_133
timestamp 1688980957
transform 1 0 13340 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_139
timestamp 1688980957
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_141
timestamp 1688980957
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_153
timestamp 1688980957
transform 1 0 15180 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_165
timestamp 1688980957
transform 1 0 16284 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_188
timestamp 1688980957
transform 1 0 18400 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_192
timestamp 1688980957
transform 1 0 18768 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_197
timestamp 1688980957
transform 1 0 19228 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_217
timestamp 1688980957
transform 1 0 21068 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_229
timestamp 1688980957
transform 1 0 22172 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_243
timestamp 1688980957
transform 1 0 23460 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_269
timestamp 1688980957
transform 1 0 25852 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_278
timestamp 1688980957
transform 1 0 26680 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_298
timestamp 1688980957
transform 1 0 28520 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_341
timestamp 1688980957
transform 1 0 32476 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_353
timestamp 1688980957
transform 1 0 33580 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_361
timestamp 1688980957
transform 1 0 34316 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_3
timestamp 1688980957
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_15
timestamp 1688980957
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_27
timestamp 1688980957
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_39
timestamp 1688980957
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_51
timestamp 1688980957
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_55
timestamp 1688980957
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_57
timestamp 1688980957
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_69
timestamp 1688980957
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_81
timestamp 1688980957
transform 1 0 8556 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_93
timestamp 1688980957
transform 1 0 9660 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_105
timestamp 1688980957
transform 1 0 10764 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_111
timestamp 1688980957
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_113
timestamp 1688980957
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_125
timestamp 1688980957
transform 1 0 12604 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_137
timestamp 1688980957
transform 1 0 13708 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_149
timestamp 1688980957
transform 1 0 14812 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_161
timestamp 1688980957
transform 1 0 15916 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_167
timestamp 1688980957
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_169
timestamp 1688980957
transform 1 0 16652 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_185
timestamp 1688980957
transform 1 0 18124 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_191
timestamp 1688980957
transform 1 0 18676 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_195
timestamp 1688980957
transform 1 0 19044 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_203
timestamp 1688980957
transform 1 0 19780 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_215
timestamp 1688980957
transform 1 0 20884 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_223
timestamp 1688980957
transform 1 0 21620 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_225
timestamp 1688980957
transform 1 0 21804 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_229
timestamp 1688980957
transform 1 0 22172 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_262
timestamp 1688980957
transform 1 0 25208 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_308
timestamp 1688980957
transform 1 0 29440 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_316
timestamp 1688980957
transform 1 0 30176 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_329
timestamp 1688980957
transform 1 0 31372 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_344
timestamp 1688980957
transform 1 0 32752 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_356
timestamp 1688980957
transform 1 0 33856 0 -1 28288
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_3
timestamp 1688980957
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_15
timestamp 1688980957
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_27
timestamp 1688980957
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_29
timestamp 1688980957
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_41
timestamp 1688980957
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_53
timestamp 1688980957
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_65
timestamp 1688980957
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_77
timestamp 1688980957
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_83
timestamp 1688980957
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_85
timestamp 1688980957
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_97
timestamp 1688980957
transform 1 0 10028 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_109
timestamp 1688980957
transform 1 0 11132 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_121
timestamp 1688980957
transform 1 0 12236 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_133
timestamp 1688980957
transform 1 0 13340 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_139
timestamp 1688980957
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_141
timestamp 1688980957
transform 1 0 14076 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_153
timestamp 1688980957
transform 1 0 15180 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_48_193
timestamp 1688980957
transform 1 0 18860 0 1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_197
timestamp 1688980957
transform 1 0 19228 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_209
timestamp 1688980957
transform 1 0 20332 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_48_235
timestamp 1688980957
transform 1 0 22724 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_241
timestamp 1688980957
transform 1 0 23276 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_250
timestamp 1688980957
transform 1 0 24104 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_48_253
timestamp 1688980957
transform 1 0 24380 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_259
timestamp 1688980957
transform 1 0 24932 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_270
timestamp 1688980957
transform 1 0 25944 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_282
timestamp 1688980957
transform 1 0 27048 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_288
timestamp 1688980957
transform 1 0 27600 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_294
timestamp 1688980957
transform 1 0 28152 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_306
timestamp 1688980957
transform 1 0 29256 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_309
timestamp 1688980957
transform 1 0 29532 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_313
timestamp 1688980957
transform 1 0 29900 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_330
timestamp 1688980957
transform 1 0 31464 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_347
timestamp 1688980957
transform 1 0 33028 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_359
timestamp 1688980957
transform 1 0 34132 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_363
timestamp 1688980957
transform 1 0 34500 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_3
timestamp 1688980957
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_15
timestamp 1688980957
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_27
timestamp 1688980957
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_39
timestamp 1688980957
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_51
timestamp 1688980957
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_55
timestamp 1688980957
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_57
timestamp 1688980957
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_69
timestamp 1688980957
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_81
timestamp 1688980957
transform 1 0 8556 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_93
timestamp 1688980957
transform 1 0 9660 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_105
timestamp 1688980957
transform 1 0 10764 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_111
timestamp 1688980957
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_113
timestamp 1688980957
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_125
timestamp 1688980957
transform 1 0 12604 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_137
timestamp 1688980957
transform 1 0 13708 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_149
timestamp 1688980957
transform 1 0 14812 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_161
timestamp 1688980957
transform 1 0 15916 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_167
timestamp 1688980957
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_169
timestamp 1688980957
transform 1 0 16652 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_176
timestamp 1688980957
transform 1 0 17296 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_188
timestamp 1688980957
transform 1 0 18400 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_197
timestamp 1688980957
transform 1 0 19228 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_228
timestamp 1688980957
transform 1 0 22080 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_236
timestamp 1688980957
transform 1 0 22816 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_240
timestamp 1688980957
transform 1 0 23184 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_252
timestamp 1688980957
transform 1 0 24288 0 -1 29376
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_263
timestamp 1688980957
transform 1 0 25300 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_275
timestamp 1688980957
transform 1 0 26404 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_279
timestamp 1688980957
transform 1 0 26772 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_281
timestamp 1688980957
transform 1 0 26956 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_293
timestamp 1688980957
transform 1 0 28060 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_303
timestamp 1688980957
transform 1 0 28980 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_315
timestamp 1688980957
transform 1 0 30084 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_327
timestamp 1688980957
transform 1 0 31188 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_334
timestamp 1688980957
transform 1 0 31832 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_342
timestamp 1688980957
transform 1 0 32568 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_354
timestamp 1688980957
transform 1 0 33672 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_362
timestamp 1688980957
transform 1 0 34408 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_3
timestamp 1688980957
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_15
timestamp 1688980957
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_27
timestamp 1688980957
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_29
timestamp 1688980957
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_41
timestamp 1688980957
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_53
timestamp 1688980957
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_65
timestamp 1688980957
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_77
timestamp 1688980957
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_83
timestamp 1688980957
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_85
timestamp 1688980957
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_97
timestamp 1688980957
transform 1 0 10028 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_109
timestamp 1688980957
transform 1 0 11132 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_121
timestamp 1688980957
transform 1 0 12236 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_133
timestamp 1688980957
transform 1 0 13340 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_139
timestamp 1688980957
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_141
timestamp 1688980957
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_153
timestamp 1688980957
transform 1 0 15180 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_165
timestamp 1688980957
transform 1 0 16284 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_180
timestamp 1688980957
transform 1 0 17664 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_184
timestamp 1688980957
transform 1 0 18032 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_194
timestamp 1688980957
transform 1 0 18952 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_204
timestamp 1688980957
transform 1 0 19872 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_223
timestamp 1688980957
transform 1 0 21620 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_50_231
timestamp 1688980957
transform 1 0 22356 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_240
timestamp 1688980957
transform 1 0 23184 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_253
timestamp 1688980957
transform 1 0 24380 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_257
timestamp 1688980957
transform 1 0 24748 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_269
timestamp 1688980957
transform 1 0 25852 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_290
timestamp 1688980957
transform 1 0 27784 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_50_325
timestamp 1688980957
transform 1 0 31004 0 1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_344
timestamp 1688980957
transform 1 0 32752 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_356
timestamp 1688980957
transform 1 0 33856 0 1 29376
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_9
timestamp 1688980957
transform 1 0 1932 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_21
timestamp 1688980957
transform 1 0 3036 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_33
timestamp 1688980957
transform 1 0 4140 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_45
timestamp 1688980957
transform 1 0 5244 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_51_53
timestamp 1688980957
transform 1 0 5980 0 -1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_57
timestamp 1688980957
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_69
timestamp 1688980957
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_81
timestamp 1688980957
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_93
timestamp 1688980957
transform 1 0 9660 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_105
timestamp 1688980957
transform 1 0 10764 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_111
timestamp 1688980957
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_113
timestamp 1688980957
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_125
timestamp 1688980957
transform 1 0 12604 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_137
timestamp 1688980957
transform 1 0 13708 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_149
timestamp 1688980957
transform 1 0 14812 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_161
timestamp 1688980957
transform 1 0 15916 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_185
timestamp 1688980957
transform 1 0 18124 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_198
timestamp 1688980957
transform 1 0 19320 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_206
timestamp 1688980957
transform 1 0 20056 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_222
timestamp 1688980957
transform 1 0 21528 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_260
timestamp 1688980957
transform 1 0 25024 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_279
timestamp 1688980957
transform 1 0 26772 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_302
timestamp 1688980957
transform 1 0 28888 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_310
timestamp 1688980957
transform 1 0 29624 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_325
timestamp 1688980957
transform 1 0 31004 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_330
timestamp 1688980957
transform 1 0 31464 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_335
timestamp 1688980957
transform 1 0 31924 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_337
timestamp 1688980957
transform 1 0 32108 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_349
timestamp 1688980957
transform 1 0 33212 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_51_361
timestamp 1688980957
transform 1 0 34316 0 -1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_3
timestamp 1688980957
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_15
timestamp 1688980957
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_27
timestamp 1688980957
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_29
timestamp 1688980957
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_41
timestamp 1688980957
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_53
timestamp 1688980957
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_65
timestamp 1688980957
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_77
timestamp 1688980957
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_83
timestamp 1688980957
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_85
timestamp 1688980957
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_97
timestamp 1688980957
transform 1 0 10028 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_109
timestamp 1688980957
transform 1 0 11132 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_121
timestamp 1688980957
transform 1 0 12236 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_133
timestamp 1688980957
transform 1 0 13340 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_139
timestamp 1688980957
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_141
timestamp 1688980957
transform 1 0 14076 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_153
timestamp 1688980957
transform 1 0 15180 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52_165
timestamp 1688980957
transform 1 0 16284 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_169
timestamp 1688980957
transform 1 0 16652 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_176
timestamp 1688980957
transform 1 0 17296 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_185
timestamp 1688980957
transform 1 0 18124 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_206
timestamp 1688980957
transform 1 0 20056 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_52_218
timestamp 1688980957
transform 1 0 21160 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_226
timestamp 1688980957
transform 1 0 21896 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_251
timestamp 1688980957
transform 1 0 24196 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_257
timestamp 1688980957
transform 1 0 24748 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_274
timestamp 1688980957
transform 1 0 26312 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_282
timestamp 1688980957
transform 1 0 27048 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52_303
timestamp 1688980957
transform 1 0 28980 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_307
timestamp 1688980957
transform 1 0 29348 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_344
timestamp 1688980957
transform 1 0 32752 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_52_356
timestamp 1688980957
transform 1 0 33856 0 1 30464
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_3
timestamp 1688980957
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_15
timestamp 1688980957
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_27
timestamp 1688980957
transform 1 0 3588 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_39
timestamp 1688980957
transform 1 0 4692 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_51
timestamp 1688980957
transform 1 0 5796 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_55
timestamp 1688980957
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_57
timestamp 1688980957
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_69
timestamp 1688980957
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_81
timestamp 1688980957
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_93
timestamp 1688980957
transform 1 0 9660 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_105
timestamp 1688980957
transform 1 0 10764 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_111
timestamp 1688980957
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_113
timestamp 1688980957
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_125
timestamp 1688980957
transform 1 0 12604 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_137
timestamp 1688980957
transform 1 0 13708 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_149
timestamp 1688980957
transform 1 0 14812 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_161
timestamp 1688980957
transform 1 0 15916 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_167
timestamp 1688980957
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_53_189
timestamp 1688980957
transform 1 0 18492 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53_222
timestamp 1688980957
transform 1 0 21528 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_225
timestamp 1688980957
transform 1 0 21804 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_237
timestamp 1688980957
transform 1 0 22908 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_267
timestamp 1688980957
transform 1 0 25668 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_279
timestamp 1688980957
transform 1 0 26772 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_53_281
timestamp 1688980957
transform 1 0 26956 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53_289
timestamp 1688980957
transform 1 0 27692 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_294
timestamp 1688980957
transform 1 0 28152 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_306
timestamp 1688980957
transform 1 0 29256 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_310
timestamp 1688980957
transform 1 0 29624 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_314
timestamp 1688980957
transform 1 0 29992 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_53_353
timestamp 1688980957
transform 1 0 33580 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53_361
timestamp 1688980957
transform 1 0 34316 0 -1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_3
timestamp 1688980957
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_15
timestamp 1688980957
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_27
timestamp 1688980957
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_29
timestamp 1688980957
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_41
timestamp 1688980957
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_53
timestamp 1688980957
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_65
timestamp 1688980957
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_77
timestamp 1688980957
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_83
timestamp 1688980957
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_85
timestamp 1688980957
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_97
timestamp 1688980957
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_109
timestamp 1688980957
transform 1 0 11132 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_121
timestamp 1688980957
transform 1 0 12236 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_133
timestamp 1688980957
transform 1 0 13340 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_139
timestamp 1688980957
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_141
timestamp 1688980957
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_153
timestamp 1688980957
transform 1 0 15180 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_54_165
timestamp 1688980957
transform 1 0 16284 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_54_189
timestamp 1688980957
transform 1 0 18492 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_195
timestamp 1688980957
transform 1 0 19044 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_197
timestamp 1688980957
transform 1 0 19228 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_228
timestamp 1688980957
transform 1 0 22080 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_240
timestamp 1688980957
transform 1 0 23184 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_253
timestamp 1688980957
transform 1 0 24380 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_54_265
timestamp 1688980957
transform 1 0 25484 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_269
timestamp 1688980957
transform 1 0 25852 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_275
timestamp 1688980957
transform 1 0 26404 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_287
timestamp 1688980957
transform 1 0 27508 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_299
timestamp 1688980957
transform 1 0 28612 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_54_305
timestamp 1688980957
transform 1 0 29164 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_54_309
timestamp 1688980957
transform 1 0 29532 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_327
timestamp 1688980957
transform 1 0 31188 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_339
timestamp 1688980957
transform 1 0 32292 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_351
timestamp 1688980957
transform 1 0 33396 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_363
timestamp 1688980957
transform 1 0 34500 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_3
timestamp 1688980957
transform 1 0 1380 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_15
timestamp 1688980957
transform 1 0 2484 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_27
timestamp 1688980957
transform 1 0 3588 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_39
timestamp 1688980957
transform 1 0 4692 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_55_51
timestamp 1688980957
transform 1 0 5796 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_55
timestamp 1688980957
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_57
timestamp 1688980957
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_69
timestamp 1688980957
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_81
timestamp 1688980957
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_93
timestamp 1688980957
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_105
timestamp 1688980957
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_111
timestamp 1688980957
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_113
timestamp 1688980957
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_125
timestamp 1688980957
transform 1 0 12604 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_137
timestamp 1688980957
transform 1 0 13708 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_149
timestamp 1688980957
transform 1 0 14812 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_161
timestamp 1688980957
transform 1 0 15916 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_167
timestamp 1688980957
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_55_169
timestamp 1688980957
transform 1 0 16652 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_55_183
timestamp 1688980957
transform 1 0 17940 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_187
timestamp 1688980957
transform 1 0 18308 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_55_204
timestamp 1688980957
transform 1 0 19872 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_55_211
timestamp 1688980957
transform 1 0 20516 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_55_219
timestamp 1688980957
transform 1 0 21252 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_223
timestamp 1688980957
transform 1 0 21620 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_55_241
timestamp 1688980957
transform 1 0 23276 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_55_249
timestamp 1688980957
transform 1 0 24012 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_55_289
timestamp 1688980957
transform 1 0 27692 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_55_308
timestamp 1688980957
transform 1 0 29440 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_318
timestamp 1688980957
transform 1 0 30360 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_335
timestamp 1688980957
transform 1 0 31924 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_337
timestamp 1688980957
transform 1 0 32108 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_349
timestamp 1688980957
transform 1 0 33212 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_3
timestamp 1688980957
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_15
timestamp 1688980957
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_27
timestamp 1688980957
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_29
timestamp 1688980957
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_41
timestamp 1688980957
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_53
timestamp 1688980957
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_65
timestamp 1688980957
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_77
timestamp 1688980957
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_83
timestamp 1688980957
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_85
timestamp 1688980957
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_97
timestamp 1688980957
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_109
timestamp 1688980957
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_121
timestamp 1688980957
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_133
timestamp 1688980957
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_139
timestamp 1688980957
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_141
timestamp 1688980957
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_153
timestamp 1688980957
transform 1 0 15180 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_165
timestamp 1688980957
transform 1 0 16284 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_177
timestamp 1688980957
transform 1 0 17388 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_189
timestamp 1688980957
transform 1 0 18492 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_195
timestamp 1688980957
transform 1 0 19044 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_197
timestamp 1688980957
transform 1 0 19228 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_209
timestamp 1688980957
transform 1 0 20332 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_221
timestamp 1688980957
transform 1 0 21436 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_56_233
timestamp 1688980957
transform 1 0 22540 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_56_241
timestamp 1688980957
transform 1 0 23276 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_283
timestamp 1688980957
transform 1 0 27140 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_331
timestamp 1688980957
transform 1 0 31556 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_343
timestamp 1688980957
transform 1 0 32660 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_56_355
timestamp 1688980957
transform 1 0 33764 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_363
timestamp 1688980957
transform 1 0 34500 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_3
timestamp 1688980957
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_15
timestamp 1688980957
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_27
timestamp 1688980957
transform 1 0 3588 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_39
timestamp 1688980957
transform 1 0 4692 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57_51
timestamp 1688980957
transform 1 0 5796 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_55
timestamp 1688980957
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_57
timestamp 1688980957
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_69
timestamp 1688980957
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_81
timestamp 1688980957
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_93
timestamp 1688980957
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_105
timestamp 1688980957
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_111
timestamp 1688980957
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_113
timestamp 1688980957
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_125
timestamp 1688980957
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_137
timestamp 1688980957
transform 1 0 13708 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_149
timestamp 1688980957
transform 1 0 14812 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_161
timestamp 1688980957
transform 1 0 15916 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_167
timestamp 1688980957
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_169
timestamp 1688980957
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_181
timestamp 1688980957
transform 1 0 17756 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_193
timestamp 1688980957
transform 1 0 18860 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_205
timestamp 1688980957
transform 1 0 19964 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_217
timestamp 1688980957
transform 1 0 21068 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_223
timestamp 1688980957
transform 1 0 21620 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_225
timestamp 1688980957
transform 1 0 21804 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_242
timestamp 1688980957
transform 1 0 23368 0 -1 33728
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_251
timestamp 1688980957
transform 1 0 24196 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57_263
timestamp 1688980957
transform 1 0 25300 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57_286
timestamp 1688980957
transform 1 0 27416 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57_294
timestamp 1688980957
transform 1 0 28152 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57_326
timestamp 1688980957
transform 1 0 31096 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57_334
timestamp 1688980957
transform 1 0 31832 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_337
timestamp 1688980957
transform 1 0 32108 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_349
timestamp 1688980957
transform 1 0 33212 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_57_361
timestamp 1688980957
transform 1 0 34316 0 -1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_3
timestamp 1688980957
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_15
timestamp 1688980957
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_27
timestamp 1688980957
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_29
timestamp 1688980957
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_41
timestamp 1688980957
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_53
timestamp 1688980957
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_65
timestamp 1688980957
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_77
timestamp 1688980957
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_83
timestamp 1688980957
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_85
timestamp 1688980957
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_97
timestamp 1688980957
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_109
timestamp 1688980957
transform 1 0 11132 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_121
timestamp 1688980957
transform 1 0 12236 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_133
timestamp 1688980957
transform 1 0 13340 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_139
timestamp 1688980957
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_141
timestamp 1688980957
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_153
timestamp 1688980957
transform 1 0 15180 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_165
timestamp 1688980957
transform 1 0 16284 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_177
timestamp 1688980957
transform 1 0 17388 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_189
timestamp 1688980957
transform 1 0 18492 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_195
timestamp 1688980957
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_197
timestamp 1688980957
transform 1 0 19228 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_209
timestamp 1688980957
transform 1 0 20332 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_221
timestamp 1688980957
transform 1 0 21436 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_233
timestamp 1688980957
transform 1 0 22540 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_245
timestamp 1688980957
transform 1 0 23644 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_251
timestamp 1688980957
transform 1 0 24196 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_253
timestamp 1688980957
transform 1 0 24380 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_58_265
timestamp 1688980957
transform 1 0 25484 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_273
timestamp 1688980957
transform 1 0 26220 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_277
timestamp 1688980957
transform 1 0 26588 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_289
timestamp 1688980957
transform 1 0 27692 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_301
timestamp 1688980957
transform 1 0 28796 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_307
timestamp 1688980957
transform 1 0 29348 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_309
timestamp 1688980957
transform 1 0 29532 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_321
timestamp 1688980957
transform 1 0 30636 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_333
timestamp 1688980957
transform 1 0 31740 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_345
timestamp 1688980957
transform 1 0 32844 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_357
timestamp 1688980957
transform 1 0 33948 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_363
timestamp 1688980957
transform 1 0 34500 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_3
timestamp 1688980957
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_15
timestamp 1688980957
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_27
timestamp 1688980957
transform 1 0 3588 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_39
timestamp 1688980957
transform 1 0 4692 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_59_51
timestamp 1688980957
transform 1 0 5796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_55
timestamp 1688980957
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_57
timestamp 1688980957
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_69
timestamp 1688980957
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_81
timestamp 1688980957
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_93
timestamp 1688980957
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_105
timestamp 1688980957
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_111
timestamp 1688980957
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_113
timestamp 1688980957
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_125
timestamp 1688980957
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_137
timestamp 1688980957
transform 1 0 13708 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_149
timestamp 1688980957
transform 1 0 14812 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_161
timestamp 1688980957
transform 1 0 15916 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_167
timestamp 1688980957
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_169
timestamp 1688980957
transform 1 0 16652 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_181
timestamp 1688980957
transform 1 0 17756 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_193
timestamp 1688980957
transform 1 0 18860 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_205
timestamp 1688980957
transform 1 0 19964 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_217
timestamp 1688980957
transform 1 0 21068 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_223
timestamp 1688980957
transform 1 0 21620 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_225
timestamp 1688980957
transform 1 0 21804 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_237
timestamp 1688980957
transform 1 0 22908 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_249
timestamp 1688980957
transform 1 0 24012 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_261
timestamp 1688980957
transform 1 0 25116 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_273
timestamp 1688980957
transform 1 0 26220 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_279
timestamp 1688980957
transform 1 0 26772 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_281
timestamp 1688980957
transform 1 0 26956 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_293
timestamp 1688980957
transform 1 0 28060 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_305
timestamp 1688980957
transform 1 0 29164 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_317
timestamp 1688980957
transform 1 0 30268 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_329
timestamp 1688980957
transform 1 0 31372 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_335
timestamp 1688980957
transform 1 0 31924 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_337
timestamp 1688980957
transform 1 0 32108 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_349
timestamp 1688980957
transform 1 0 33212 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_59_361
timestamp 1688980957
transform 1 0 34316 0 -1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_3
timestamp 1688980957
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_15
timestamp 1688980957
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_27
timestamp 1688980957
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_29
timestamp 1688980957
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_41
timestamp 1688980957
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_53
timestamp 1688980957
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_65
timestamp 1688980957
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_77
timestamp 1688980957
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_83
timestamp 1688980957
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_85
timestamp 1688980957
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_97
timestamp 1688980957
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_109
timestamp 1688980957
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_121
timestamp 1688980957
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_133
timestamp 1688980957
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_139
timestamp 1688980957
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_141
timestamp 1688980957
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_153
timestamp 1688980957
transform 1 0 15180 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_165
timestamp 1688980957
transform 1 0 16284 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_177
timestamp 1688980957
transform 1 0 17388 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_189
timestamp 1688980957
transform 1 0 18492 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_195
timestamp 1688980957
transform 1 0 19044 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_197
timestamp 1688980957
transform 1 0 19228 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_209
timestamp 1688980957
transform 1 0 20332 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_221
timestamp 1688980957
transform 1 0 21436 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_233
timestamp 1688980957
transform 1 0 22540 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_245
timestamp 1688980957
transform 1 0 23644 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_251
timestamp 1688980957
transform 1 0 24196 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_253
timestamp 1688980957
transform 1 0 24380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_265
timestamp 1688980957
transform 1 0 25484 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_277
timestamp 1688980957
transform 1 0 26588 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_289
timestamp 1688980957
transform 1 0 27692 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_301
timestamp 1688980957
transform 1 0 28796 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_307
timestamp 1688980957
transform 1 0 29348 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_309
timestamp 1688980957
transform 1 0 29532 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_321
timestamp 1688980957
transform 1 0 30636 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_333
timestamp 1688980957
transform 1 0 31740 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_345
timestamp 1688980957
transform 1 0 32844 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_357
timestamp 1688980957
transform 1 0 33948 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_363
timestamp 1688980957
transform 1 0 34500 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_3
timestamp 1688980957
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_15
timestamp 1688980957
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_27
timestamp 1688980957
transform 1 0 3588 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_39
timestamp 1688980957
transform 1 0 4692 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_61_51
timestamp 1688980957
transform 1 0 5796 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_55
timestamp 1688980957
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_57
timestamp 1688980957
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_69
timestamp 1688980957
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_81
timestamp 1688980957
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_93
timestamp 1688980957
transform 1 0 9660 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_105
timestamp 1688980957
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_111
timestamp 1688980957
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_113
timestamp 1688980957
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_125
timestamp 1688980957
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_137
timestamp 1688980957
transform 1 0 13708 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_149
timestamp 1688980957
transform 1 0 14812 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_161
timestamp 1688980957
transform 1 0 15916 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_167
timestamp 1688980957
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_169
timestamp 1688980957
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_181
timestamp 1688980957
transform 1 0 17756 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_193
timestamp 1688980957
transform 1 0 18860 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_205
timestamp 1688980957
transform 1 0 19964 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_217
timestamp 1688980957
transform 1 0 21068 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_223
timestamp 1688980957
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_225
timestamp 1688980957
transform 1 0 21804 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_237
timestamp 1688980957
transform 1 0 22908 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_249
timestamp 1688980957
transform 1 0 24012 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_261
timestamp 1688980957
transform 1 0 25116 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_273
timestamp 1688980957
transform 1 0 26220 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_279
timestamp 1688980957
transform 1 0 26772 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_281
timestamp 1688980957
transform 1 0 26956 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_293
timestamp 1688980957
transform 1 0 28060 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_305
timestamp 1688980957
transform 1 0 29164 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_317
timestamp 1688980957
transform 1 0 30268 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_329
timestamp 1688980957
transform 1 0 31372 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_335
timestamp 1688980957
transform 1 0 31924 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_337
timestamp 1688980957
transform 1 0 32108 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_349
timestamp 1688980957
transform 1 0 33212 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_61_361
timestamp 1688980957
transform 1 0 34316 0 -1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_3
timestamp 1688980957
transform 1 0 1380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_15
timestamp 1688980957
transform 1 0 2484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_27
timestamp 1688980957
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_29
timestamp 1688980957
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_41
timestamp 1688980957
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_53
timestamp 1688980957
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_65
timestamp 1688980957
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_77
timestamp 1688980957
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_83
timestamp 1688980957
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_85
timestamp 1688980957
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_97
timestamp 1688980957
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_109
timestamp 1688980957
transform 1 0 11132 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_121
timestamp 1688980957
transform 1 0 12236 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_133
timestamp 1688980957
transform 1 0 13340 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_139
timestamp 1688980957
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_141
timestamp 1688980957
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_153
timestamp 1688980957
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_165
timestamp 1688980957
transform 1 0 16284 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_177
timestamp 1688980957
transform 1 0 17388 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_189
timestamp 1688980957
transform 1 0 18492 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_195
timestamp 1688980957
transform 1 0 19044 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_197
timestamp 1688980957
transform 1 0 19228 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_209
timestamp 1688980957
transform 1 0 20332 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_221
timestamp 1688980957
transform 1 0 21436 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_233
timestamp 1688980957
transform 1 0 22540 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_245
timestamp 1688980957
transform 1 0 23644 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_251
timestamp 1688980957
transform 1 0 24196 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_253
timestamp 1688980957
transform 1 0 24380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_265
timestamp 1688980957
transform 1 0 25484 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_277
timestamp 1688980957
transform 1 0 26588 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_289
timestamp 1688980957
transform 1 0 27692 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_301
timestamp 1688980957
transform 1 0 28796 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_307
timestamp 1688980957
transform 1 0 29348 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_309
timestamp 1688980957
transform 1 0 29532 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_321
timestamp 1688980957
transform 1 0 30636 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_333
timestamp 1688980957
transform 1 0 31740 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_345
timestamp 1688980957
transform 1 0 32844 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_357
timestamp 1688980957
transform 1 0 33948 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_363
timestamp 1688980957
transform 1 0 34500 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_3
timestamp 1688980957
transform 1 0 1380 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_15
timestamp 1688980957
transform 1 0 2484 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_27
timestamp 1688980957
transform 1 0 3588 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_39
timestamp 1688980957
transform 1 0 4692 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_63_51
timestamp 1688980957
transform 1 0 5796 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_55
timestamp 1688980957
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_57
timestamp 1688980957
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_69
timestamp 1688980957
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_81
timestamp 1688980957
transform 1 0 8556 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_93
timestamp 1688980957
transform 1 0 9660 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_105
timestamp 1688980957
transform 1 0 10764 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_111
timestamp 1688980957
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_113
timestamp 1688980957
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_125
timestamp 1688980957
transform 1 0 12604 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_137
timestamp 1688980957
transform 1 0 13708 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_149
timestamp 1688980957
transform 1 0 14812 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_161
timestamp 1688980957
transform 1 0 15916 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_167
timestamp 1688980957
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_169
timestamp 1688980957
transform 1 0 16652 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_181
timestamp 1688980957
transform 1 0 17756 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_193
timestamp 1688980957
transform 1 0 18860 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_205
timestamp 1688980957
transform 1 0 19964 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_217
timestamp 1688980957
transform 1 0 21068 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_223
timestamp 1688980957
transform 1 0 21620 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_225
timestamp 1688980957
transform 1 0 21804 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_237
timestamp 1688980957
transform 1 0 22908 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_249
timestamp 1688980957
transform 1 0 24012 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_261
timestamp 1688980957
transform 1 0 25116 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_273
timestamp 1688980957
transform 1 0 26220 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_279
timestamp 1688980957
transform 1 0 26772 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_281
timestamp 1688980957
transform 1 0 26956 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_293
timestamp 1688980957
transform 1 0 28060 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_305
timestamp 1688980957
transform 1 0 29164 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_317
timestamp 1688980957
transform 1 0 30268 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_329
timestamp 1688980957
transform 1 0 31372 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_335
timestamp 1688980957
transform 1 0 31924 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_337
timestamp 1688980957
transform 1 0 32108 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_349
timestamp 1688980957
transform 1 0 33212 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_63_361
timestamp 1688980957
transform 1 0 34316 0 -1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_3
timestamp 1688980957
transform 1 0 1380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_15
timestamp 1688980957
transform 1 0 2484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_27
timestamp 1688980957
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_29
timestamp 1688980957
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_41
timestamp 1688980957
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_53
timestamp 1688980957
transform 1 0 5980 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_65
timestamp 1688980957
transform 1 0 7084 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_77
timestamp 1688980957
transform 1 0 8188 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_83
timestamp 1688980957
transform 1 0 8740 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_85
timestamp 1688980957
transform 1 0 8924 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_97
timestamp 1688980957
transform 1 0 10028 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_109
timestamp 1688980957
transform 1 0 11132 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_121
timestamp 1688980957
transform 1 0 12236 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_133
timestamp 1688980957
transform 1 0 13340 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_139
timestamp 1688980957
transform 1 0 13892 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_141
timestamp 1688980957
transform 1 0 14076 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_153
timestamp 1688980957
transform 1 0 15180 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_165
timestamp 1688980957
transform 1 0 16284 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_177
timestamp 1688980957
transform 1 0 17388 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_189
timestamp 1688980957
transform 1 0 18492 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_195
timestamp 1688980957
transform 1 0 19044 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_197
timestamp 1688980957
transform 1 0 19228 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_209
timestamp 1688980957
transform 1 0 20332 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_221
timestamp 1688980957
transform 1 0 21436 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_233
timestamp 1688980957
transform 1 0 22540 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_245
timestamp 1688980957
transform 1 0 23644 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_251
timestamp 1688980957
transform 1 0 24196 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_253
timestamp 1688980957
transform 1 0 24380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_265
timestamp 1688980957
transform 1 0 25484 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_277
timestamp 1688980957
transform 1 0 26588 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_289
timestamp 1688980957
transform 1 0 27692 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_301
timestamp 1688980957
transform 1 0 28796 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_307
timestamp 1688980957
transform 1 0 29348 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_309
timestamp 1688980957
transform 1 0 29532 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_321
timestamp 1688980957
transform 1 0 30636 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_333
timestamp 1688980957
transform 1 0 31740 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_345
timestamp 1688980957
transform 1 0 32844 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_357
timestamp 1688980957
transform 1 0 33948 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_363
timestamp 1688980957
transform 1 0 34500 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_3
timestamp 1688980957
transform 1 0 1380 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_15
timestamp 1688980957
transform 1 0 2484 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_27
timestamp 1688980957
transform 1 0 3588 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_39
timestamp 1688980957
transform 1 0 4692 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_65_51
timestamp 1688980957
transform 1 0 5796 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_55
timestamp 1688980957
transform 1 0 6164 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_57
timestamp 1688980957
transform 1 0 6348 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_69
timestamp 1688980957
transform 1 0 7452 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_81
timestamp 1688980957
transform 1 0 8556 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_93
timestamp 1688980957
transform 1 0 9660 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_65_105
timestamp 1688980957
transform 1 0 10764 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_111
timestamp 1688980957
transform 1 0 11316 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_113
timestamp 1688980957
transform 1 0 11500 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_125
timestamp 1688980957
transform 1 0 12604 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_137
timestamp 1688980957
transform 1 0 13708 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_149
timestamp 1688980957
transform 1 0 14812 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_65_161
timestamp 1688980957
transform 1 0 15916 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_167
timestamp 1688980957
transform 1 0 16468 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_169
timestamp 1688980957
transform 1 0 16652 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_181
timestamp 1688980957
transform 1 0 17756 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_193
timestamp 1688980957
transform 1 0 18860 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_205
timestamp 1688980957
transform 1 0 19964 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_65_217
timestamp 1688980957
transform 1 0 21068 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_223
timestamp 1688980957
transform 1 0 21620 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_225
timestamp 1688980957
transform 1 0 21804 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_237
timestamp 1688980957
transform 1 0 22908 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_249
timestamp 1688980957
transform 1 0 24012 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_261
timestamp 1688980957
transform 1 0 25116 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_65_273
timestamp 1688980957
transform 1 0 26220 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_279
timestamp 1688980957
transform 1 0 26772 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_281
timestamp 1688980957
transform 1 0 26956 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_293
timestamp 1688980957
transform 1 0 28060 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_305
timestamp 1688980957
transform 1 0 29164 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_317
timestamp 1688980957
transform 1 0 30268 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_65_329
timestamp 1688980957
transform 1 0 31372 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_335
timestamp 1688980957
transform 1 0 31924 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_337
timestamp 1688980957
transform 1 0 32108 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_349
timestamp 1688980957
transform 1 0 33212 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_65_361
timestamp 1688980957
transform 1 0 34316 0 -1 38080
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_3
timestamp 1688980957
transform 1 0 1380 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_15
timestamp 1688980957
transform 1 0 2484 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_27
timestamp 1688980957
transform 1 0 3588 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_29
timestamp 1688980957
transform 1 0 3772 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_41
timestamp 1688980957
transform 1 0 4876 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_53
timestamp 1688980957
transform 1 0 5980 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_65
timestamp 1688980957
transform 1 0 7084 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_77
timestamp 1688980957
transform 1 0 8188 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_83
timestamp 1688980957
transform 1 0 8740 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_85
timestamp 1688980957
transform 1 0 8924 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_97
timestamp 1688980957
transform 1 0 10028 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_109
timestamp 1688980957
transform 1 0 11132 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_121
timestamp 1688980957
transform 1 0 12236 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_133
timestamp 1688980957
transform 1 0 13340 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_139
timestamp 1688980957
transform 1 0 13892 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_141
timestamp 1688980957
transform 1 0 14076 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_153
timestamp 1688980957
transform 1 0 15180 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_165
timestamp 1688980957
transform 1 0 16284 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_177
timestamp 1688980957
transform 1 0 17388 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_189
timestamp 1688980957
transform 1 0 18492 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_195
timestamp 1688980957
transform 1 0 19044 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_197
timestamp 1688980957
transform 1 0 19228 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_209
timestamp 1688980957
transform 1 0 20332 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_221
timestamp 1688980957
transform 1 0 21436 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_233
timestamp 1688980957
transform 1 0 22540 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_245
timestamp 1688980957
transform 1 0 23644 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_251
timestamp 1688980957
transform 1 0 24196 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_253
timestamp 1688980957
transform 1 0 24380 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_265
timestamp 1688980957
transform 1 0 25484 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_277
timestamp 1688980957
transform 1 0 26588 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_289
timestamp 1688980957
transform 1 0 27692 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_301
timestamp 1688980957
transform 1 0 28796 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_307
timestamp 1688980957
transform 1 0 29348 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_309
timestamp 1688980957
transform 1 0 29532 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_321
timestamp 1688980957
transform 1 0 30636 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_333
timestamp 1688980957
transform 1 0 31740 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_345
timestamp 1688980957
transform 1 0 32844 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_357
timestamp 1688980957
transform 1 0 33948 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_363
timestamp 1688980957
transform 1 0 34500 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_3
timestamp 1688980957
transform 1 0 1380 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_15
timestamp 1688980957
transform 1 0 2484 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_27
timestamp 1688980957
transform 1 0 3588 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_39
timestamp 1688980957
transform 1 0 4692 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_67_51
timestamp 1688980957
transform 1 0 5796 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_55
timestamp 1688980957
transform 1 0 6164 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_57
timestamp 1688980957
transform 1 0 6348 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_69
timestamp 1688980957
transform 1 0 7452 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_81
timestamp 1688980957
transform 1 0 8556 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_93
timestamp 1688980957
transform 1 0 9660 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_105
timestamp 1688980957
transform 1 0 10764 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_111
timestamp 1688980957
transform 1 0 11316 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_113
timestamp 1688980957
transform 1 0 11500 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_125
timestamp 1688980957
transform 1 0 12604 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_137
timestamp 1688980957
transform 1 0 13708 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_149
timestamp 1688980957
transform 1 0 14812 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_161
timestamp 1688980957
transform 1 0 15916 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_167
timestamp 1688980957
transform 1 0 16468 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_169
timestamp 1688980957
transform 1 0 16652 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_181
timestamp 1688980957
transform 1 0 17756 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_193
timestamp 1688980957
transform 1 0 18860 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_205
timestamp 1688980957
transform 1 0 19964 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_217
timestamp 1688980957
transform 1 0 21068 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_223
timestamp 1688980957
transform 1 0 21620 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_225
timestamp 1688980957
transform 1 0 21804 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_237
timestamp 1688980957
transform 1 0 22908 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_249
timestamp 1688980957
transform 1 0 24012 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_261
timestamp 1688980957
transform 1 0 25116 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_273
timestamp 1688980957
transform 1 0 26220 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_279
timestamp 1688980957
transform 1 0 26772 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_281
timestamp 1688980957
transform 1 0 26956 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_293
timestamp 1688980957
transform 1 0 28060 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_305
timestamp 1688980957
transform 1 0 29164 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_317
timestamp 1688980957
transform 1 0 30268 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_329
timestamp 1688980957
transform 1 0 31372 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_335
timestamp 1688980957
transform 1 0 31924 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_337
timestamp 1688980957
transform 1 0 32108 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_349
timestamp 1688980957
transform 1 0 33212 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_67_361
timestamp 1688980957
transform 1 0 34316 0 -1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_6
timestamp 1688980957
transform 1 0 1656 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_68_18
timestamp 1688980957
transform 1 0 2760 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_68_26
timestamp 1688980957
transform 1 0 3496 0 1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_29
timestamp 1688980957
transform 1 0 3772 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_41
timestamp 1688980957
transform 1 0 4876 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_68_53
timestamp 1688980957
transform 1 0 5980 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_68_57
timestamp 1688980957
transform 1 0 6348 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_65
timestamp 1688980957
transform 1 0 7084 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_70
timestamp 1688980957
transform 1 0 7544 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_68_82
timestamp 1688980957
transform 1 0 8648 0 1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_85
timestamp 1688980957
transform 1 0 8924 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_97
timestamp 1688980957
transform 1 0 10028 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_68_109
timestamp 1688980957
transform 1 0 11132 0 1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_113
timestamp 1688980957
transform 1 0 11500 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_125
timestamp 1688980957
transform 1 0 12604 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_68_137
timestamp 1688980957
transform 1 0 13708 0 1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_141
timestamp 1688980957
transform 1 0 14076 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_153
timestamp 1688980957
transform 1 0 15180 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_68_165
timestamp 1688980957
transform 1 0 16284 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_68_169
timestamp 1688980957
transform 1 0 16652 0 1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_174
timestamp 1688980957
transform 1 0 17112 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_68_186
timestamp 1688980957
transform 1 0 18216 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_68_194
timestamp 1688980957
transform 1 0 18952 0 1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_197
timestamp 1688980957
transform 1 0 19228 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_209
timestamp 1688980957
transform 1 0 20332 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_68_221
timestamp 1688980957
transform 1 0 21436 0 1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_225
timestamp 1688980957
transform 1 0 21804 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_237
timestamp 1688980957
transform 1 0 22908 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_68_249
timestamp 1688980957
transform 1 0 24012 0 1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_253
timestamp 1688980957
transform 1 0 24380 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_68_265
timestamp 1688980957
transform 1 0 25484 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_68_273
timestamp 1688980957
transform 1 0 26220 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_279
timestamp 1688980957
transform 1 0 26772 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_281
timestamp 1688980957
transform 1 0 26956 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_293
timestamp 1688980957
transform 1 0 28060 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_68_305
timestamp 1688980957
transform 1 0 29164 0 1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_309
timestamp 1688980957
transform 1 0 29532 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_321
timestamp 1688980957
transform 1 0 30636 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_68_333
timestamp 1688980957
transform 1 0 31740 0 1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_337
timestamp 1688980957
transform 1 0 32108 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_68_349
timestamp 1688980957
transform 1 0 33212 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_357
timestamp 1688980957
transform 1 0 33948 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input1
timestamp 1688980957
transform -1 0 34592 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input2
timestamp 1688980957
transform 1 0 1380 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1688980957
transform 1 0 34316 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input4
timestamp 1688980957
transform -1 0 34592 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input5
timestamp 1688980957
transform 1 0 16836 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input6 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1380 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1688980957
transform 1 0 28428 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input8
timestamp 1688980957
transform 1 0 7176 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output9
timestamp 1688980957
transform 1 0 34040 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output10
timestamp 1688980957
transform -1 0 19780 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output11
timestamp 1688980957
transform -1 0 1932 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output12
timestamp 1688980957
transform 1 0 34040 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1688980957
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1688980957
transform -1 0 34868 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1688980957
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1688980957
transform -1 0 34868 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1688980957
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1688980957
transform -1 0 34868 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1688980957
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1688980957
transform -1 0 34868 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1688980957
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1688980957
transform -1 0 34868 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1688980957
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1688980957
transform -1 0 34868 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1688980957
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1688980957
transform -1 0 34868 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1688980957
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1688980957
transform -1 0 34868 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1688980957
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1688980957
transform -1 0 34868 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1688980957
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1688980957
transform -1 0 34868 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1688980957
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1688980957
transform -1 0 34868 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1688980957
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1688980957
transform -1 0 34868 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1688980957
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1688980957
transform -1 0 34868 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1688980957
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1688980957
transform -1 0 34868 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1688980957
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1688980957
transform -1 0 34868 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1688980957
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1688980957
transform -1 0 34868 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1688980957
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1688980957
transform -1 0 34868 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1688980957
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1688980957
transform -1 0 34868 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1688980957
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1688980957
transform -1 0 34868 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1688980957
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1688980957
transform -1 0 34868 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1688980957
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1688980957
transform -1 0 34868 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1688980957
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1688980957
transform -1 0 34868 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1688980957
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1688980957
transform -1 0 34868 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1688980957
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1688980957
transform -1 0 34868 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1688980957
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1688980957
transform -1 0 34868 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1688980957
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1688980957
transform -1 0 34868 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1688980957
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1688980957
transform -1 0 34868 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1688980957
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1688980957
transform -1 0 34868 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1688980957
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1688980957
transform -1 0 34868 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1688980957
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1688980957
transform -1 0 34868 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1688980957
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1688980957
transform -1 0 34868 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1688980957
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1688980957
transform -1 0 34868 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1688980957
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1688980957
transform -1 0 34868 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1688980957
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1688980957
transform -1 0 34868 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1688980957
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1688980957
transform -1 0 34868 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1688980957
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1688980957
transform -1 0 34868 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1688980957
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1688980957
transform -1 0 34868 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1688980957
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1688980957
transform -1 0 34868 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1688980957
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1688980957
transform -1 0 34868 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1688980957
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1688980957
transform -1 0 34868 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1688980957
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1688980957
transform -1 0 34868 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1688980957
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1688980957
transform -1 0 34868 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1688980957
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1688980957
transform -1 0 34868 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1688980957
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1688980957
transform -1 0 34868 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1688980957
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1688980957
transform -1 0 34868 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1688980957
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1688980957
transform -1 0 34868 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1688980957
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1688980957
transform -1 0 34868 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1688980957
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1688980957
transform -1 0 34868 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1688980957
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1688980957
transform -1 0 34868 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1688980957
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1688980957
transform -1 0 34868 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1688980957
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1688980957
transform -1 0 34868 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1688980957
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1688980957
transform -1 0 34868 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1688980957
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1688980957
transform -1 0 34868 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1688980957
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1688980957
transform -1 0 34868 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1688980957
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1688980957
transform -1 0 34868 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1688980957
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1688980957
transform -1 0 34868 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1688980957
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1688980957
transform -1 0 34868 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1688980957
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1688980957
transform -1 0 34868 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1688980957
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1688980957
transform -1 0 34868 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1688980957
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1688980957
transform -1 0 34868 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1688980957
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1688980957
transform -1 0 34868 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1688980957
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1688980957
transform -1 0 34868 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1688980957
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1688980957
transform -1 0 34868 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1688980957
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1688980957
transform -1 0 34868 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1688980957
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1688980957
transform -1 0 34868 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1688980957
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1688980957
transform -1 0 34868 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1688980957
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1688980957
transform -1 0 34868 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1688980957
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1688980957
transform -1 0 34868 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1688980957
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1688980957
transform -1 0 34868 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rgb_mixer_28
timestamp 1688980957
transform -1 0 9384 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rgb_mixer_29
timestamp 1688980957
transform -1 0 26772 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rgb_mixer_30
timestamp 1688980957
transform -1 0 1656 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rgb_mixer_31
timestamp 1688980957
transform -1 0 1656 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1688980957
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1688980957
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1688980957
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1688980957
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1688980957
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1688980957
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1688980957
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1688980957
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1688980957
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1688980957
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1688980957
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1688980957
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1688980957
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1688980957
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1688980957
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1688980957
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1688980957
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1688980957
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1688980957
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1688980957
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1688980957
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1688980957
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1688980957
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1688980957
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1688980957
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1688980957
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1688980957
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1688980957
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1688980957
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1688980957
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1688980957
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1688980957
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1688980957
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1688980957
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1688980957
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1688980957
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1688980957
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1688980957
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1688980957
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1688980957
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1688980957
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1688980957
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1688980957
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1688980957
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1688980957
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1688980957
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1688980957
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1688980957
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1688980957
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1688980957
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1688980957
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1688980957
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1688980957
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1688980957
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1688980957
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1688980957
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1688980957
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1688980957
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1688980957
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1688980957
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1688980957
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1688980957
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1688980957
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1688980957
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1688980957
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1688980957
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1688980957
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1688980957
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1688980957
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1688980957
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1688980957
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1688980957
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1688980957
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1688980957
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1688980957
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1688980957
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1688980957
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1688980957
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1688980957
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1688980957
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1688980957
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1688980957
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1688980957
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1688980957
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1688980957
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1688980957
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1688980957
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1688980957
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1688980957
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1688980957
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1688980957
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1688980957
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1688980957
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1688980957
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1688980957
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1688980957
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1688980957
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1688980957
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1688980957
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1688980957
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1688980957
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1688980957
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1688980957
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1688980957
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1688980957
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1688980957
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1688980957
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1688980957
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1688980957
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1688980957
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1688980957
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1688980957
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1688980957
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1688980957
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1688980957
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1688980957
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1688980957
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1688980957
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1688980957
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1688980957
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1688980957
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1688980957
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1688980957
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1688980957
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1688980957
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1688980957
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1688980957
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1688980957
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1688980957
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1688980957
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1688980957
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1688980957
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1688980957
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1688980957
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1688980957
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1688980957
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1688980957
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1688980957
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1688980957
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1688980957
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1688980957
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1688980957
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1688980957
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1688980957
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1688980957
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1688980957
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1688980957
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1688980957
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1688980957
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1688980957
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1688980957
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1688980957
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1688980957
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1688980957
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1688980957
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1688980957
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1688980957
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1688980957
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1688980957
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1688980957
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1688980957
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1688980957
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1688980957
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1688980957
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1688980957
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1688980957
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1688980957
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1688980957
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1688980957
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1688980957
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1688980957
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1688980957
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1688980957
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1688980957
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1688980957
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1688980957
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1688980957
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1688980957
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1688980957
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1688980957
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1688980957
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1688980957
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1688980957
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1688980957
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1688980957
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1688980957
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1688980957
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1688980957
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1688980957
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1688980957
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1688980957
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1688980957
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1688980957
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1688980957
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1688980957
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1688980957
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1688980957
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1688980957
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1688980957
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1688980957
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1688980957
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1688980957
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1688980957
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1688980957
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1688980957
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1688980957
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1688980957
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1688980957
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1688980957
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1688980957
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1688980957
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1688980957
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1688980957
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1688980957
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1688980957
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1688980957
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1688980957
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1688980957
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1688980957
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1688980957
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1688980957
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1688980957
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1688980957
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1688980957
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1688980957
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1688980957
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1688980957
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1688980957
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1688980957
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1688980957
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1688980957
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1688980957
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1688980957
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1688980957
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1688980957
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1688980957
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1688980957
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1688980957
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1688980957
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1688980957
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1688980957
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1688980957
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1688980957
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1688980957
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1688980957
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1688980957
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1688980957
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1688980957
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1688980957
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1688980957
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1688980957
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1688980957
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1688980957
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1688980957
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1688980957
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1688980957
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1688980957
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1688980957
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1688980957
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1688980957
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1688980957
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1688980957
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1688980957
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1688980957
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1688980957
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1688980957
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1688980957
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1688980957
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1688980957
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1688980957
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1688980957
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1688980957
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1688980957
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1688980957
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1688980957
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1688980957
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1688980957
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1688980957
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1688980957
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1688980957
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1688980957
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1688980957
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1688980957
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1688980957
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1688980957
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1688980957
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1688980957
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1688980957
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1688980957
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1688980957
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1688980957
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1688980957
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1688980957
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1688980957
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1688980957
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1688980957
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1688980957
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1688980957
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1688980957
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1688980957
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1688980957
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1688980957
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1688980957
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1688980957
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1688980957
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1688980957
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1688980957
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1688980957
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1688980957
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1688980957
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1688980957
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1688980957
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1688980957
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1688980957
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1688980957
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1688980957
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1688980957
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1688980957
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1688980957
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1688980957
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1688980957
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1688980957
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1688980957
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1688980957
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1688980957
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1688980957
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1688980957
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1688980957
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1688980957
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1688980957
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1688980957
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1688980957
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1688980957
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1688980957
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1688980957
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1688980957
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1688980957
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1688980957
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1688980957
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1688980957
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1688980957
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1688980957
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1688980957
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1688980957
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1688980957
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1688980957
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1688980957
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1688980957
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1688980957
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1688980957
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1688980957
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1688980957
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1688980957
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1688980957
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1688980957
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1688980957
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1688980957
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1688980957
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1688980957
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1688980957
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1688980957
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1688980957
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1688980957
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1688980957
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1688980957
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1688980957
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1688980957
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1688980957
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1688980957
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1688980957
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1688980957
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1688980957
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1688980957
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1688980957
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1688980957
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1688980957
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1688980957
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1688980957
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1688980957
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1688980957
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1688980957
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1688980957
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1688980957
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1688980957
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1688980957
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1688980957
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1688980957
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1688980957
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1688980957
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1688980957
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1688980957
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1688980957
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1688980957
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1688980957
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1688980957
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1688980957
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1688980957
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1688980957
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1688980957
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1688980957
transform 1 0 26864 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1688980957
transform 1 0 32016 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1688980957
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1688980957
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1688980957
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1688980957
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1688980957
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1688980957
transform 1 0 29440 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1688980957
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1688980957
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1688980957
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1688980957
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1688980957
transform 1 0 26864 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1688980957
transform 1 0 32016 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1688980957
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1688980957
transform 1 0 6256 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1688980957
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1688980957
transform 1 0 11408 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1688980957
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1688980957
transform 1 0 16560 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1688980957
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1688980957
transform 1 0 21712 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1688980957
transform 1 0 24288 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1688980957
transform 1 0 26864 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1688980957
transform 1 0 29440 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1688980957
transform 1 0 32016 0 1 39168
box -38 -48 130 592
<< labels >>
flabel metal3 s 35200 21708 36000 21948 0 FreeSans 960 0 0 0 clk
port 0 nsew signal input
flabel metal3 s 0 39388 800 39628 0 FreeSans 960 0 0 0 enc0_a
port 1 nsew signal input
flabel metal3 s 35200 31908 36000 32148 0 FreeSans 960 0 0 0 enc0_b
port 2 nsew signal input
flabel metal3 s 35200 1988 36000 2228 0 FreeSans 960 0 0 0 enc1_a
port 3 nsew signal input
flabel metal2 s 16734 41200 16846 42000 0 FreeSans 448 90 0 0 enc1_b
port 4 nsew signal input
flabel metal2 s -10 0 102 800 0 FreeSans 448 90 0 0 enc2_a
port 5 nsew signal input
flabel metal2 s 28326 0 28438 800 0 FreeSans 448 90 0 0 enc2_b
port 6 nsew signal input
flabel metal2 s 9006 0 9118 800 0 FreeSans 448 90 0 0 io_oeb[0]
port 7 nsew signal tristate
flabel metal2 s 26394 41200 26506 42000 0 FreeSans 448 90 0 0 io_oeb[1]
port 8 nsew signal tristate
flabel metal3 s 0 9468 800 9708 0 FreeSans 960 0 0 0 io_oeb[2]
port 9 nsew signal tristate
flabel metal3 s 0 19668 800 19908 0 FreeSans 960 0 0 0 io_oeb[3]
port 10 nsew signal tristate
flabel metal2 s 35410 41200 35522 42000 0 FreeSans 448 90 0 0 pwm0_out
port 11 nsew signal tristate
flabel metal2 s 18666 0 18778 800 0 FreeSans 448 90 0 0 pwm1_out
port 12 nsew signal tristate
flabel metal3 s 0 29868 800 30108 0 FreeSans 960 0 0 0 pwm2_out
port 13 nsew signal tristate
flabel metal2 s 7074 41200 7186 42000 0 FreeSans 448 90 0 0 reset
port 14 nsew signal input
flabel metal3 s 35200 11508 36000 11748 0 FreeSans 960 0 0 0 sync
port 15 nsew signal tristate
flabel metal4 s 5164 2128 5484 39760 0 FreeSans 1920 90 0 0 vccd1
port 16 nsew power bidirectional
flabel metal4 s 13605 2128 13925 39760 0 FreeSans 1920 90 0 0 vccd1
port 16 nsew power bidirectional
flabel metal4 s 22046 2128 22366 39760 0 FreeSans 1920 90 0 0 vccd1
port 16 nsew power bidirectional
flabel metal4 s 30487 2128 30807 39760 0 FreeSans 1920 90 0 0 vccd1
port 16 nsew power bidirectional
flabel metal4 s 9384 2128 9704 39760 0 FreeSans 1920 90 0 0 vssd1
port 17 nsew ground bidirectional
flabel metal4 s 17825 2128 18145 39760 0 FreeSans 1920 90 0 0 vssd1
port 17 nsew ground bidirectional
flabel metal4 s 26266 2128 26586 39760 0 FreeSans 1920 90 0 0 vssd1
port 17 nsew ground bidirectional
flabel metal4 s 34707 2128 35027 39760 0 FreeSans 1920 90 0 0 vssd1
port 17 nsew ground bidirectional
rlabel metal1 17986 39712 17986 39712 0 vccd1
rlabel via1 18065 39168 18065 39168 0 vssd1
rlabel metal1 16192 17306 16192 17306 0 _000_
rlabel via1 29849 29614 29849 29614 0 _001_
rlabel metal1 25652 32810 25652 32810 0 _002_
rlabel via1 29128 32402 29128 32402 0 _003_
rlabel metal2 29578 33286 29578 33286 0 _004_
rlabel metal1 31157 32810 31157 32810 0 _005_
rlabel metal1 30815 32470 30815 32470 0 _006_
rlabel via1 29849 30702 29849 30702 0 _007_
rlabel metal2 31418 30498 31418 30498 0 _008_
rlabel metal2 32706 31110 32706 31110 0 _009_
rlabel metal2 31786 25058 31786 25058 0 _010_
rlabel via1 31597 29614 31597 29614 0 _011_
rlabel via1 31873 28526 31873 28526 0 _012_
rlabel metal2 30406 28322 30406 28322 0 _013_
rlabel via1 31321 27438 31321 27438 0 _014_
rlabel via1 32241 26350 32241 26350 0 _015_
rlabel metal1 30677 25262 30677 25262 0 _016_
rlabel metal1 31091 23766 31091 23766 0 _017_
rlabel metal2 32614 23970 32614 23970 0 _018_
rlabel via1 30861 20910 30861 20910 0 _019_
rlabel metal2 31510 16082 31510 16082 0 _020_
rlabel metal1 31367 19754 31367 19754 0 _021_
rlabel metal1 30666 19414 30666 19414 0 _022_
rlabel metal1 32839 19414 32839 19414 0 _023_
rlabel metal2 33350 20706 33350 20706 0 _024_
rlabel metal1 30176 21862 30176 21862 0 _025_
rlabel metal1 30907 22678 30907 22678 0 _026_
rlabel metal1 33023 21930 33023 21930 0 _027_
rlabel metal2 27094 21318 27094 21318 0 _028_
rlabel metal1 24876 24174 24876 24174 0 _029_
rlabel metal1 26261 23018 26261 23018 0 _030_
rlabel metal1 27032 23766 27032 23766 0 _031_
rlabel metal2 29026 22882 29026 22882 0 _032_
rlabel metal2 28382 21726 28382 21726 0 _033_
rlabel metal1 26077 19822 26077 19822 0 _034_
rlabel metal1 27084 19822 27084 19822 0 _035_
rlabel metal1 28888 20570 28888 20570 0 _036_
rlabel metal2 25530 18870 25530 18870 0 _037_
rlabel metal1 23368 14586 23368 14586 0 _038_
rlabel metal1 24656 14586 24656 14586 0 _039_
rlabel metal1 24502 15062 24502 15062 0 _040_
rlabel metal2 26726 15266 26726 15266 0 _041_
rlabel metal1 27466 16150 27466 16150 0 _042_
rlabel via1 24697 17646 24697 17646 0 _043_
rlabel metal1 25806 17272 25806 17272 0 _044_
rlabel metal1 28202 17646 28202 17646 0 _045_
rlabel metal2 29394 19618 29394 19618 0 _046_
rlabel via1 16969 24854 16969 24854 0 _047_
rlabel via1 17337 24174 17337 24174 0 _048_
rlabel metal1 16739 26350 16739 26350 0 _049_
rlabel metal1 17245 27438 17245 27438 0 _050_
rlabel metal2 16882 28322 16882 28322 0 _051_
rlabel metal1 16744 29818 16744 29818 0 _052_
rlabel metal2 16790 31110 16790 31110 0 _053_
rlabel via1 17337 31790 17337 31790 0 _054_
rlabel metal1 29895 23018 29895 23018 0 _055_
rlabel metal1 27963 15062 27963 15062 0 _056_
rlabel metal1 28596 16150 28596 16150 0 _057_
rlabel metal2 29762 15878 29762 15878 0 _058_
rlabel metal1 30314 15130 30314 15130 0 _059_
rlabel metal2 30866 17442 30866 17442 0 _060_
rlabel metal1 27600 18394 27600 18394 0 _061_
rlabel viali 28561 18258 28561 18258 0 _062_
rlabel metal1 30130 17850 30130 17850 0 _063_
rlabel metal1 25944 24922 25944 24922 0 _064_
rlabel metal1 27641 25262 27641 25262 0 _065_
rlabel metal1 30042 27370 30042 27370 0 _066_
rlabel metal2 25990 27846 25990 27846 0 _067_
rlabel metal2 28934 29410 28934 29410 0 _068_
rlabel metal1 26914 29614 26914 29614 0 _069_
rlabel metal1 24600 32878 24600 32878 0 _070_
rlabel metal1 25458 32470 25458 32470 0 _071_
rlabel metal1 25852 21658 25852 21658 0 _072_
rlabel metal1 29026 24378 29026 24378 0 _073_
rlabel metal2 20378 21794 20378 21794 0 _074_
rlabel metal1 21932 21998 21932 21998 0 _075_
rlabel via1 23133 19822 23133 19822 0 _076_
rlabel metal2 20194 19142 20194 19142 0 _077_
rlabel metal2 23874 19142 23874 19142 0 _078_
rlabel metal1 24108 17170 24108 17170 0 _079_
rlabel metal1 19499 16150 19499 16150 0 _080_
rlabel via1 20097 14994 20097 14994 0 _081_
rlabel metal2 24426 23494 24426 23494 0 _082_
rlabel metal2 24426 21726 24426 21726 0 _083_
rlabel metal2 19274 24582 19274 24582 0 _084_
rlabel metal1 20270 23766 20270 23766 0 _085_
rlabel metal2 22494 26758 22494 26758 0 _086_
rlabel via1 19462 27030 19462 27030 0 _087_
rlabel metal1 21808 28458 21808 28458 0 _088_
rlabel metal1 22222 30226 22222 30226 0 _089_
rlabel metal1 18860 31994 18860 31994 0 _090_
rlabel metal2 21758 32198 21758 32198 0 _091_
rlabel metal1 22356 23290 22356 23290 0 _092_
rlabel metal1 22816 25466 22816 25466 0 _093_
rlabel metal2 24702 25670 24702 25670 0 _094_
rlabel metal1 23036 26350 23036 26350 0 _095_
rlabel metal1 24150 27642 24150 27642 0 _096_
rlabel metal2 22954 27846 22954 27846 0 _097_
rlabel metal2 22678 30226 22678 30226 0 _098_
rlabel metal1 23368 29818 23368 29818 0 _099_
rlabel metal1 24283 31314 24283 31314 0 _100_
rlabel metal1 17337 22678 17337 22678 0 _101_
rlabel metal1 19500 22746 19500 22746 0 _102_
rlabel metal1 17521 21930 17521 21930 0 _103_
rlabel metal1 18022 20434 18022 20434 0 _104_
rlabel metal1 17633 19754 17633 19754 0 _105_
rlabel metal1 17015 18666 17015 18666 0 _106_
rlabel metal1 17061 17238 17061 17238 0 _107_
rlabel metal1 17802 16150 17802 16150 0 _108_
rlabel metal1 25254 30804 25254 30804 0 _109_
rlabel metal1 25530 30124 25530 30124 0 _110_
rlabel metal1 25714 30736 25714 30736 0 _111_
rlabel metal1 25346 30260 25346 30260 0 _112_
rlabel metal2 25530 29070 25530 29070 0 _113_
rlabel metal1 25346 28560 25346 28560 0 _114_
rlabel metal1 24886 27098 24886 27098 0 _115_
rlabel metal1 25622 27472 25622 27472 0 _116_
rlabel metal2 25714 25636 25714 25636 0 _117_
rlabel metal1 25714 26554 25714 26554 0 _118_
rlabel metal1 25024 25398 25024 25398 0 _119_
rlabel metal1 25300 26554 25300 26554 0 _120_
rlabel metal1 25852 27098 25852 27098 0 _121_
rlabel metal1 25208 27642 25208 27642 0 _122_
rlabel metal1 25852 28730 25852 28730 0 _123_
rlabel metal2 25162 30022 25162 30022 0 _124_
rlabel metal1 25852 30362 25852 30362 0 _125_
rlabel metal1 17250 19278 17250 19278 0 _126_
rlabel metal1 26404 21998 26404 21998 0 _127_
rlabel metal2 29578 23392 29578 23392 0 _128_
rlabel metal1 25760 23834 25760 23834 0 _129_
rlabel metal1 19412 16422 19412 16422 0 _130_
rlabel metal1 18906 17204 18906 17204 0 _131_
rlabel viali 19089 18258 19089 18258 0 _132_
rlabel metal2 18998 19142 18998 19142 0 _133_
rlabel metal1 19872 20026 19872 20026 0 _134_
rlabel metal1 19090 19448 19090 19448 0 _135_
rlabel metal1 20010 20570 20010 20570 0 _136_
rlabel metal1 20010 21114 20010 21114 0 _137_
rlabel metal1 19458 21454 19458 21454 0 _138_
rlabel metal2 19918 21692 19918 21692 0 _139_
rlabel metal1 20102 21556 20102 21556 0 _140_
rlabel metal1 20194 20434 20194 20434 0 _141_
rlabel metal1 19366 19346 19366 19346 0 _142_
rlabel metal1 19228 18734 19228 18734 0 _143_
rlabel metal1 19596 18258 19596 18258 0 _144_
rlabel metal1 18630 17204 18630 17204 0 _145_
rlabel metal1 19458 16762 19458 16762 0 _146_
rlabel metal1 20010 16592 20010 16592 0 _147_
rlabel metal1 19918 30702 19918 30702 0 _148_
rlabel metal2 19550 30498 19550 30498 0 _149_
rlabel metal1 18354 29648 18354 29648 0 _150_
rlabel metal1 18860 29274 18860 29274 0 _151_
rlabel metal2 18998 27166 18998 27166 0 _152_
rlabel metal1 18538 28186 18538 28186 0 _153_
rlabel metal1 18032 25874 18032 25874 0 _154_
rlabel metal1 18768 25262 18768 25262 0 _155_
rlabel metal1 19826 25738 19826 25738 0 _156_
rlabel metal1 18584 25466 18584 25466 0 _157_
rlabel metal1 18308 25262 18308 25262 0 _158_
rlabel metal1 18170 25466 18170 25466 0 _159_
rlabel metal2 18262 27812 18262 27812 0 _160_
rlabel metal1 18860 28730 18860 28730 0 _161_
rlabel metal1 18262 29818 18262 29818 0 _162_
rlabel metal1 19044 30362 19044 30362 0 _163_
rlabel metal2 19274 30617 19274 30617 0 _164_
rlabel metal1 30360 33286 30360 33286 0 _165_
rlabel metal1 30222 30260 30222 30260 0 _166_
rlabel metal1 30728 32198 30728 32198 0 _167_
rlabel metal1 30314 30260 30314 30260 0 _168_
rlabel metal1 26450 20842 26450 20842 0 _169_
rlabel metal1 27922 14348 27922 14348 0 _170_
rlabel metal1 23552 32878 23552 32878 0 _171_
rlabel metal1 29256 32878 29256 32878 0 _172_
rlabel metal1 29440 31994 29440 31994 0 _173_
rlabel metal1 31418 32878 31418 32878 0 _174_
rlabel metal1 31786 26928 31786 26928 0 _175_
rlabel metal1 31096 31994 31096 31994 0 _176_
rlabel metal1 30130 31314 30130 31314 0 _177_
rlabel metal1 31096 30226 31096 30226 0 _178_
rlabel metal1 32338 30702 32338 30702 0 _179_
rlabel metal1 32246 27846 32246 27846 0 _180_
rlabel metal1 31418 24752 31418 24752 0 _181_
rlabel metal2 32798 26826 32798 26826 0 _182_
rlabel metal1 31326 24718 31326 24718 0 _183_
rlabel metal2 31878 31008 31878 31008 0 _184_
rlabel metal1 31878 29138 31878 29138 0 _185_
rlabel metal1 30636 28050 30636 28050 0 _186_
rlabel metal1 31188 27098 31188 27098 0 _187_
rlabel metal1 32246 26962 32246 26962 0 _188_
rlabel metal1 31004 25874 31004 25874 0 _189_
rlabel metal1 31510 24208 31510 24208 0 _190_
rlabel metal1 30498 22032 30498 22032 0 _191_
rlabel metal1 32660 23698 32660 23698 0 _192_
rlabel metal1 32568 20570 32568 20570 0 _193_
rlabel metal2 31142 21828 31142 21828 0 _194_
rlabel metal1 33350 19754 33350 19754 0 _195_
rlabel metal1 31234 21522 31234 21522 0 _196_
rlabel metal2 31694 15300 31694 15300 0 _197_
rlabel metal1 31464 20434 31464 20434 0 _198_
rlabel metal2 31234 19142 31234 19142 0 _199_
rlabel metal1 32936 18938 32936 18938 0 _200_
rlabel metal2 33534 20230 33534 20230 0 _201_
rlabel metal1 29992 21114 29992 21114 0 _202_
rlabel metal1 30958 22202 30958 22202 0 _203_
rlabel metal1 33074 21998 33074 21998 0 _204_
rlabel metal1 27462 21114 27462 21114 0 _205_
rlabel metal1 26726 20944 26726 20944 0 _206_
rlabel metal2 27922 21257 27922 21257 0 _207_
rlabel metal1 26956 20570 26956 20570 0 _208_
rlabel metal1 23966 24786 23966 24786 0 _209_
rlabel metal1 26588 22746 26588 22746 0 _210_
rlabel metal1 26910 22066 26910 22066 0 _211_
rlabel metal2 28198 19924 28198 19924 0 _212_
rlabel metal1 28842 22576 28842 22576 0 _213_
rlabel metal2 28198 22039 28198 22039 0 _214_
rlabel metal1 26496 20434 26496 20434 0 _215_
rlabel metal1 27278 19482 27278 19482 0 _216_
rlabel metal1 28474 20434 28474 20434 0 _217_
rlabel metal1 26542 15130 26542 15130 0 _218_
rlabel metal2 25898 17782 25898 17782 0 _219_
rlabel metal2 26174 16371 26174 16371 0 _220_
rlabel metal1 25990 16762 25990 16762 0 _221_
rlabel metal1 23046 14382 23046 14382 0 _222_
rlabel metal1 24472 14382 24472 14382 0 _223_
rlabel metal1 24058 15572 24058 15572 0 _224_
rlabel metal1 26358 14586 26358 14586 0 _225_
rlabel metal1 26772 16082 26772 16082 0 _226_
rlabel metal1 25024 17306 25024 17306 0 _227_
rlabel metal1 28014 21930 28014 21930 0 _228_
rlabel metal1 25852 17170 25852 17170 0 _229_
rlabel metal2 27002 17782 27002 17782 0 _230_
rlabel metal1 29072 16422 29072 16422 0 _231_
rlabel metal1 29302 18938 29302 18938 0 _232_
rlabel metal1 30038 16762 30038 16762 0 _233_
rlabel metal2 29302 18360 29302 18360 0 _234_
rlabel metal1 20930 17238 20930 17238 0 _235_
rlabel metal1 18216 24922 18216 24922 0 _236_
rlabel metal1 17296 26826 17296 26826 0 _237_
rlabel metal1 17434 25772 17434 25772 0 _238_
rlabel metal1 17664 28118 17664 28118 0 _239_
rlabel metal1 18216 27642 18216 27642 0 _240_
rlabel metal1 20976 21522 20976 21522 0 _241_
rlabel metal1 17066 29172 17066 29172 0 _242_
rlabel metal2 17066 28492 17066 28492 0 _243_
rlabel metal1 17204 29818 17204 29818 0 _244_
rlabel metal1 16698 29614 16698 29614 0 _245_
rlabel metal2 17802 31969 17802 31969 0 _246_
rlabel metal1 16974 30736 16974 30736 0 _247_
rlabel metal1 17986 32402 17986 32402 0 _248_
rlabel metal1 29992 23698 29992 23698 0 _249_
rlabel metal1 28244 14586 28244 14586 0 _250_
rlabel metal1 28336 15674 28336 15674 0 _251_
rlabel metal1 29394 15470 29394 15470 0 _252_
rlabel metal1 30636 14994 30636 14994 0 _253_
rlabel metal1 30498 16694 30498 16694 0 _254_
rlabel metal1 27784 18258 27784 18258 0 _255_
rlabel metal1 28566 18938 28566 18938 0 _256_
rlabel metal1 29992 17646 29992 17646 0 _257_
rlabel metal1 29992 25874 29992 25874 0 _258_
rlabel metal1 29854 25874 29854 25874 0 _259_
rlabel metal1 30038 25738 30038 25738 0 _260_
rlabel metal1 30176 25874 30176 25874 0 _261_
rlabel metal1 26956 31994 26956 31994 0 _262_
rlabel metal1 26358 27472 26358 27472 0 _263_
rlabel metal2 26082 25228 26082 25228 0 _264_
rlabel metal1 28842 25840 28842 25840 0 _265_
rlabel metal1 27830 26282 27830 26282 0 _266_
rlabel metal1 28512 26010 28512 26010 0 _267_
rlabel metal1 26772 25738 26772 25738 0 _268_
rlabel metal1 27324 25738 27324 25738 0 _269_
rlabel metal1 27324 26010 27324 26010 0 _270_
rlabel metal1 27922 28050 27922 28050 0 _271_
rlabel metal1 29164 27098 29164 27098 0 _272_
rlabel via1 27738 28594 27738 28594 0 _273_
rlabel metal2 29026 28390 29026 28390 0 _274_
rlabel metal1 28934 27982 28934 27982 0 _275_
rlabel metal1 29394 27030 29394 27030 0 _276_
rlabel metal1 29118 27030 29118 27030 0 _277_
rlabel metal1 27692 27914 27692 27914 0 _278_
rlabel metal1 27968 27642 27968 27642 0 _279_
rlabel metal1 27278 27404 27278 27404 0 _280_
rlabel metal1 26450 27404 26450 27404 0 _281_
rlabel metal1 27646 28050 27646 28050 0 _282_
rlabel metal2 28842 29444 28842 29444 0 _283_
rlabel metal1 28336 30838 28336 30838 0 _284_
rlabel metal2 28566 30396 28566 30396 0 _285_
rlabel metal1 28060 30226 28060 30226 0 _286_
rlabel metal1 28417 29141 28417 29141 0 _287_
rlabel metal1 27416 30226 27416 30226 0 _288_
rlabel metal1 28658 30158 28658 30158 0 _289_
rlabel metal1 26174 30260 26174 30260 0 _290_
rlabel metal1 26266 30124 26266 30124 0 _291_
rlabel metal1 26542 31790 26542 31790 0 _292_
rlabel metal1 27002 33558 27002 33558 0 _293_
rlabel via1 27002 33014 27002 33014 0 _294_
rlabel metal1 26956 32946 26956 32946 0 _295_
rlabel metal1 27692 29818 27692 29818 0 _296_
rlabel metal2 27416 32402 27416 32402 0 _297_
rlabel via1 26266 32861 26266 32861 0 _298_
rlabel metal2 26174 32300 26174 32300 0 _299_
rlabel metal1 24196 32878 24196 32878 0 _300_
rlabel metal1 24104 33082 24104 33082 0 _301_
rlabel metal1 26404 33354 26404 33354 0 _302_
rlabel metal1 25990 32436 25990 32436 0 _303_
rlabel metal1 26082 32436 26082 32436 0 _304_
rlabel metal1 25438 21522 25438 21522 0 _305_
rlabel metal1 28934 24174 28934 24174 0 _306_
rlabel metal1 25116 20978 25116 20978 0 _307_
rlabel metal1 24564 21658 24564 21658 0 _308_
rlabel metal1 24656 20842 24656 20842 0 _309_
rlabel metal1 25019 20910 25019 20910 0 _310_
rlabel metal2 21206 21148 21206 21148 0 _311_
rlabel metal1 20792 21318 20792 21318 0 _312_
rlabel metal1 20562 21454 20562 21454 0 _313_
rlabel metal2 23046 21318 23046 21318 0 _314_
rlabel metal1 21528 21318 21528 21318 0 _315_
rlabel metal1 21896 21454 21896 21454 0 _316_
rlabel metal2 21390 22406 21390 22406 0 _317_
rlabel metal2 21666 21869 21666 21869 0 _318_
rlabel metal1 22310 22644 22310 22644 0 _319_
rlabel metal2 22402 20740 22402 20740 0 _320_
rlabel metal1 22770 19924 22770 19924 0 _321_
rlabel metal1 22632 16626 22632 16626 0 _322_
rlabel metal1 21574 19822 21574 19822 0 _323_
rlabel metal1 22172 19210 22172 19210 0 _324_
rlabel metal1 22448 20026 22448 20026 0 _325_
rlabel metal1 23598 20400 23598 20400 0 _326_
rlabel metal1 21528 19482 21528 19482 0 _327_
rlabel metal1 21666 19686 21666 19686 0 _328_
rlabel metal1 21390 18598 21390 18598 0 _329_
rlabel metal1 20700 18734 20700 18734 0 _330_
rlabel metal1 21436 18938 21436 18938 0 _331_
rlabel metal1 22540 18258 22540 18258 0 _332_
rlabel metal1 22310 17578 22310 17578 0 _333_
rlabel metal1 23230 17612 23230 17612 0 _334_
rlabel metal2 22310 17340 22310 17340 0 _335_
rlabel metal1 23736 17646 23736 17646 0 _336_
rlabel metal1 22954 17850 22954 17850 0 _337_
rlabel metal2 23966 18258 23966 18258 0 _338_
rlabel metal1 22678 17034 22678 17034 0 _339_
rlabel metal1 22954 17204 22954 17204 0 _340_
rlabel metal1 23000 16762 23000 16762 0 _341_
rlabel metal1 21528 16558 21528 16558 0 _342_
rlabel metal1 21298 17612 21298 17612 0 _343_
rlabel metal1 21298 17068 21298 17068 0 _344_
rlabel metal1 22540 16762 22540 16762 0 _345_
rlabel metal1 21620 17170 21620 17170 0 _346_
rlabel metal1 20171 17782 20171 17782 0 _347_
rlabel metal1 19872 17170 19872 17170 0 _348_
rlabel metal1 19826 16592 19826 16592 0 _349_
rlabel metal1 21022 17680 21022 17680 0 _350_
rlabel metal1 20792 17170 20792 17170 0 _351_
rlabel metal1 20654 17204 20654 17204 0 _352_
rlabel metal1 24380 23086 24380 23086 0 _353_
rlabel metal1 24472 21998 24472 21998 0 _354_
rlabel metal2 23598 23732 23598 23732 0 _355_
rlabel metal1 23322 24106 23322 24106 0 _356_
rlabel metal1 22586 24208 22586 24208 0 _357_
rlabel metal1 22678 24140 22678 24140 0 _358_
rlabel metal1 20838 31858 20838 31858 0 _359_
rlabel metal2 21436 31756 21436 31756 0 _360_
rlabel metal1 19412 24174 19412 24174 0 _361_
rlabel metal2 21482 25534 21482 25534 0 _362_
rlabel metal1 21022 25126 21022 25126 0 _363_
rlabel metal1 20286 24684 20286 24684 0 _364_
rlabel metal2 20930 24786 20930 24786 0 _365_
rlabel metal1 21068 24378 21068 24378 0 _366_
rlabel metal1 20654 24140 20654 24140 0 _367_
rlabel metal1 20608 26350 20608 26350 0 _368_
rlabel metal1 21022 26010 21022 26010 0 _369_
rlabel metal1 19780 27982 19780 27982 0 _370_
rlabel metal1 21206 26894 21206 26894 0 _371_
rlabel metal1 21022 26758 21022 26758 0 _372_
rlabel metal1 22310 26418 22310 26418 0 _373_
rlabel metal1 21574 26384 21574 26384 0 _374_
rlabel metal1 20010 27914 20010 27914 0 _375_
rlabel metal1 20976 27438 20976 27438 0 _376_
rlabel metal1 20378 27404 20378 27404 0 _377_
rlabel metal1 19918 27404 19918 27404 0 _378_
rlabel metal1 20286 26996 20286 26996 0 _379_
rlabel metal1 20838 27098 20838 27098 0 _380_
rlabel metal1 20102 29274 20102 29274 0 _381_
rlabel metal1 20332 29138 20332 29138 0 _382_
rlabel metal2 20378 29886 20378 29886 0 _383_
rlabel metal1 21344 29138 21344 29138 0 _384_
rlabel metal1 20677 29002 20677 29002 0 _385_
rlabel metal1 20746 28560 20746 28560 0 _386_
rlabel metal1 20148 29750 20148 29750 0 _387_
rlabel metal1 21068 29818 21068 29818 0 _388_
rlabel metal1 20930 29274 20930 29274 0 _389_
rlabel metal1 21620 31382 21620 31382 0 _390_
rlabel metal1 20654 32266 20654 32266 0 _391_
rlabel metal1 20378 31348 20378 31348 0 _392_
rlabel viali 20562 29619 20562 29619 0 _393_
rlabel metal2 20194 30430 20194 30430 0 _394_
rlabel metal1 20746 32198 20746 32198 0 _395_
rlabel metal1 19642 31314 19642 31314 0 _396_
rlabel metal1 19136 31450 19136 31450 0 _397_
rlabel metal1 20884 31994 20884 31994 0 _398_
rlabel metal1 21206 31892 21206 31892 0 _399_
rlabel metal1 20976 31926 20976 31926 0 _400_
rlabel metal1 22908 23086 22908 23086 0 _401_
rlabel metal1 24886 25364 24886 25364 0 _402_
rlabel metal1 23552 26554 23552 26554 0 _403_
rlabel metal1 23966 25772 23966 25772 0 _404_
rlabel metal1 23460 27506 23460 27506 0 _405_
rlabel metal1 24242 27404 24242 27404 0 _406_
rlabel metal1 23230 29614 23230 29614 0 _407_
rlabel metal2 23138 27914 23138 27914 0 _408_
rlabel metal1 23598 29818 23598 29818 0 _409_
rlabel metal1 22954 29274 22954 29274 0 _410_
rlabel metal1 24426 30736 24426 30736 0 _411_
rlabel metal1 23552 29614 23552 29614 0 _412_
rlabel metal1 25070 31280 25070 31280 0 _413_
rlabel metal1 19090 22678 19090 22678 0 _414_
rlabel metal1 18262 20910 18262 20910 0 _415_
rlabel metal1 17710 21488 17710 21488 0 _416_
rlabel metal1 17848 20230 17848 20230 0 _417_
rlabel metal1 17434 20468 17434 20468 0 _418_
rlabel metal1 18170 18938 18170 18938 0 _419_
rlabel metal1 17802 19278 17802 19278 0 _420_
rlabel metal1 17434 18054 17434 18054 0 _421_
rlabel metal1 17204 18394 17204 18394 0 _422_
rlabel via1 18444 17170 18444 17170 0 _423_
rlabel metal1 17342 17680 17342 17680 0 _424_
rlabel metal1 18170 16082 18170 16082 0 _425_
rlabel metal1 34730 21998 34730 21998 0 clk
rlabel metal2 29946 32912 29946 32912 0 debounce0_a.button_hist\[0\]
rlabel metal1 29992 32470 29992 32470 0 debounce0_a.button_hist\[1\]
rlabel metal1 29946 33354 29946 33354 0 debounce0_a.button_hist\[2\]
rlabel metal2 30038 32130 30038 32130 0 debounce0_a.button_hist\[3\]
rlabel metal1 31372 31994 31372 31994 0 debounce0_a.button_hist\[4\]
rlabel metal2 30682 30396 30682 30396 0 debounce0_a.button_hist\[5\]
rlabel metal1 31556 31858 31556 31858 0 debounce0_a.button_hist\[6\]
rlabel metal1 31004 31450 31004 31450 0 debounce0_a.button_hist\[7\]
rlabel metal1 30912 29478 30912 29478 0 debounce0_a.debounced
rlabel metal1 17411 17578 17411 17578 0 debounce0_a.reset
rlabel metal1 32062 28186 32062 28186 0 debounce0_b.button_hist\[0\]
rlabel metal2 32154 28220 32154 28220 0 debounce0_b.button_hist\[1\]
rlabel metal1 31234 28118 31234 28118 0 debounce0_b.button_hist\[2\]
rlabel metal2 32430 27846 32430 27846 0 debounce0_b.button_hist\[3\]
rlabel metal1 32706 25874 32706 25874 0 debounce0_b.button_hist\[4\]
rlabel metal1 31556 24786 31556 24786 0 debounce0_b.button_hist\[5\]
rlabel metal1 32660 24786 32660 24786 0 debounce0_b.button_hist\[6\]
rlabel metal1 33028 24582 33028 24582 0 debounce0_b.button_hist\[7\]
rlabel metal1 28382 24718 28382 24718 0 debounce0_b.debounced
rlabel metal1 32200 16422 32200 16422 0 debounce1_a.button_hist\[0\]
rlabel metal1 31878 18802 31878 18802 0 debounce1_a.button_hist\[1\]
rlabel metal1 32108 18734 32108 18734 0 debounce1_a.button_hist\[2\]
rlabel metal1 32522 19822 32522 19822 0 debounce1_a.button_hist\[3\]
rlabel metal1 30406 21046 30406 21046 0 debounce1_a.button_hist\[4\]
rlabel metal1 31050 21964 31050 21964 0 debounce1_a.button_hist\[5\]
rlabel metal2 31786 22236 31786 22236 0 debounce1_a.button_hist\[6\]
rlabel metal1 33488 21658 33488 21658 0 debounce1_a.button_hist\[7\]
rlabel metal2 25622 21182 25622 21182 0 debounce1_a.debounced
rlabel metal1 26128 22610 26128 22610 0 debounce1_b.button_hist\[0\]
rlabel metal1 27324 22066 27324 22066 0 debounce1_b.button_hist\[1\]
rlabel metal1 27876 23086 27876 23086 0 debounce1_b.button_hist\[2\]
rlabel metal1 28106 22746 28106 22746 0 debounce1_b.button_hist\[3\]
rlabel metal1 27968 20910 27968 20910 0 debounce1_b.button_hist\[4\]
rlabel metal2 26818 20468 26818 20468 0 debounce1_b.button_hist\[5\]
rlabel metal2 27830 20740 27830 20740 0 debounce1_b.button_hist\[6\]
rlabel metal1 27876 21046 27876 21046 0 debounce1_b.button_hist\[7\]
rlabel via1 25254 21403 25254 21403 0 debounce1_b.debounced
rlabel metal2 25806 15436 25806 15436 0 debounce2_a.button_hist\[0\]
rlabel metal1 25806 15368 25806 15368 0 debounce2_a.button_hist\[1\]
rlabel metal2 25990 15572 25990 15572 0 debounce2_a.button_hist\[2\]
rlabel metal1 25990 16218 25990 16218 0 debounce2_a.button_hist\[3\]
rlabel metal1 26818 17170 26818 17170 0 debounce2_a.button_hist\[4\]
rlabel viali 25806 18259 25806 18259 0 debounce2_a.button_hist\[5\]
rlabel metal1 27278 17238 27278 17238 0 debounce2_a.button_hist\[6\]
rlabel metal1 26910 16966 26910 16966 0 debounce2_a.button_hist\[7\]
rlabel metal1 25622 19482 25622 19482 0 debounce2_a.debounced
rlabel metal1 29578 16762 29578 16762 0 debounce2_b.button_hist\[0\]
rlabel metal2 29118 16048 29118 16048 0 debounce2_b.button_hist\[1\]
rlabel metal1 29670 16422 29670 16422 0 debounce2_b.button_hist\[2\]
rlabel metal1 29946 16558 29946 16558 0 debounce2_b.button_hist\[3\]
rlabel metal1 29808 17782 29808 17782 0 debounce2_b.button_hist\[4\]
rlabel metal1 29164 18802 29164 18802 0 debounce2_b.button_hist\[5\]
rlabel metal1 30406 18938 30406 18938 0 debounce2_b.button_hist\[6\]
rlabel metal1 29946 18394 29946 18394 0 debounce2_b.button_hist\[7\]
rlabel metal1 29394 20026 29394 20026 0 debounce2_b.debounced
rlabel metal3 820 39508 820 39508 0 enc0_a
rlabel metal1 34730 32402 34730 32402 0 enc0_b
rlabel metal1 34868 2414 34868 2414 0 enc1_a
rlabel metal1 16836 39406 16836 39406 0 enc1_b
rlabel metal2 46 1588 46 1588 0 enc2_a
rlabel metal2 28382 1588 28382 1588 0 enc2_b
rlabel viali 30315 24786 30315 24786 0 encoder0.old_a
rlabel metal1 29624 24922 29624 24922 0 encoder0.old_b
rlabel metal1 28244 25874 28244 25874 0 encoder0.value\[0\]
rlabel metal1 25806 26282 25806 26282 0 encoder0.value\[1\]
rlabel metal1 25622 26928 25622 26928 0 encoder0.value\[2\]
rlabel metal2 25530 27948 25530 27948 0 encoder0.value\[3\]
rlabel via1 25713 29614 25713 29614 0 encoder0.value\[4\]
rlabel metal1 26818 30226 26818 30226 0 encoder0.value\[5\]
rlabel metal2 25714 30396 25714 30396 0 encoder0.value\[6\]
rlabel metal1 26542 32402 26542 32402 0 encoder0.value\[7\]
rlabel metal2 25346 21386 25346 21386 0 encoder1.old_a
rlabel metal1 25438 20842 25438 20842 0 encoder1.old_b
rlabel metal1 20792 21454 20792 21454 0 encoder1.value\[0\]
rlabel metal1 21206 20910 21206 20910 0 encoder1.value\[1\]
rlabel metal1 21298 18836 21298 18836 0 encoder1.value\[2\]
rlabel metal1 20562 19482 20562 19482 0 encoder1.value\[3\]
rlabel metal2 21666 18496 21666 18496 0 encoder1.value\[4\]
rlabel metal1 19458 17748 19458 17748 0 encoder1.value\[5\]
rlabel metal1 21206 16524 21206 16524 0 encoder1.value\[6\]
rlabel metal1 20470 16048 20470 16048 0 encoder1.value\[7\]
rlabel metal1 23138 24786 23138 24786 0 encoder2.old_a
rlabel metal1 22034 24106 22034 24106 0 encoder2.old_b
rlabel metal1 19320 25262 19320 25262 0 encoder2.value\[0\]
rlabel metal1 20470 24106 20470 24106 0 encoder2.value\[1\]
rlabel metal1 19688 26758 19688 26758 0 encoder2.value\[2\]
rlabel metal1 19228 27438 19228 27438 0 encoder2.value\[3\]
rlabel metal1 21390 28730 21390 28730 0 encoder2.value\[4\]
rlabel metal1 19366 29614 19366 29614 0 encoder2.value\[5\]
rlabel metal1 20378 32334 20378 32334 0 encoder2.value\[6\]
rlabel metal1 21574 31824 21574 31824 0 encoder2.value\[7\]
rlabel metal1 23874 26894 23874 26894 0 net1
rlabel metal2 19642 4657 19642 4657 0 net10
rlabel metal2 18262 30430 18262 30430 0 net11
rlabel metal1 34178 11798 34178 11798 0 net12
rlabel metal1 19688 19346 19688 19346 0 net13
rlabel metal2 17894 20366 17894 20366 0 net14
rlabel metal1 19826 15028 19826 15028 0 net15
rlabel metal1 24380 17646 24380 17646 0 net16
rlabel metal1 31142 18122 31142 18122 0 net17
rlabel metal1 29348 20910 29348 20910 0 net18
rlabel metal1 29992 21522 29992 21522 0 net19
rlabel metal2 1610 36380 1610 36380 0 net2
rlabel metal1 27094 18734 27094 18734 0 net20
rlabel metal1 19826 26894 19826 26894 0 net21
rlabel metal1 17112 31790 17112 31790 0 net22
rlabel metal1 23368 31314 23368 31314 0 net23
rlabel metal1 25484 25874 25484 25874 0 net24
rlabel metal1 29348 32402 29348 32402 0 net25
rlabel metal1 31924 31314 31924 31314 0 net26
rlabel metal1 15594 17238 15594 17238 0 net27
rlabel metal2 9062 1027 9062 1027 0 net28
rlabel metal1 26496 39610 26496 39610 0 net29
rlabel via1 32069 31790 32069 31790 0 net3
rlabel metal3 1050 9588 1050 9588 0 net30
rlabel metal3 820 19788 820 19788 0 net31
rlabel metal1 32936 2618 32936 2618 0 net4
rlabel metal1 17342 39270 17342 39270 0 net5
rlabel metal2 1702 8398 1702 8398 0 net6
rlabel metal1 28290 14382 28290 14382 0 net7
rlabel metal1 25024 12206 25024 12206 0 net8
rlabel metal2 34178 34952 34178 34952 0 net9
rlabel metal2 23598 25432 23598 25432 0 pwm0.count\[0\]
rlabel via1 24614 26554 24614 26554 0 pwm0.count\[1\]
rlabel metal2 24794 26622 24794 26622 0 pwm0.count\[2\]
rlabel metal1 25116 28186 25116 28186 0 pwm0.count\[3\]
rlabel metal1 24058 28492 24058 28492 0 pwm0.count\[4\]
rlabel metal1 24058 29784 24058 29784 0 pwm0.count\[5\]
rlabel metal1 24794 29614 24794 29614 0 pwm0.count\[6\]
rlabel metal2 24794 30906 24794 30906 0 pwm0.count\[7\]
rlabel metal1 34960 39610 34960 39610 0 pwm0_out
rlabel metal1 18860 21998 18860 21998 0 pwm1.count\[0\]
rlabel via1 18631 21998 18631 21998 0 pwm1.count\[1\]
rlabel metal2 19642 20944 19642 20944 0 pwm1.count\[2\]
rlabel metal1 17894 20332 17894 20332 0 pwm1.count\[3\]
rlabel metal1 19412 18734 19412 18734 0 pwm1.count\[4\]
rlabel metal1 18906 18360 18906 18360 0 pwm1.count\[5\]
rlabel metal1 18400 17306 18400 17306 0 pwm1.count\[6\]
rlabel metal1 18676 17102 18676 17102 0 pwm1.count\[7\]
rlabel metal2 18722 959 18722 959 0 pwm1_out
rlabel metal1 18254 26010 18254 26010 0 pwm2.count\[0\]
rlabel metal1 18446 25806 18446 25806 0 pwm2.count\[1\]
rlabel metal1 17802 26554 17802 26554 0 pwm2.count\[2\]
rlabel metal1 18308 28050 18308 28050 0 pwm2.count\[3\]
rlabel metal1 18676 28526 18676 28526 0 pwm2.count\[4\]
rlabel metal1 17848 30362 17848 30362 0 pwm2.count\[5\]
rlabel metal2 19366 30753 19366 30753 0 pwm2.count\[6\]
rlabel metal1 18308 31994 18308 31994 0 pwm2.count\[7\]
rlabel metal3 820 29988 820 29988 0 pwm2_out
rlabel metal1 7176 39406 7176 39406 0 reset
rlabel metal1 34500 11594 34500 11594 0 sync
<< properties >>
string FIXED_BBOX 0 0 36000 42000
<< end >>
